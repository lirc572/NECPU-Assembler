`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Company: lirc572
// Engineer: lirc572
// 
// Create Date: 
// Design Name: NECPU
// Module Name: InstMem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module instMem (
    input  [31:0]  address,
    output reg [31:0] inst
  );
  always @ (address) begin
    inst = 32'd0;
    case (address)
      0: inst = 32'd268468224;
      1: inst = 32'd201342944;
      2: inst = 32'd203486871;
      3: inst = 32'd136314880;
      4: inst = 32'd268468224;
      5: inst = 32'd201342945;
      6: inst = 32'd203484855;
      7: inst = 32'd136314880;
      8: inst = 32'd268468224;
      9: inst = 32'd201342946;
      10: inst = 32'd203484854;
      11: inst = 32'd136314880;
      12: inst = 32'd268468224;
      13: inst = 32'd201342947;
      14: inst = 32'd203484886;
      15: inst = 32'd136314880;
      16: inst = 32'd268468224;
      17: inst = 32'd201342948;
      18: inst = 32'd203482837;
      19: inst = 32'd136314880;
      20: inst = 32'd268468224;
      21: inst = 32'd201342949;
      22: inst = 32'd203482837;
      23: inst = 32'd136314880;
      24: inst = 32'd268468224;
      25: inst = 32'd201342950;
      26: inst = 32'd203484885;
      27: inst = 32'd136314880;
      28: inst = 32'd268468224;
      29: inst = 32'd201342951;
      30: inst = 32'd203484854;
      31: inst = 32'd136314880;
      32: inst = 32'd268468224;
      33: inst = 32'd201342952;
      34: inst = 32'd203486902;
      35: inst = 32'd136314880;
      36: inst = 32'd268468224;
      37: inst = 32'd201342953;
      38: inst = 32'd203486871;
      39: inst = 32'd136314880;
      40: inst = 32'd268468224;
      41: inst = 32'd201342954;
      42: inst = 32'd203486871;
      43: inst = 32'd136314880;
      44: inst = 32'd268468224;
      45: inst = 32'd201342955;
      46: inst = 32'd203469934;
      47: inst = 32'd136314880;
      48: inst = 32'd268468224;
      49: inst = 32'd201342956;
      50: inst = 32'd203486870;
      51: inst = 32'd136314880;
      52: inst = 32'd268468224;
      53: inst = 32'd201342957;
      54: inst = 32'd203484854;
      55: inst = 32'd136314880;
      56: inst = 32'd268468224;
      57: inst = 32'd201342958;
      58: inst = 32'd203484853;
      59: inst = 32'd136314880;
      60: inst = 32'd268468224;
      61: inst = 32'd201342959;
      62: inst = 32'd203484885;
      63: inst = 32'd136314880;
      64: inst = 32'd268468224;
      65: inst = 32'd201342960;
      66: inst = 32'd203484854;
      67: inst = 32'd136314880;
      68: inst = 32'd268468224;
      69: inst = 32'd201342961;
      70: inst = 32'd203484854;
      71: inst = 32'd136314880;
      72: inst = 32'd268468224;
      73: inst = 32'd201342962;
      74: inst = 32'd203484854;
      75: inst = 32'd136314880;
      76: inst = 32'd268468224;
      77: inst = 32'd201342963;
      78: inst = 32'd203484855;
      79: inst = 32'd136314880;
      80: inst = 32'd268468224;
      81: inst = 32'd201342964;
      82: inst = 32'd203484855;
      83: inst = 32'd136314880;
      84: inst = 32'd268468224;
      85: inst = 32'd201342965;
      86: inst = 32'd203484855;
      87: inst = 32'd136314880;
      88: inst = 32'd268468224;
      89: inst = 32'd201342966;
      90: inst = 32'd203484854;
      91: inst = 32'd136314880;
      92: inst = 32'd268468224;
      93: inst = 32'd201342967;
      94: inst = 32'd203484854;
      95: inst = 32'd136314880;
      96: inst = 32'd268468224;
      97: inst = 32'd201342968;
      98: inst = 32'd203486934;
      99: inst = 32'd136314880;
      100: inst = 32'd268468224;
      101: inst = 32'd201342969;
      102: inst = 32'd203484821;
      103: inst = 32'd136314880;
      104: inst = 32'd268468224;
      105: inst = 32'd201342970;
      106: inst = 32'd203486934;
      107: inst = 32'd136314880;
      108: inst = 32'd268468224;
      109: inst = 32'd201342971;
      110: inst = 32'd203484821;
      111: inst = 32'd136314880;
      112: inst = 32'd268468224;
      113: inst = 32'd201342972;
      114: inst = 32'd203484853;
      115: inst = 32'd136314880;
      116: inst = 32'd268468224;
      117: inst = 32'd201342973;
      118: inst = 32'd203484821;
      119: inst = 32'd136314880;
      120: inst = 32'd268468224;
      121: inst = 32'd201342974;
      122: inst = 32'd203484887;
      123: inst = 32'd136314880;
      124: inst = 32'd268468224;
      125: inst = 32'd201342975;
      126: inst = 32'd203484886;
      127: inst = 32'd136314880;
      128: inst = 32'd268468224;
      129: inst = 32'd201342976;
      130: inst = 32'd203484823;
      131: inst = 32'd136314880;
      132: inst = 32'd268468224;
      133: inst = 32'd201342977;
      134: inst = 32'd203484823;
      135: inst = 32'd136314880;
      136: inst = 32'd268468224;
      137: inst = 32'd201342978;
      138: inst = 32'd203484823;
      139: inst = 32'd136314880;
      140: inst = 32'd268468224;
      141: inst = 32'd201342979;
      142: inst = 32'd203484823;
      143: inst = 32'd136314880;
      144: inst = 32'd268468224;
      145: inst = 32'd201342980;
      146: inst = 32'd203484823;
      147: inst = 32'd136314880;
      148: inst = 32'd268468224;
      149: inst = 32'd201342981;
      150: inst = 32'd203484823;
      151: inst = 32'd136314880;
      152: inst = 32'd268468224;
      153: inst = 32'd201342982;
      154: inst = 32'd203484823;
      155: inst = 32'd136314880;
      156: inst = 32'd268468224;
      157: inst = 32'd201342983;
      158: inst = 32'd203484823;
      159: inst = 32'd136314880;
      160: inst = 32'd268468224;
      161: inst = 32'd201342984;
      162: inst = 32'd203484823;
      163: inst = 32'd136314880;
      164: inst = 32'd268468224;
      165: inst = 32'd201342985;
      166: inst = 32'd203484823;
      167: inst = 32'd136314880;
      168: inst = 32'd268468224;
      169: inst = 32'd201342986;
      170: inst = 32'd203484823;
      171: inst = 32'd136314880;
      172: inst = 32'd268468224;
      173: inst = 32'd201342987;
      174: inst = 32'd203484823;
      175: inst = 32'd136314880;
      176: inst = 32'd268468224;
      177: inst = 32'd201342988;
      178: inst = 32'd203484823;
      179: inst = 32'd136314880;
      180: inst = 32'd268468224;
      181: inst = 32'd201342989;
      182: inst = 32'd203484823;
      183: inst = 32'd136314880;
      184: inst = 32'd268468224;
      185: inst = 32'd201342990;
      186: inst = 32'd203484823;
      187: inst = 32'd136314880;
      188: inst = 32'd268468224;
      189: inst = 32'd201342991;
      190: inst = 32'd203484823;
      191: inst = 32'd136314880;
      192: inst = 32'd268468224;
      193: inst = 32'd201342992;
      194: inst = 32'd203484823;
      195: inst = 32'd136314880;
      196: inst = 32'd268468224;
      197: inst = 32'd201342993;
      198: inst = 32'd203484823;
      199: inst = 32'd136314880;
      200: inst = 32'd268468224;
      201: inst = 32'd201342994;
      202: inst = 32'd203484823;
      203: inst = 32'd136314880;
      204: inst = 32'd268468224;
      205: inst = 32'd201342995;
      206: inst = 32'd203484823;
      207: inst = 32'd136314880;
      208: inst = 32'd268468224;
      209: inst = 32'd201342996;
      210: inst = 32'd203484823;
      211: inst = 32'd136314880;
      212: inst = 32'd268468224;
      213: inst = 32'd201342997;
      214: inst = 32'd203484823;
      215: inst = 32'd136314880;
      216: inst = 32'd268468224;
      217: inst = 32'd201342998;
      218: inst = 32'd203484823;
      219: inst = 32'd136314880;
      220: inst = 32'd268468224;
      221: inst = 32'd201342999;
      222: inst = 32'd203484823;
      223: inst = 32'd136314880;
      224: inst = 32'd268468224;
      225: inst = 32'd201343000;
      226: inst = 32'd203484823;
      227: inst = 32'd136314880;
      228: inst = 32'd268468224;
      229: inst = 32'd201343001;
      230: inst = 32'd203484823;
      231: inst = 32'd136314880;
      232: inst = 32'd268468224;
      233: inst = 32'd201343002;
      234: inst = 32'd203484823;
      235: inst = 32'd136314880;
      236: inst = 32'd268468224;
      237: inst = 32'd201343003;
      238: inst = 32'd203484823;
      239: inst = 32'd136314880;
      240: inst = 32'd268468224;
      241: inst = 32'd201343004;
      242: inst = 32'd203484823;
      243: inst = 32'd136314880;
      244: inst = 32'd268468224;
      245: inst = 32'd201343005;
      246: inst = 32'd203484823;
      247: inst = 32'd136314880;
      248: inst = 32'd268468224;
      249: inst = 32'd201343006;
      250: inst = 32'd203484823;
      251: inst = 32'd136314880;
      252: inst = 32'd268468224;
      253: inst = 32'd201343007;
      254: inst = 32'd203484823;
      255: inst = 32'd136314880;
      256: inst = 32'd268468224;
      257: inst = 32'd201343008;
      258: inst = 32'd203484886;
      259: inst = 32'd136314880;
      260: inst = 32'd268468224;
      261: inst = 32'd201343009;
      262: inst = 32'd203484887;
      263: inst = 32'd136314880;
      264: inst = 32'd268468224;
      265: inst = 32'd201343010;
      266: inst = 32'd203484821;
      267: inst = 32'd136314880;
      268: inst = 32'd268468224;
      269: inst = 32'd201343011;
      270: inst = 32'd203484853;
      271: inst = 32'd136314880;
      272: inst = 32'd268468224;
      273: inst = 32'd201343012;
      274: inst = 32'd203484821;
      275: inst = 32'd136314880;
      276: inst = 32'd268468224;
      277: inst = 32'd201343013;
      278: inst = 32'd203486934;
      279: inst = 32'd136314880;
      280: inst = 32'd268468224;
      281: inst = 32'd201343014;
      282: inst = 32'd203484821;
      283: inst = 32'd136314880;
      284: inst = 32'd268468224;
      285: inst = 32'd201343015;
      286: inst = 32'd203486902;
      287: inst = 32'd136314880;
      288: inst = 32'd268468224;
      289: inst = 32'd201343016;
      290: inst = 32'd203484854;
      291: inst = 32'd136314880;
      292: inst = 32'd268468224;
      293: inst = 32'd201343017;
      294: inst = 32'd203484854;
      295: inst = 32'd136314880;
      296: inst = 32'd268468224;
      297: inst = 32'd201343018;
      298: inst = 32'd203484855;
      299: inst = 32'd136314880;
      300: inst = 32'd268468224;
      301: inst = 32'd201343019;
      302: inst = 32'd203484855;
      303: inst = 32'd136314880;
      304: inst = 32'd268468224;
      305: inst = 32'd201343020;
      306: inst = 32'd203484855;
      307: inst = 32'd136314880;
      308: inst = 32'd268468224;
      309: inst = 32'd201343021;
      310: inst = 32'd203484854;
      311: inst = 32'd136314880;
      312: inst = 32'd268468224;
      313: inst = 32'd201343022;
      314: inst = 32'd203484854;
      315: inst = 32'd136314880;
      316: inst = 32'd268468224;
      317: inst = 32'd201343023;
      318: inst = 32'd203484854;
      319: inst = 32'd136314880;
      320: inst = 32'd268468224;
      321: inst = 32'd201343024;
      322: inst = 32'd203484854;
      323: inst = 32'd136314880;
      324: inst = 32'd268468224;
      325: inst = 32'd201343025;
      326: inst = 32'd203484854;
      327: inst = 32'd136314880;
      328: inst = 32'd268468224;
      329: inst = 32'd201343026;
      330: inst = 32'd203484854;
      331: inst = 32'd136314880;
      332: inst = 32'd268468224;
      333: inst = 32'd201343027;
      334: inst = 32'd203484854;
      335: inst = 32'd136314880;
      336: inst = 32'd268468224;
      337: inst = 32'd201343028;
      338: inst = 32'd203484854;
      339: inst = 32'd136314880;
      340: inst = 32'd268468224;
      341: inst = 32'd201343029;
      342: inst = 32'd203484854;
      343: inst = 32'd136314880;
      344: inst = 32'd268468224;
      345: inst = 32'd201343030;
      346: inst = 32'd203484854;
      347: inst = 32'd136314880;
      348: inst = 32'd268468224;
      349: inst = 32'd201343031;
      350: inst = 32'd203484854;
      351: inst = 32'd136314880;
      352: inst = 32'd268468224;
      353: inst = 32'd201343032;
      354: inst = 32'd203484854;
      355: inst = 32'd136314880;
      356: inst = 32'd268468224;
      357: inst = 32'd201343033;
      358: inst = 32'd203484854;
      359: inst = 32'd136314880;
      360: inst = 32'd268468224;
      361: inst = 32'd201343034;
      362: inst = 32'd203484854;
      363: inst = 32'd136314880;
      364: inst = 32'd268468224;
      365: inst = 32'd201343035;
      366: inst = 32'd203484854;
      367: inst = 32'd136314880;
      368: inst = 32'd268468224;
      369: inst = 32'd201343036;
      370: inst = 32'd203484854;
      371: inst = 32'd136314880;
      372: inst = 32'd268468224;
      373: inst = 32'd201343037;
      374: inst = 32'd203484854;
      375: inst = 32'd136314880;
      376: inst = 32'd268468224;
      377: inst = 32'd201343038;
      378: inst = 32'd203484854;
      379: inst = 32'd136314880;
      380: inst = 32'd268468224;
      381: inst = 32'd201343039;
      382: inst = 32'd203484854;
      383: inst = 32'd136314880;
      384: inst = 32'd268468224;
      385: inst = 32'd201343040;
      386: inst = 32'd203484823;
      387: inst = 32'd136314880;
      388: inst = 32'd268468224;
      389: inst = 32'd201343041;
      390: inst = 32'd203484855;
      391: inst = 32'd136314880;
      392: inst = 32'd268468224;
      393: inst = 32'd201343042;
      394: inst = 32'd203484854;
      395: inst = 32'd136314880;
      396: inst = 32'd268468224;
      397: inst = 32'd201343043;
      398: inst = 32'd203484886;
      399: inst = 32'd136314880;
      400: inst = 32'd268468224;
      401: inst = 32'd201343044;
      402: inst = 32'd203484885;
      403: inst = 32'd136314880;
      404: inst = 32'd268468224;
      405: inst = 32'd201343045;
      406: inst = 32'd203482837;
      407: inst = 32'd136314880;
      408: inst = 32'd268468224;
      409: inst = 32'd201343046;
      410: inst = 32'd203482838;
      411: inst = 32'd136314880;
      412: inst = 32'd268468224;
      413: inst = 32'd201343047;
      414: inst = 32'd203484886;
      415: inst = 32'd136314880;
      416: inst = 32'd268468224;
      417: inst = 32'd201343048;
      418: inst = 32'd203484887;
      419: inst = 32'd136314880;
      420: inst = 32'd268468224;
      421: inst = 32'd201343049;
      422: inst = 32'd203484855;
      423: inst = 32'd136314880;
      424: inst = 32'd268468224;
      425: inst = 32'd201343050;
      426: inst = 32'd203484855;
      427: inst = 32'd136314880;
      428: inst = 32'd268468224;
      429: inst = 32'd201343051;
      430: inst = 32'd203465871;
      431: inst = 32'd136314880;
      432: inst = 32'd268468224;
      433: inst = 32'd201343052;
      434: inst = 32'd203482839;
      435: inst = 32'd136314880;
      436: inst = 32'd268468224;
      437: inst = 32'd201343053;
      438: inst = 32'd203482838;
      439: inst = 32'd136314880;
      440: inst = 32'd268468224;
      441: inst = 32'd201343054;
      442: inst = 32'd203482838;
      443: inst = 32'd136314880;
      444: inst = 32'd268468224;
      445: inst = 32'd201343055;
      446: inst = 32'd203482870;
      447: inst = 32'd136314880;
      448: inst = 32'd268468224;
      449: inst = 32'd201343056;
      450: inst = 32'd203484854;
      451: inst = 32'd136314880;
      452: inst = 32'd268468224;
      453: inst = 32'd201343057;
      454: inst = 32'd203484854;
      455: inst = 32'd136314880;
      456: inst = 32'd268468224;
      457: inst = 32'd201343058;
      458: inst = 32'd203484854;
      459: inst = 32'd136314880;
      460: inst = 32'd268468224;
      461: inst = 32'd201343059;
      462: inst = 32'd203484855;
      463: inst = 32'd136314880;
      464: inst = 32'd268468224;
      465: inst = 32'd201343060;
      466: inst = 32'd203484855;
      467: inst = 32'd136314880;
      468: inst = 32'd268468224;
      469: inst = 32'd201343061;
      470: inst = 32'd203484855;
      471: inst = 32'd136314880;
      472: inst = 32'd268468224;
      473: inst = 32'd201343062;
      474: inst = 32'd203484854;
      475: inst = 32'd136314880;
      476: inst = 32'd268468224;
      477: inst = 32'd201343063;
      478: inst = 32'd203484854;
      479: inst = 32'd136314880;
      480: inst = 32'd268468224;
      481: inst = 32'd201343064;
      482: inst = 32'd203484854;
      483: inst = 32'd136314880;
      484: inst = 32'd268468224;
      485: inst = 32'd201343065;
      486: inst = 32'd203484821;
      487: inst = 32'd136314880;
      488: inst = 32'd268468224;
      489: inst = 32'd201343066;
      490: inst = 32'd203486934;
      491: inst = 32'd136314880;
      492: inst = 32'd268468224;
      493: inst = 32'd201343067;
      494: inst = 32'd203486934;
      495: inst = 32'd136314880;
      496: inst = 32'd268468224;
      497: inst = 32'd201343068;
      498: inst = 32'd203486934;
      499: inst = 32'd136314880;
      500: inst = 32'd268468224;
      501: inst = 32'd201343069;
      502: inst = 32'd203484854;
      503: inst = 32'd136314880;
      504: inst = 32'd268468224;
      505: inst = 32'd201343070;
      506: inst = 32'd203484854;
      507: inst = 32'd136314880;
      508: inst = 32'd268468224;
      509: inst = 32'd201343071;
      510: inst = 32'd203482806;
      511: inst = 32'd136314880;
      512: inst = 32'd268468224;
      513: inst = 32'd201343072;
      514: inst = 32'd203484854;
      515: inst = 32'd136314880;
      516: inst = 32'd268468224;
      517: inst = 32'd201343073;
      518: inst = 32'd203484854;
      519: inst = 32'd136314880;
      520: inst = 32'd268468224;
      521: inst = 32'd201343074;
      522: inst = 32'd203484854;
      523: inst = 32'd136314880;
      524: inst = 32'd268468224;
      525: inst = 32'd201343075;
      526: inst = 32'd203484854;
      527: inst = 32'd136314880;
      528: inst = 32'd268468224;
      529: inst = 32'd201343076;
      530: inst = 32'd203484854;
      531: inst = 32'd136314880;
      532: inst = 32'd268468224;
      533: inst = 32'd201343077;
      534: inst = 32'd203484854;
      535: inst = 32'd136314880;
      536: inst = 32'd268468224;
      537: inst = 32'd201343078;
      538: inst = 32'd203484854;
      539: inst = 32'd136314880;
      540: inst = 32'd268468224;
      541: inst = 32'd201343079;
      542: inst = 32'd203484854;
      543: inst = 32'd136314880;
      544: inst = 32'd268468224;
      545: inst = 32'd201343080;
      546: inst = 32'd203484854;
      547: inst = 32'd136314880;
      548: inst = 32'd268468224;
      549: inst = 32'd201343081;
      550: inst = 32'd203484854;
      551: inst = 32'd136314880;
      552: inst = 32'd268468224;
      553: inst = 32'd201343082;
      554: inst = 32'd203484854;
      555: inst = 32'd136314880;
      556: inst = 32'd268468224;
      557: inst = 32'd201343083;
      558: inst = 32'd203484854;
      559: inst = 32'd136314880;
      560: inst = 32'd268468224;
      561: inst = 32'd201343084;
      562: inst = 32'd203484854;
      563: inst = 32'd136314880;
      564: inst = 32'd268468224;
      565: inst = 32'd201343085;
      566: inst = 32'd203484854;
      567: inst = 32'd136314880;
      568: inst = 32'd268468224;
      569: inst = 32'd201343086;
      570: inst = 32'd203484854;
      571: inst = 32'd136314880;
      572: inst = 32'd268468224;
      573: inst = 32'd201343087;
      574: inst = 32'd203484854;
      575: inst = 32'd136314880;
      576: inst = 32'd268468224;
      577: inst = 32'd201343088;
      578: inst = 32'd203484854;
      579: inst = 32'd136314880;
      580: inst = 32'd268468224;
      581: inst = 32'd201343089;
      582: inst = 32'd203484854;
      583: inst = 32'd136314880;
      584: inst = 32'd268468224;
      585: inst = 32'd201343090;
      586: inst = 32'd203484854;
      587: inst = 32'd136314880;
      588: inst = 32'd268468224;
      589: inst = 32'd201343091;
      590: inst = 32'd203484854;
      591: inst = 32'd136314880;
      592: inst = 32'd268468224;
      593: inst = 32'd201343092;
      594: inst = 32'd203484854;
      595: inst = 32'd136314880;
      596: inst = 32'd268468224;
      597: inst = 32'd201343093;
      598: inst = 32'd203484854;
      599: inst = 32'd136314880;
      600: inst = 32'd268468224;
      601: inst = 32'd201343094;
      602: inst = 32'd203484854;
      603: inst = 32'd136314880;
      604: inst = 32'd268468224;
      605: inst = 32'd201343095;
      606: inst = 32'd203484854;
      607: inst = 32'd136314880;
      608: inst = 32'd268468224;
      609: inst = 32'd201343096;
      610: inst = 32'd203484854;
      611: inst = 32'd136314880;
      612: inst = 32'd268468224;
      613: inst = 32'd201343097;
      614: inst = 32'd203484854;
      615: inst = 32'd136314880;
      616: inst = 32'd268468224;
      617: inst = 32'd201343098;
      618: inst = 32'd203484854;
      619: inst = 32'd136314880;
      620: inst = 32'd268468224;
      621: inst = 32'd201343099;
      622: inst = 32'd203484854;
      623: inst = 32'd136314880;
      624: inst = 32'd268468224;
      625: inst = 32'd201343100;
      626: inst = 32'd203484854;
      627: inst = 32'd136314880;
      628: inst = 32'd268468224;
      629: inst = 32'd201343101;
      630: inst = 32'd203484854;
      631: inst = 32'd136314880;
      632: inst = 32'd268468224;
      633: inst = 32'd201343102;
      634: inst = 32'd203484854;
      635: inst = 32'd136314880;
      636: inst = 32'd268468224;
      637: inst = 32'd201343103;
      638: inst = 32'd203484854;
      639: inst = 32'd136314880;
      640: inst = 32'd268468224;
      641: inst = 32'd201343104;
      642: inst = 32'd203482806;
      643: inst = 32'd136314880;
      644: inst = 32'd268468224;
      645: inst = 32'd201343105;
      646: inst = 32'd203484854;
      647: inst = 32'd136314880;
      648: inst = 32'd268468224;
      649: inst = 32'd201343106;
      650: inst = 32'd203484854;
      651: inst = 32'd136314880;
      652: inst = 32'd268468224;
      653: inst = 32'd201343107;
      654: inst = 32'd203486934;
      655: inst = 32'd136314880;
      656: inst = 32'd268468224;
      657: inst = 32'd201343108;
      658: inst = 32'd203486934;
      659: inst = 32'd136314880;
      660: inst = 32'd268468224;
      661: inst = 32'd201343109;
      662: inst = 32'd203486934;
      663: inst = 32'd136314880;
      664: inst = 32'd268468224;
      665: inst = 32'd201343110;
      666: inst = 32'd203484821;
      667: inst = 32'd136314880;
      668: inst = 32'd268468224;
      669: inst = 32'd201343111;
      670: inst = 32'd203484822;
      671: inst = 32'd136314880;
      672: inst = 32'd268468224;
      673: inst = 32'd201343112;
      674: inst = 32'd203484854;
      675: inst = 32'd136314880;
      676: inst = 32'd268468224;
      677: inst = 32'd201343113;
      678: inst = 32'd203484854;
      679: inst = 32'd136314880;
      680: inst = 32'd268468224;
      681: inst = 32'd201343114;
      682: inst = 32'd203484855;
      683: inst = 32'd136314880;
      684: inst = 32'd268468224;
      685: inst = 32'd201343115;
      686: inst = 32'd203484855;
      687: inst = 32'd136314880;
      688: inst = 32'd268468224;
      689: inst = 32'd201343116;
      690: inst = 32'd203484855;
      691: inst = 32'd136314880;
      692: inst = 32'd268468224;
      693: inst = 32'd201343117;
      694: inst = 32'd203484854;
      695: inst = 32'd136314880;
      696: inst = 32'd268468224;
      697: inst = 32'd201343118;
      698: inst = 32'd203484854;
      699: inst = 32'd136314880;
      700: inst = 32'd268468224;
      701: inst = 32'd201343119;
      702: inst = 32'd203484854;
      703: inst = 32'd136314880;
      704: inst = 32'd268468224;
      705: inst = 32'd201343120;
      706: inst = 32'd203484854;
      707: inst = 32'd136314880;
      708: inst = 32'd268468224;
      709: inst = 32'd201343121;
      710: inst = 32'd203484854;
      711: inst = 32'd136314880;
      712: inst = 32'd268468224;
      713: inst = 32'd201343122;
      714: inst = 32'd203484854;
      715: inst = 32'd136314880;
      716: inst = 32'd268468224;
      717: inst = 32'd201343123;
      718: inst = 32'd203484854;
      719: inst = 32'd136314880;
      720: inst = 32'd268468224;
      721: inst = 32'd201343124;
      722: inst = 32'd203484854;
      723: inst = 32'd136314880;
      724: inst = 32'd268468224;
      725: inst = 32'd201343125;
      726: inst = 32'd203484854;
      727: inst = 32'd136314880;
      728: inst = 32'd268468224;
      729: inst = 32'd201343126;
      730: inst = 32'd203484854;
      731: inst = 32'd136314880;
      732: inst = 32'd268468224;
      733: inst = 32'd201343127;
      734: inst = 32'd203484854;
      735: inst = 32'd136314880;
      736: inst = 32'd268468224;
      737: inst = 32'd201343128;
      738: inst = 32'd203484854;
      739: inst = 32'd136314880;
      740: inst = 32'd268468224;
      741: inst = 32'd201343129;
      742: inst = 32'd203484854;
      743: inst = 32'd136314880;
      744: inst = 32'd268468224;
      745: inst = 32'd201343130;
      746: inst = 32'd203484854;
      747: inst = 32'd136314880;
      748: inst = 32'd268468224;
      749: inst = 32'd201343131;
      750: inst = 32'd203484854;
      751: inst = 32'd136314880;
      752: inst = 32'd268468224;
      753: inst = 32'd201343132;
      754: inst = 32'd203484854;
      755: inst = 32'd136314880;
      756: inst = 32'd268468224;
      757: inst = 32'd201343133;
      758: inst = 32'd203484854;
      759: inst = 32'd136314880;
      760: inst = 32'd268468224;
      761: inst = 32'd201343134;
      762: inst = 32'd203484854;
      763: inst = 32'd136314880;
      764: inst = 32'd268468224;
      765: inst = 32'd201343135;
      766: inst = 32'd203484854;
      767: inst = 32'd136314880;
      768: inst = 32'd268468224;
      769: inst = 32'd201343136;
      770: inst = 32'd203484855;
      771: inst = 32'd136314880;
      772: inst = 32'd268468224;
      773: inst = 32'd201343137;
      774: inst = 32'd203484855;
      775: inst = 32'd136314880;
      776: inst = 32'd268468224;
      777: inst = 32'd201343138;
      778: inst = 32'd203484854;
      779: inst = 32'd136314880;
      780: inst = 32'd268468224;
      781: inst = 32'd201343139;
      782: inst = 32'd203484854;
      783: inst = 32'd136314880;
      784: inst = 32'd268468224;
      785: inst = 32'd201343140;
      786: inst = 32'd203484854;
      787: inst = 32'd136314880;
      788: inst = 32'd268468224;
      789: inst = 32'd201343141;
      790: inst = 32'd203484886;
      791: inst = 32'd136314880;
      792: inst = 32'd268468224;
      793: inst = 32'd201343142;
      794: inst = 32'd203484886;
      795: inst = 32'd136314880;
      796: inst = 32'd268468224;
      797: inst = 32'd201343143;
      798: inst = 32'd203482838;
      799: inst = 32'd136314880;
      800: inst = 32'd268468224;
      801: inst = 32'd201343144;
      802: inst = 32'd203482839;
      803: inst = 32'd136314880;
      804: inst = 32'd268468224;
      805: inst = 32'd201343145;
      806: inst = 32'd203482839;
      807: inst = 32'd136314880;
      808: inst = 32'd268468224;
      809: inst = 32'd201343146;
      810: inst = 32'd203482840;
      811: inst = 32'd136314880;
      812: inst = 32'd268468224;
      813: inst = 32'd201343147;
      814: inst = 32'd203463855;
      815: inst = 32'd136314880;
      816: inst = 32'd268468224;
      817: inst = 32'd201343148;
      818: inst = 32'd203480791;
      819: inst = 32'd136314880;
      820: inst = 32'd268468224;
      821: inst = 32'd201343149;
      822: inst = 32'd203480791;
      823: inst = 32'd136314880;
      824: inst = 32'd268468224;
      825: inst = 32'd201343150;
      826: inst = 32'd203480822;
      827: inst = 32'd136314880;
      828: inst = 32'd268468224;
      829: inst = 32'd201343151;
      830: inst = 32'd203482870;
      831: inst = 32'd136314880;
      832: inst = 32'd268468224;
      833: inst = 32'd201343152;
      834: inst = 32'd203484854;
      835: inst = 32'd136314880;
      836: inst = 32'd268468224;
      837: inst = 32'd201343153;
      838: inst = 32'd203484854;
      839: inst = 32'd136314880;
      840: inst = 32'd268468224;
      841: inst = 32'd201343154;
      842: inst = 32'd203484854;
      843: inst = 32'd136314880;
      844: inst = 32'd268468224;
      845: inst = 32'd201343155;
      846: inst = 32'd203484854;
      847: inst = 32'd136314880;
      848: inst = 32'd268468224;
      849: inst = 32'd201343156;
      850: inst = 32'd203484855;
      851: inst = 32'd136314880;
      852: inst = 32'd268468224;
      853: inst = 32'd201343157;
      854: inst = 32'd203484855;
      855: inst = 32'd136314880;
      856: inst = 32'd268468224;
      857: inst = 32'd201343158;
      858: inst = 32'd203484854;
      859: inst = 32'd136314880;
      860: inst = 32'd268468224;
      861: inst = 32'd201343159;
      862: inst = 32'd203484854;
      863: inst = 32'd136314880;
      864: inst = 32'd268468224;
      865: inst = 32'd201343160;
      866: inst = 32'd203486934;
      867: inst = 32'd136314880;
      868: inst = 32'd268468224;
      869: inst = 32'd201343161;
      870: inst = 32'd203486934;
      871: inst = 32'd136314880;
      872: inst = 32'd268468224;
      873: inst = 32'd201343162;
      874: inst = 32'd203484821;
      875: inst = 32'd136314880;
      876: inst = 32'd268468224;
      877: inst = 32'd201343163;
      878: inst = 32'd203484821;
      879: inst = 32'd136314880;
      880: inst = 32'd268468224;
      881: inst = 32'd201343164;
      882: inst = 32'd203482741;
      883: inst = 32'd136314880;
      884: inst = 32'd268468224;
      885: inst = 32'd201343165;
      886: inst = 32'd203482806;
      887: inst = 32'd136314880;
      888: inst = 32'd268468224;
      889: inst = 32'd201343166;
      890: inst = 32'd203482806;
      891: inst = 32'd136314880;
      892: inst = 32'd268468224;
      893: inst = 32'd201343167;
      894: inst = 32'd203484887;
      895: inst = 32'd136314880;
      896: inst = 32'd268468224;
      897: inst = 32'd201343168;
      898: inst = 32'd203484853;
      899: inst = 32'd136314880;
      900: inst = 32'd268468224;
      901: inst = 32'd201343169;
      902: inst = 32'd203484853;
      903: inst = 32'd136314880;
      904: inst = 32'd268468224;
      905: inst = 32'd201343170;
      906: inst = 32'd203484853;
      907: inst = 32'd136314880;
      908: inst = 32'd268468224;
      909: inst = 32'd201343171;
      910: inst = 32'd203484853;
      911: inst = 32'd136314880;
      912: inst = 32'd268468224;
      913: inst = 32'd201343172;
      914: inst = 32'd203484853;
      915: inst = 32'd136314880;
      916: inst = 32'd268468224;
      917: inst = 32'd201343173;
      918: inst = 32'd203484853;
      919: inst = 32'd136314880;
      920: inst = 32'd268468224;
      921: inst = 32'd201343174;
      922: inst = 32'd203484853;
      923: inst = 32'd136314880;
      924: inst = 32'd268468224;
      925: inst = 32'd201343175;
      926: inst = 32'd203484853;
      927: inst = 32'd136314880;
      928: inst = 32'd268468224;
      929: inst = 32'd201343176;
      930: inst = 32'd203484853;
      931: inst = 32'd136314880;
      932: inst = 32'd268468224;
      933: inst = 32'd201343177;
      934: inst = 32'd203484853;
      935: inst = 32'd136314880;
      936: inst = 32'd268468224;
      937: inst = 32'd201343178;
      938: inst = 32'd203484853;
      939: inst = 32'd136314880;
      940: inst = 32'd268468224;
      941: inst = 32'd201343179;
      942: inst = 32'd203484853;
      943: inst = 32'd136314880;
      944: inst = 32'd268468224;
      945: inst = 32'd201343180;
      946: inst = 32'd203484853;
      947: inst = 32'd136314880;
      948: inst = 32'd268468224;
      949: inst = 32'd201343181;
      950: inst = 32'd203484853;
      951: inst = 32'd136314880;
      952: inst = 32'd268468224;
      953: inst = 32'd201343182;
      954: inst = 32'd203484853;
      955: inst = 32'd136314880;
      956: inst = 32'd268468224;
      957: inst = 32'd201343183;
      958: inst = 32'd203484853;
      959: inst = 32'd136314880;
      960: inst = 32'd268468224;
      961: inst = 32'd201343184;
      962: inst = 32'd203484853;
      963: inst = 32'd136314880;
      964: inst = 32'd268468224;
      965: inst = 32'd201343185;
      966: inst = 32'd203484853;
      967: inst = 32'd136314880;
      968: inst = 32'd268468224;
      969: inst = 32'd201343186;
      970: inst = 32'd203484853;
      971: inst = 32'd136314880;
      972: inst = 32'd268468224;
      973: inst = 32'd201343187;
      974: inst = 32'd203484853;
      975: inst = 32'd136314880;
      976: inst = 32'd268468224;
      977: inst = 32'd201343188;
      978: inst = 32'd203484853;
      979: inst = 32'd136314880;
      980: inst = 32'd268468224;
      981: inst = 32'd201343189;
      982: inst = 32'd203484853;
      983: inst = 32'd136314880;
      984: inst = 32'd268468224;
      985: inst = 32'd201343190;
      986: inst = 32'd203484853;
      987: inst = 32'd136314880;
      988: inst = 32'd268468224;
      989: inst = 32'd201343191;
      990: inst = 32'd203484853;
      991: inst = 32'd136314880;
      992: inst = 32'd268468224;
      993: inst = 32'd201343192;
      994: inst = 32'd203484853;
      995: inst = 32'd136314880;
      996: inst = 32'd268468224;
      997: inst = 32'd201343193;
      998: inst = 32'd203484853;
      999: inst = 32'd136314880;
      1000: inst = 32'd268468224;
      1001: inst = 32'd201343194;
      1002: inst = 32'd203484853;
      1003: inst = 32'd136314880;
      1004: inst = 32'd268468224;
      1005: inst = 32'd201343195;
      1006: inst = 32'd203484853;
      1007: inst = 32'd136314880;
      1008: inst = 32'd268468224;
      1009: inst = 32'd201343196;
      1010: inst = 32'd203484853;
      1011: inst = 32'd136314880;
      1012: inst = 32'd268468224;
      1013: inst = 32'd201343197;
      1014: inst = 32'd203484853;
      1015: inst = 32'd136314880;
      1016: inst = 32'd268468224;
      1017: inst = 32'd201343198;
      1018: inst = 32'd203484853;
      1019: inst = 32'd136314880;
      1020: inst = 32'd268468224;
      1021: inst = 32'd201343199;
      1022: inst = 32'd203484853;
      1023: inst = 32'd136314880;
      1024: inst = 32'd268468224;
      1025: inst = 32'd201343200;
      1026: inst = 32'd203484887;
      1027: inst = 32'd136314880;
      1028: inst = 32'd268468224;
      1029: inst = 32'd201343201;
      1030: inst = 32'd203482806;
      1031: inst = 32'd136314880;
      1032: inst = 32'd268468224;
      1033: inst = 32'd201343202;
      1034: inst = 32'd203482806;
      1035: inst = 32'd136314880;
      1036: inst = 32'd268468224;
      1037: inst = 32'd201343203;
      1038: inst = 32'd203482741;
      1039: inst = 32'd136314880;
      1040: inst = 32'd268468224;
      1041: inst = 32'd201343204;
      1042: inst = 32'd203484821;
      1043: inst = 32'd136314880;
      1044: inst = 32'd268468224;
      1045: inst = 32'd201343205;
      1046: inst = 32'd203484821;
      1047: inst = 32'd136314880;
      1048: inst = 32'd268468224;
      1049: inst = 32'd201343206;
      1050: inst = 32'd203486902;
      1051: inst = 32'd136314880;
      1052: inst = 32'd268468224;
      1053: inst = 32'd201343207;
      1054: inst = 32'd203486934;
      1055: inst = 32'd136314880;
      1056: inst = 32'd268468224;
      1057: inst = 32'd201343208;
      1058: inst = 32'd203484854;
      1059: inst = 32'd136314880;
      1060: inst = 32'd268468224;
      1061: inst = 32'd201343209;
      1062: inst = 32'd203484854;
      1063: inst = 32'd136314880;
      1064: inst = 32'd268468224;
      1065: inst = 32'd201343210;
      1066: inst = 32'd203484855;
      1067: inst = 32'd136314880;
      1068: inst = 32'd268468224;
      1069: inst = 32'd201343211;
      1070: inst = 32'd203484855;
      1071: inst = 32'd136314880;
      1072: inst = 32'd268468224;
      1073: inst = 32'd201343212;
      1074: inst = 32'd203484854;
      1075: inst = 32'd136314880;
      1076: inst = 32'd268468224;
      1077: inst = 32'd201343213;
      1078: inst = 32'd203484854;
      1079: inst = 32'd136314880;
      1080: inst = 32'd268468224;
      1081: inst = 32'd201343214;
      1082: inst = 32'd203484854;
      1083: inst = 32'd136314880;
      1084: inst = 32'd268468224;
      1085: inst = 32'd201343215;
      1086: inst = 32'd203484854;
      1087: inst = 32'd136314880;
      1088: inst = 32'd268468224;
      1089: inst = 32'd201343216;
      1090: inst = 32'd203484854;
      1091: inst = 32'd136314880;
      1092: inst = 32'd268468224;
      1093: inst = 32'd201343217;
      1094: inst = 32'd203484854;
      1095: inst = 32'd136314880;
      1096: inst = 32'd268468224;
      1097: inst = 32'd201343218;
      1098: inst = 32'd203484854;
      1099: inst = 32'd136314880;
      1100: inst = 32'd268468224;
      1101: inst = 32'd201343219;
      1102: inst = 32'd203484854;
      1103: inst = 32'd136314880;
      1104: inst = 32'd268468224;
      1105: inst = 32'd201343220;
      1106: inst = 32'd203484854;
      1107: inst = 32'd136314880;
      1108: inst = 32'd268468224;
      1109: inst = 32'd201343221;
      1110: inst = 32'd203484854;
      1111: inst = 32'd136314880;
      1112: inst = 32'd268468224;
      1113: inst = 32'd201343222;
      1114: inst = 32'd203484854;
      1115: inst = 32'd136314880;
      1116: inst = 32'd268468224;
      1117: inst = 32'd201343223;
      1118: inst = 32'd203484854;
      1119: inst = 32'd136314880;
      1120: inst = 32'd268468224;
      1121: inst = 32'd201343224;
      1122: inst = 32'd203484854;
      1123: inst = 32'd136314880;
      1124: inst = 32'd268468224;
      1125: inst = 32'd201343225;
      1126: inst = 32'd203484854;
      1127: inst = 32'd136314880;
      1128: inst = 32'd268468224;
      1129: inst = 32'd201343226;
      1130: inst = 32'd203484854;
      1131: inst = 32'd136314880;
      1132: inst = 32'd268468224;
      1133: inst = 32'd201343227;
      1134: inst = 32'd203484854;
      1135: inst = 32'd136314880;
      1136: inst = 32'd268468224;
      1137: inst = 32'd201343228;
      1138: inst = 32'd203484854;
      1139: inst = 32'd136314880;
      1140: inst = 32'd268468224;
      1141: inst = 32'd201343229;
      1142: inst = 32'd203484854;
      1143: inst = 32'd136314880;
      1144: inst = 32'd268468224;
      1145: inst = 32'd201343230;
      1146: inst = 32'd203484854;
      1147: inst = 32'd136314880;
      1148: inst = 32'd268468224;
      1149: inst = 32'd201343231;
      1150: inst = 32'd203484854;
      1151: inst = 32'd136314880;
      1152: inst = 32'd268468224;
      1153: inst = 32'd201343232;
      1154: inst = 32'd203482839;
      1155: inst = 32'd136314880;
      1156: inst = 32'd268468224;
      1157: inst = 32'd201343233;
      1158: inst = 32'd203484855;
      1159: inst = 32'd136314880;
      1160: inst = 32'd268468224;
      1161: inst = 32'd201343234;
      1162: inst = 32'd203484854;
      1163: inst = 32'd136314880;
      1164: inst = 32'd268468224;
      1165: inst = 32'd201343235;
      1166: inst = 32'd203484854;
      1167: inst = 32'd136314880;
      1168: inst = 32'd268468224;
      1169: inst = 32'd201343236;
      1170: inst = 32'd203486902;
      1171: inst = 32'd136314880;
      1172: inst = 32'd268468224;
      1173: inst = 32'd201343237;
      1174: inst = 32'd203486902;
      1175: inst = 32'd136314880;
      1176: inst = 32'd268468224;
      1177: inst = 32'd201343238;
      1178: inst = 32'd203484854;
      1179: inst = 32'd136314880;
      1180: inst = 32'd268468224;
      1181: inst = 32'd201343239;
      1182: inst = 32'd203484855;
      1183: inst = 32'd136314880;
      1184: inst = 32'd268468224;
      1185: inst = 32'd201343240;
      1186: inst = 32'd203484855;
      1187: inst = 32'd136314880;
      1188: inst = 32'd268468224;
      1189: inst = 32'd201343241;
      1190: inst = 32'd203482808;
      1191: inst = 32'd136314880;
      1192: inst = 32'd268468224;
      1193: inst = 32'd201343242;
      1194: inst = 32'd203482840;
      1195: inst = 32'd136314880;
      1196: inst = 32'd268468224;
      1197: inst = 32'd201343243;
      1198: inst = 32'd203463856;
      1199: inst = 32'd136314880;
      1200: inst = 32'd268468224;
      1201: inst = 32'd201343244;
      1202: inst = 32'd203482808;
      1203: inst = 32'd136314880;
      1204: inst = 32'd268468224;
      1205: inst = 32'd201343245;
      1206: inst = 32'd203482807;
      1207: inst = 32'd136314880;
      1208: inst = 32'd268468224;
      1209: inst = 32'd201343246;
      1210: inst = 32'd203484855;
      1211: inst = 32'd136314880;
      1212: inst = 32'd268468224;
      1213: inst = 32'd201343247;
      1214: inst = 32'd203484855;
      1215: inst = 32'd136314880;
      1216: inst = 32'd268468224;
      1217: inst = 32'd201343248;
      1218: inst = 32'd203484854;
      1219: inst = 32'd136314880;
      1220: inst = 32'd268468224;
      1221: inst = 32'd201343249;
      1222: inst = 32'd203484854;
      1223: inst = 32'd136314880;
      1224: inst = 32'd268468224;
      1225: inst = 32'd201343250;
      1226: inst = 32'd203484854;
      1227: inst = 32'd136314880;
      1228: inst = 32'd268468224;
      1229: inst = 32'd201343251;
      1230: inst = 32'd203484854;
      1231: inst = 32'd136314880;
      1232: inst = 32'd268468224;
      1233: inst = 32'd201343252;
      1234: inst = 32'd203484855;
      1235: inst = 32'd136314880;
      1236: inst = 32'd268468224;
      1237: inst = 32'd201343253;
      1238: inst = 32'd203484855;
      1239: inst = 32'd136314880;
      1240: inst = 32'd268468224;
      1241: inst = 32'd201343254;
      1242: inst = 32'd203484854;
      1243: inst = 32'd136314880;
      1244: inst = 32'd268468224;
      1245: inst = 32'd201343255;
      1246: inst = 32'd203484854;
      1247: inst = 32'd136314880;
      1248: inst = 32'd268468224;
      1249: inst = 32'd201343256;
      1250: inst = 32'd203484822;
      1251: inst = 32'd136314880;
      1252: inst = 32'd268468224;
      1253: inst = 32'd201343257;
      1254: inst = 32'd203484854;
      1255: inst = 32'd136314880;
      1256: inst = 32'd268468224;
      1257: inst = 32'd201343258;
      1258: inst = 32'd203484854;
      1259: inst = 32'd136314880;
      1260: inst = 32'd268468224;
      1261: inst = 32'd201343259;
      1262: inst = 32'd203486967;
      1263: inst = 32'd136314880;
      1264: inst = 32'd268468224;
      1265: inst = 32'd201343260;
      1266: inst = 32'd203484887;
      1267: inst = 32'd136314880;
      1268: inst = 32'd268468224;
      1269: inst = 32'd201343261;
      1270: inst = 32'd203484920;
      1271: inst = 32'd136314880;
      1272: inst = 32'd268468224;
      1273: inst = 32'd201343262;
      1274: inst = 32'd203482807;
      1275: inst = 32'd136314880;
      1276: inst = 32'd268468224;
      1277: inst = 32'd201343263;
      1278: inst = 32'd203482807;
      1279: inst = 32'd136314880;
      1280: inst = 32'd268468224;
      1281: inst = 32'd201343264;
      1282: inst = 32'd203484917;
      1283: inst = 32'd136314880;
      1284: inst = 32'd268468224;
      1285: inst = 32'd201343265;
      1286: inst = 32'd203484917;
      1287: inst = 32'd136314880;
      1288: inst = 32'd268468224;
      1289: inst = 32'd201343266;
      1290: inst = 32'd203484917;
      1291: inst = 32'd136314880;
      1292: inst = 32'd268468224;
      1293: inst = 32'd201343267;
      1294: inst = 32'd203484917;
      1295: inst = 32'd136314880;
      1296: inst = 32'd268468224;
      1297: inst = 32'd201343268;
      1298: inst = 32'd203484917;
      1299: inst = 32'd136314880;
      1300: inst = 32'd268468224;
      1301: inst = 32'd201343269;
      1302: inst = 32'd203484917;
      1303: inst = 32'd136314880;
      1304: inst = 32'd268468224;
      1305: inst = 32'd201343270;
      1306: inst = 32'd203484917;
      1307: inst = 32'd136314880;
      1308: inst = 32'd268468224;
      1309: inst = 32'd201343271;
      1310: inst = 32'd203484917;
      1311: inst = 32'd136314880;
      1312: inst = 32'd268468224;
      1313: inst = 32'd201343272;
      1314: inst = 32'd203484917;
      1315: inst = 32'd136314880;
      1316: inst = 32'd268468224;
      1317: inst = 32'd201343273;
      1318: inst = 32'd203484917;
      1319: inst = 32'd136314880;
      1320: inst = 32'd268468224;
      1321: inst = 32'd201343274;
      1322: inst = 32'd203484917;
      1323: inst = 32'd136314880;
      1324: inst = 32'd268468224;
      1325: inst = 32'd201343275;
      1326: inst = 32'd203484917;
      1327: inst = 32'd136314880;
      1328: inst = 32'd268468224;
      1329: inst = 32'd201343276;
      1330: inst = 32'd203484917;
      1331: inst = 32'd136314880;
      1332: inst = 32'd268468224;
      1333: inst = 32'd201343277;
      1334: inst = 32'd203484917;
      1335: inst = 32'd136314880;
      1336: inst = 32'd268468224;
      1337: inst = 32'd201343278;
      1338: inst = 32'd203484917;
      1339: inst = 32'd136314880;
      1340: inst = 32'd268468224;
      1341: inst = 32'd201343279;
      1342: inst = 32'd203484917;
      1343: inst = 32'd136314880;
      1344: inst = 32'd268468224;
      1345: inst = 32'd201343280;
      1346: inst = 32'd203484917;
      1347: inst = 32'd136314880;
      1348: inst = 32'd268468224;
      1349: inst = 32'd201343281;
      1350: inst = 32'd203484917;
      1351: inst = 32'd136314880;
      1352: inst = 32'd268468224;
      1353: inst = 32'd201343282;
      1354: inst = 32'd203484917;
      1355: inst = 32'd136314880;
      1356: inst = 32'd268468224;
      1357: inst = 32'd201343283;
      1358: inst = 32'd203484917;
      1359: inst = 32'd136314880;
      1360: inst = 32'd268468224;
      1361: inst = 32'd201343284;
      1362: inst = 32'd203484917;
      1363: inst = 32'd136314880;
      1364: inst = 32'd268468224;
      1365: inst = 32'd201343285;
      1366: inst = 32'd203484917;
      1367: inst = 32'd136314880;
      1368: inst = 32'd268468224;
      1369: inst = 32'd201343286;
      1370: inst = 32'd203484917;
      1371: inst = 32'd136314880;
      1372: inst = 32'd268468224;
      1373: inst = 32'd201343287;
      1374: inst = 32'd203484917;
      1375: inst = 32'd136314880;
      1376: inst = 32'd268468224;
      1377: inst = 32'd201343288;
      1378: inst = 32'd203484917;
      1379: inst = 32'd136314880;
      1380: inst = 32'd268468224;
      1381: inst = 32'd201343289;
      1382: inst = 32'd203484917;
      1383: inst = 32'd136314880;
      1384: inst = 32'd268468224;
      1385: inst = 32'd201343290;
      1386: inst = 32'd203484917;
      1387: inst = 32'd136314880;
      1388: inst = 32'd268468224;
      1389: inst = 32'd201343291;
      1390: inst = 32'd203484917;
      1391: inst = 32'd136314880;
      1392: inst = 32'd268468224;
      1393: inst = 32'd201343292;
      1394: inst = 32'd203484917;
      1395: inst = 32'd136314880;
      1396: inst = 32'd268468224;
      1397: inst = 32'd201343293;
      1398: inst = 32'd203484917;
      1399: inst = 32'd136314880;
      1400: inst = 32'd268468224;
      1401: inst = 32'd201343294;
      1402: inst = 32'd203484917;
      1403: inst = 32'd136314880;
      1404: inst = 32'd268468224;
      1405: inst = 32'd201343295;
      1406: inst = 32'd203484917;
      1407: inst = 32'd136314880;
      1408: inst = 32'd268468224;
      1409: inst = 32'd201343296;
      1410: inst = 32'd203482807;
      1411: inst = 32'd136314880;
      1412: inst = 32'd268468224;
      1413: inst = 32'd201343297;
      1414: inst = 32'd203482807;
      1415: inst = 32'd136314880;
      1416: inst = 32'd268468224;
      1417: inst = 32'd201343298;
      1418: inst = 32'd203484920;
      1419: inst = 32'd136314880;
      1420: inst = 32'd268468224;
      1421: inst = 32'd201343299;
      1422: inst = 32'd203484855;
      1423: inst = 32'd136314880;
      1424: inst = 32'd268468224;
      1425: inst = 32'd201343300;
      1426: inst = 32'd203486935;
      1427: inst = 32'd136314880;
      1428: inst = 32'd268468224;
      1429: inst = 32'd201343301;
      1430: inst = 32'd203484822;
      1431: inst = 32'd136314880;
      1432: inst = 32'd268468224;
      1433: inst = 32'd201343302;
      1434: inst = 32'd203486902;
      1435: inst = 32'd136314880;
      1436: inst = 32'd268468224;
      1437: inst = 32'd201343303;
      1438: inst = 32'd203484822;
      1439: inst = 32'd136314880;
      1440: inst = 32'd268468224;
      1441: inst = 32'd201343304;
      1442: inst = 32'd203484854;
      1443: inst = 32'd136314880;
      1444: inst = 32'd268468224;
      1445: inst = 32'd201343305;
      1446: inst = 32'd203484854;
      1447: inst = 32'd136314880;
      1448: inst = 32'd268468224;
      1449: inst = 32'd201343306;
      1450: inst = 32'd203484855;
      1451: inst = 32'd136314880;
      1452: inst = 32'd268468224;
      1453: inst = 32'd201343307;
      1454: inst = 32'd203484855;
      1455: inst = 32'd136314880;
      1456: inst = 32'd268468224;
      1457: inst = 32'd201343308;
      1458: inst = 32'd203484854;
      1459: inst = 32'd136314880;
      1460: inst = 32'd268468224;
      1461: inst = 32'd201343309;
      1462: inst = 32'd203484854;
      1463: inst = 32'd136314880;
      1464: inst = 32'd268468224;
      1465: inst = 32'd201343310;
      1466: inst = 32'd203484854;
      1467: inst = 32'd136314880;
      1468: inst = 32'd268468224;
      1469: inst = 32'd201343311;
      1470: inst = 32'd203484854;
      1471: inst = 32'd136314880;
      1472: inst = 32'd268468224;
      1473: inst = 32'd201343312;
      1474: inst = 32'd203484854;
      1475: inst = 32'd136314880;
      1476: inst = 32'd268468224;
      1477: inst = 32'd201343313;
      1478: inst = 32'd203484854;
      1479: inst = 32'd136314880;
      1480: inst = 32'd268468224;
      1481: inst = 32'd201343314;
      1482: inst = 32'd203484854;
      1483: inst = 32'd136314880;
      1484: inst = 32'd268468224;
      1485: inst = 32'd201343315;
      1486: inst = 32'd203484854;
      1487: inst = 32'd136314880;
      1488: inst = 32'd268468224;
      1489: inst = 32'd201343316;
      1490: inst = 32'd203484854;
      1491: inst = 32'd136314880;
      1492: inst = 32'd268468224;
      1493: inst = 32'd201343317;
      1494: inst = 32'd203484854;
      1495: inst = 32'd136314880;
      1496: inst = 32'd268468224;
      1497: inst = 32'd201343318;
      1498: inst = 32'd203484854;
      1499: inst = 32'd136314880;
      1500: inst = 32'd268468224;
      1501: inst = 32'd201343319;
      1502: inst = 32'd203484854;
      1503: inst = 32'd136314880;
      1504: inst = 32'd268468224;
      1505: inst = 32'd201343320;
      1506: inst = 32'd203484854;
      1507: inst = 32'd136314880;
      1508: inst = 32'd268468224;
      1509: inst = 32'd201343321;
      1510: inst = 32'd203484854;
      1511: inst = 32'd136314880;
      1512: inst = 32'd268468224;
      1513: inst = 32'd201343322;
      1514: inst = 32'd203484854;
      1515: inst = 32'd136314880;
      1516: inst = 32'd268468224;
      1517: inst = 32'd201343323;
      1518: inst = 32'd203484854;
      1519: inst = 32'd136314880;
      1520: inst = 32'd268468224;
      1521: inst = 32'd201343324;
      1522: inst = 32'd203484854;
      1523: inst = 32'd136314880;
      1524: inst = 32'd268468224;
      1525: inst = 32'd201343325;
      1526: inst = 32'd203484854;
      1527: inst = 32'd136314880;
      1528: inst = 32'd268468224;
      1529: inst = 32'd201343326;
      1530: inst = 32'd203484854;
      1531: inst = 32'd136314880;
      1532: inst = 32'd268468224;
      1533: inst = 32'd201343327;
      1534: inst = 32'd203484854;
      1535: inst = 32'd136314880;
      1536: inst = 32'd268468224;
      1537: inst = 32'd201343328;
      1538: inst = 32'd203482839;
      1539: inst = 32'd136314880;
      1540: inst = 32'd268468224;
      1541: inst = 32'd201343329;
      1542: inst = 32'd203482839;
      1543: inst = 32'd136314880;
      1544: inst = 32'd268468224;
      1545: inst = 32'd201343330;
      1546: inst = 32'd203484854;
      1547: inst = 32'd136314880;
      1548: inst = 32'd268468224;
      1549: inst = 32'd201343331;
      1550: inst = 32'd203484854;
      1551: inst = 32'd136314880;
      1552: inst = 32'd268468224;
      1553: inst = 32'd201343332;
      1554: inst = 32'd203486870;
      1555: inst = 32'd136314880;
      1556: inst = 32'd268468224;
      1557: inst = 32'd201343333;
      1558: inst = 32'd203486870;
      1559: inst = 32'd136314880;
      1560: inst = 32'd268468224;
      1561: inst = 32'd201343334;
      1562: inst = 32'd203486870;
      1563: inst = 32'd136314880;
      1564: inst = 32'd268468224;
      1565: inst = 32'd201343335;
      1566: inst = 32'd203486871;
      1567: inst = 32'd136314880;
      1568: inst = 32'd268468224;
      1569: inst = 32'd201343336;
      1570: inst = 32'd203484855;
      1571: inst = 32'd136314880;
      1572: inst = 32'd268468224;
      1573: inst = 32'd201343337;
      1574: inst = 32'd203484824;
      1575: inst = 32'd136314880;
      1576: inst = 32'd268468224;
      1577: inst = 32'd201343338;
      1578: inst = 32'd203484856;
      1579: inst = 32'd136314880;
      1580: inst = 32'd268468224;
      1581: inst = 32'd201343339;
      1582: inst = 32'd203467888;
      1583: inst = 32'd136314880;
      1584: inst = 32'd268468224;
      1585: inst = 32'd201343340;
      1586: inst = 32'd203486872;
      1587: inst = 32'd136314880;
      1588: inst = 32'd268468224;
      1589: inst = 32'd201343341;
      1590: inst = 32'd203486840;
      1591: inst = 32'd136314880;
      1592: inst = 32'd268468224;
      1593: inst = 32'd201343342;
      1594: inst = 32'd203488855;
      1595: inst = 32'd136314880;
      1596: inst = 32'd268468224;
      1597: inst = 32'd201343343;
      1598: inst = 32'd203488888;
      1599: inst = 32'd136314880;
      1600: inst = 32'd268468224;
      1601: inst = 32'd201343344;
      1602: inst = 32'd203486902;
      1603: inst = 32'd136314880;
      1604: inst = 32'd268468224;
      1605: inst = 32'd201343345;
      1606: inst = 32'd203484854;
      1607: inst = 32'd136314880;
      1608: inst = 32'd268468224;
      1609: inst = 32'd201343346;
      1610: inst = 32'd203484854;
      1611: inst = 32'd136314880;
      1612: inst = 32'd268468224;
      1613: inst = 32'd201343347;
      1614: inst = 32'd203484854;
      1615: inst = 32'd136314880;
      1616: inst = 32'd268468224;
      1617: inst = 32'd201343348;
      1618: inst = 32'd203484854;
      1619: inst = 32'd136314880;
      1620: inst = 32'd268468224;
      1621: inst = 32'd201343349;
      1622: inst = 32'd203484854;
      1623: inst = 32'd136314880;
      1624: inst = 32'd268468224;
      1625: inst = 32'd201343350;
      1626: inst = 32'd203484854;
      1627: inst = 32'd136314880;
      1628: inst = 32'd268468224;
      1629: inst = 32'd201343351;
      1630: inst = 32'd203484854;
      1631: inst = 32'd136314880;
      1632: inst = 32'd268468224;
      1633: inst = 32'd201343352;
      1634: inst = 32'd203484854;
      1635: inst = 32'd136314880;
      1636: inst = 32'd268468224;
      1637: inst = 32'd201343353;
      1638: inst = 32'd203486935;
      1639: inst = 32'd136314880;
      1640: inst = 32'd268468224;
      1641: inst = 32'd201343354;
      1642: inst = 32'd203482742;
      1643: inst = 32'd136314880;
      1644: inst = 32'd268468224;
      1645: inst = 32'd201343355;
      1646: inst = 32'd203484854;
      1647: inst = 32'd136314880;
      1648: inst = 32'd268468224;
      1649: inst = 32'd201343356;
      1650: inst = 32'd203482807;
      1651: inst = 32'd136314880;
      1652: inst = 32'd268468224;
      1653: inst = 32'd201343357;
      1654: inst = 32'd203484888;
      1655: inst = 32'd136314880;
      1656: inst = 32'd268468224;
      1657: inst = 32'd201343358;
      1658: inst = 32'd203480728;
      1659: inst = 32'd136314880;
      1660: inst = 32'd268468224;
      1661: inst = 32'd201343359;
      1662: inst = 32'd203482840;
      1663: inst = 32'd136314880;
      1664: inst = 32'd268468224;
      1665: inst = 32'd201343360;
      1666: inst = 32'd203482839;
      1667: inst = 32'd136314880;
      1668: inst = 32'd268468224;
      1669: inst = 32'd201343361;
      1670: inst = 32'd203482839;
      1671: inst = 32'd136314880;
      1672: inst = 32'd268468224;
      1673: inst = 32'd201343362;
      1674: inst = 32'd203482839;
      1675: inst = 32'd136314880;
      1676: inst = 32'd268468224;
      1677: inst = 32'd201343363;
      1678: inst = 32'd203482839;
      1679: inst = 32'd136314880;
      1680: inst = 32'd268468224;
      1681: inst = 32'd201343364;
      1682: inst = 32'd203482839;
      1683: inst = 32'd136314880;
      1684: inst = 32'd268468224;
      1685: inst = 32'd201343365;
      1686: inst = 32'd203482839;
      1687: inst = 32'd136314880;
      1688: inst = 32'd268468224;
      1689: inst = 32'd201343366;
      1690: inst = 32'd203482839;
      1691: inst = 32'd136314880;
      1692: inst = 32'd268468224;
      1693: inst = 32'd201343367;
      1694: inst = 32'd203482839;
      1695: inst = 32'd136314880;
      1696: inst = 32'd268468224;
      1697: inst = 32'd201343368;
      1698: inst = 32'd203482839;
      1699: inst = 32'd136314880;
      1700: inst = 32'd268468224;
      1701: inst = 32'd201343369;
      1702: inst = 32'd203482839;
      1703: inst = 32'd136314880;
      1704: inst = 32'd268468224;
      1705: inst = 32'd201343370;
      1706: inst = 32'd203482839;
      1707: inst = 32'd136314880;
      1708: inst = 32'd268468224;
      1709: inst = 32'd201343371;
      1710: inst = 32'd203482839;
      1711: inst = 32'd136314880;
      1712: inst = 32'd268468224;
      1713: inst = 32'd201343372;
      1714: inst = 32'd203482839;
      1715: inst = 32'd136314880;
      1716: inst = 32'd268468224;
      1717: inst = 32'd201343373;
      1718: inst = 32'd203482839;
      1719: inst = 32'd136314880;
      1720: inst = 32'd268468224;
      1721: inst = 32'd201343374;
      1722: inst = 32'd203482839;
      1723: inst = 32'd136314880;
      1724: inst = 32'd268468224;
      1725: inst = 32'd201343375;
      1726: inst = 32'd203482839;
      1727: inst = 32'd136314880;
      1728: inst = 32'd268468224;
      1729: inst = 32'd201343376;
      1730: inst = 32'd203482839;
      1731: inst = 32'd136314880;
      1732: inst = 32'd268468224;
      1733: inst = 32'd201343377;
      1734: inst = 32'd203482839;
      1735: inst = 32'd136314880;
      1736: inst = 32'd268468224;
      1737: inst = 32'd201343378;
      1738: inst = 32'd203482839;
      1739: inst = 32'd136314880;
      1740: inst = 32'd268468224;
      1741: inst = 32'd201343379;
      1742: inst = 32'd203482839;
      1743: inst = 32'd136314880;
      1744: inst = 32'd268468224;
      1745: inst = 32'd201343380;
      1746: inst = 32'd203482839;
      1747: inst = 32'd136314880;
      1748: inst = 32'd268468224;
      1749: inst = 32'd201343381;
      1750: inst = 32'd203482839;
      1751: inst = 32'd136314880;
      1752: inst = 32'd268468224;
      1753: inst = 32'd201343382;
      1754: inst = 32'd203482839;
      1755: inst = 32'd136314880;
      1756: inst = 32'd268468224;
      1757: inst = 32'd201343383;
      1758: inst = 32'd203482839;
      1759: inst = 32'd136314880;
      1760: inst = 32'd268468224;
      1761: inst = 32'd201343384;
      1762: inst = 32'd203482839;
      1763: inst = 32'd136314880;
      1764: inst = 32'd268468224;
      1765: inst = 32'd201343385;
      1766: inst = 32'd203482839;
      1767: inst = 32'd136314880;
      1768: inst = 32'd268468224;
      1769: inst = 32'd201343386;
      1770: inst = 32'd203482839;
      1771: inst = 32'd136314880;
      1772: inst = 32'd268468224;
      1773: inst = 32'd201343387;
      1774: inst = 32'd203482839;
      1775: inst = 32'd136314880;
      1776: inst = 32'd268468224;
      1777: inst = 32'd201343388;
      1778: inst = 32'd203482839;
      1779: inst = 32'd136314880;
      1780: inst = 32'd268468224;
      1781: inst = 32'd201343389;
      1782: inst = 32'd203482839;
      1783: inst = 32'd136314880;
      1784: inst = 32'd268468224;
      1785: inst = 32'd201343390;
      1786: inst = 32'd203482839;
      1787: inst = 32'd136314880;
      1788: inst = 32'd268468224;
      1789: inst = 32'd201343391;
      1790: inst = 32'd203482839;
      1791: inst = 32'd136314880;
      1792: inst = 32'd268468224;
      1793: inst = 32'd201343392;
      1794: inst = 32'd203482840;
      1795: inst = 32'd136314880;
      1796: inst = 32'd268468224;
      1797: inst = 32'd201343393;
      1798: inst = 32'd203480728;
      1799: inst = 32'd136314880;
      1800: inst = 32'd268468224;
      1801: inst = 32'd201343394;
      1802: inst = 32'd203484888;
      1803: inst = 32'd136314880;
      1804: inst = 32'd268468224;
      1805: inst = 32'd201343395;
      1806: inst = 32'd203482807;
      1807: inst = 32'd136314880;
      1808: inst = 32'd268468224;
      1809: inst = 32'd201343396;
      1810: inst = 32'd203484854;
      1811: inst = 32'd136314880;
      1812: inst = 32'd268468224;
      1813: inst = 32'd201343397;
      1814: inst = 32'd203482742;
      1815: inst = 32'd136314880;
      1816: inst = 32'd268468224;
      1817: inst = 32'd201343398;
      1818: inst = 32'd203486935;
      1819: inst = 32'd136314880;
      1820: inst = 32'd268468224;
      1821: inst = 32'd201343399;
      1822: inst = 32'd203484854;
      1823: inst = 32'd136314880;
      1824: inst = 32'd268468224;
      1825: inst = 32'd201343400;
      1826: inst = 32'd203484854;
      1827: inst = 32'd136314880;
      1828: inst = 32'd268468224;
      1829: inst = 32'd201343401;
      1830: inst = 32'd203484854;
      1831: inst = 32'd136314880;
      1832: inst = 32'd268468224;
      1833: inst = 32'd201343402;
      1834: inst = 32'd203484854;
      1835: inst = 32'd136314880;
      1836: inst = 32'd268468224;
      1837: inst = 32'd201343403;
      1838: inst = 32'd203484854;
      1839: inst = 32'd136314880;
      1840: inst = 32'd268468224;
      1841: inst = 32'd201343404;
      1842: inst = 32'd203484854;
      1843: inst = 32'd136314880;
      1844: inst = 32'd268468224;
      1845: inst = 32'd201343405;
      1846: inst = 32'd203484854;
      1847: inst = 32'd136314880;
      1848: inst = 32'd268468224;
      1849: inst = 32'd201343406;
      1850: inst = 32'd203484854;
      1851: inst = 32'd136314880;
      1852: inst = 32'd268468224;
      1853: inst = 32'd201343407;
      1854: inst = 32'd203484854;
      1855: inst = 32'd136314880;
      1856: inst = 32'd268468224;
      1857: inst = 32'd201343408;
      1858: inst = 32'd203484854;
      1859: inst = 32'd136314880;
      1860: inst = 32'd268468224;
      1861: inst = 32'd201343409;
      1862: inst = 32'd203484854;
      1863: inst = 32'd136314880;
      1864: inst = 32'd268468224;
      1865: inst = 32'd201343410;
      1866: inst = 32'd203484854;
      1867: inst = 32'd136314880;
      1868: inst = 32'd268468224;
      1869: inst = 32'd201343411;
      1870: inst = 32'd203484854;
      1871: inst = 32'd136314880;
      1872: inst = 32'd268468224;
      1873: inst = 32'd201343412;
      1874: inst = 32'd203484854;
      1875: inst = 32'd136314880;
      1876: inst = 32'd268468224;
      1877: inst = 32'd201343413;
      1878: inst = 32'd203484854;
      1879: inst = 32'd136314880;
      1880: inst = 32'd268468224;
      1881: inst = 32'd201343414;
      1882: inst = 32'd203484854;
      1883: inst = 32'd136314880;
      1884: inst = 32'd268468224;
      1885: inst = 32'd201343415;
      1886: inst = 32'd203484854;
      1887: inst = 32'd136314880;
      1888: inst = 32'd268468224;
      1889: inst = 32'd201343416;
      1890: inst = 32'd203484854;
      1891: inst = 32'd136314880;
      1892: inst = 32'd268468224;
      1893: inst = 32'd201343417;
      1894: inst = 32'd203484854;
      1895: inst = 32'd136314880;
      1896: inst = 32'd268468224;
      1897: inst = 32'd201343418;
      1898: inst = 32'd203484854;
      1899: inst = 32'd136314880;
      1900: inst = 32'd268468224;
      1901: inst = 32'd201343419;
      1902: inst = 32'd203484854;
      1903: inst = 32'd136314880;
      1904: inst = 32'd268468224;
      1905: inst = 32'd201343420;
      1906: inst = 32'd203484854;
      1907: inst = 32'd136314880;
      1908: inst = 32'd268468224;
      1909: inst = 32'd201343421;
      1910: inst = 32'd203484854;
      1911: inst = 32'd136314880;
      1912: inst = 32'd268468224;
      1913: inst = 32'd201343422;
      1914: inst = 32'd203484854;
      1915: inst = 32'd136314880;
      1916: inst = 32'd268468224;
      1917: inst = 32'd201343423;
      1918: inst = 32'd203484854;
      1919: inst = 32'd136314880;
      1920: inst = 32'd268468224;
      1921: inst = 32'd201343424;
      1922: inst = 32'd203482839;
      1923: inst = 32'd136314880;
      1924: inst = 32'd268468224;
      1925: inst = 32'd201343425;
      1926: inst = 32'd203482839;
      1927: inst = 32'd136314880;
      1928: inst = 32'd268468224;
      1929: inst = 32'd201343426;
      1930: inst = 32'd203484854;
      1931: inst = 32'd136314880;
      1932: inst = 32'd268468224;
      1933: inst = 32'd201343427;
      1934: inst = 32'd203486902;
      1935: inst = 32'd136314880;
      1936: inst = 32'd268468224;
      1937: inst = 32'd201343428;
      1938: inst = 32'd203486870;
      1939: inst = 32'd136314880;
      1940: inst = 32'd268468224;
      1941: inst = 32'd201343429;
      1942: inst = 32'd203488918;
      1943: inst = 32'd136314880;
      1944: inst = 32'd268468224;
      1945: inst = 32'd201343430;
      1946: inst = 32'd203486870;
      1947: inst = 32'd136314880;
      1948: inst = 32'd268468224;
      1949: inst = 32'd201343431;
      1950: inst = 32'd203486871;
      1951: inst = 32'd136314880;
      1952: inst = 32'd268468224;
      1953: inst = 32'd201343432;
      1954: inst = 32'd203486903;
      1955: inst = 32'd136314880;
      1956: inst = 32'd268468224;
      1957: inst = 32'd201343433;
      1958: inst = 32'd203484823;
      1959: inst = 32'd136314880;
      1960: inst = 32'd268468224;
      1961: inst = 32'd201343434;
      1962: inst = 32'd203484856;
      1963: inst = 32'd136314880;
      1964: inst = 32'd268468224;
      1965: inst = 32'd201343435;
      1966: inst = 32'd203467888;
      1967: inst = 32'd136314880;
      1968: inst = 32'd268468224;
      1969: inst = 32'd201343436;
      1970: inst = 32'd203486872;
      1971: inst = 32'd136314880;
      1972: inst = 32'd268468224;
      1973: inst = 32'd201343437;
      1974: inst = 32'd203488888;
      1975: inst = 32'd136314880;
      1976: inst = 32'd268468224;
      1977: inst = 32'd201343438;
      1978: inst = 32'd203488855;
      1979: inst = 32'd136314880;
      1980: inst = 32'd268468224;
      1981: inst = 32'd201343439;
      1982: inst = 32'd203488855;
      1983: inst = 32'd136314880;
      1984: inst = 32'd268468224;
      1985: inst = 32'd201343440;
      1986: inst = 32'd203486902;
      1987: inst = 32'd136314880;
      1988: inst = 32'd268468224;
      1989: inst = 32'd201343441;
      1990: inst = 32'd203484854;
      1991: inst = 32'd136314880;
      1992: inst = 32'd268468224;
      1993: inst = 32'd201343442;
      1994: inst = 32'd203484854;
      1995: inst = 32'd136314880;
      1996: inst = 32'd268468224;
      1997: inst = 32'd201343443;
      1998: inst = 32'd203484854;
      1999: inst = 32'd136314880;
      2000: inst = 32'd268468224;
      2001: inst = 32'd201343444;
      2002: inst = 32'd203484854;
      2003: inst = 32'd136314880;
      2004: inst = 32'd268468224;
      2005: inst = 32'd201343445;
      2006: inst = 32'd203484854;
      2007: inst = 32'd136314880;
      2008: inst = 32'd268468224;
      2009: inst = 32'd201343446;
      2010: inst = 32'd203484854;
      2011: inst = 32'd136314880;
      2012: inst = 32'd268468224;
      2013: inst = 32'd201343447;
      2014: inst = 32'd203484854;
      2015: inst = 32'd136314880;
      2016: inst = 32'd268468224;
      2017: inst = 32'd201343448;
      2018: inst = 32'd203484887;
      2019: inst = 32'd136314880;
      2020: inst = 32'd268468224;
      2021: inst = 32'd201343449;
      2022: inst = 32'd203482774;
      2023: inst = 32'd136314880;
      2024: inst = 32'd268468224;
      2025: inst = 32'd201343450;
      2026: inst = 32'd203476435;
      2027: inst = 32'd136314880;
      2028: inst = 32'd268468224;
      2029: inst = 32'd201343451;
      2030: inst = 32'd203474290;
      2031: inst = 32'd136314880;
      2032: inst = 32'd268468224;
      2033: inst = 32'd201343452;
      2034: inst = 32'd203472275;
      2035: inst = 32'd136314880;
      2036: inst = 32'd268468224;
      2037: inst = 32'd201343453;
      2038: inst = 32'd203472276;
      2039: inst = 32'd136314880;
      2040: inst = 32'd268468224;
      2041: inst = 32'd201343454;
      2042: inst = 32'd203470196;
      2043: inst = 32'd136314880;
      2044: inst = 32'd268468224;
      2045: inst = 32'd201343455;
      2046: inst = 32'd203472277;
      2047: inst = 32'd136314880;
      2048: inst = 32'd268468224;
      2049: inst = 32'd201343456;
      2050: inst = 32'd203472277;
      2051: inst = 32'd136314880;
      2052: inst = 32'd268468224;
      2053: inst = 32'd201343457;
      2054: inst = 32'd203472277;
      2055: inst = 32'd136314880;
      2056: inst = 32'd268468224;
      2057: inst = 32'd201343458;
      2058: inst = 32'd203472277;
      2059: inst = 32'd136314880;
      2060: inst = 32'd268468224;
      2061: inst = 32'd201343459;
      2062: inst = 32'd203472277;
      2063: inst = 32'd136314880;
      2064: inst = 32'd268468224;
      2065: inst = 32'd201343460;
      2066: inst = 32'd203472277;
      2067: inst = 32'd136314880;
      2068: inst = 32'd268468224;
      2069: inst = 32'd201343461;
      2070: inst = 32'd203472277;
      2071: inst = 32'd136314880;
      2072: inst = 32'd268468224;
      2073: inst = 32'd201343462;
      2074: inst = 32'd203472277;
      2075: inst = 32'd136314880;
      2076: inst = 32'd268468224;
      2077: inst = 32'd201343463;
      2078: inst = 32'd203472277;
      2079: inst = 32'd136314880;
      2080: inst = 32'd268468224;
      2081: inst = 32'd201343464;
      2082: inst = 32'd203472277;
      2083: inst = 32'd136314880;
      2084: inst = 32'd268468224;
      2085: inst = 32'd201343465;
      2086: inst = 32'd203472277;
      2087: inst = 32'd136314880;
      2088: inst = 32'd268468224;
      2089: inst = 32'd201343466;
      2090: inst = 32'd203472277;
      2091: inst = 32'd136314880;
      2092: inst = 32'd268468224;
      2093: inst = 32'd201343467;
      2094: inst = 32'd203472277;
      2095: inst = 32'd136314880;
      2096: inst = 32'd268468224;
      2097: inst = 32'd201343468;
      2098: inst = 32'd203472277;
      2099: inst = 32'd136314880;
      2100: inst = 32'd268468224;
      2101: inst = 32'd201343469;
      2102: inst = 32'd203472277;
      2103: inst = 32'd136314880;
      2104: inst = 32'd268468224;
      2105: inst = 32'd201343470;
      2106: inst = 32'd203472277;
      2107: inst = 32'd136314880;
      2108: inst = 32'd268468224;
      2109: inst = 32'd201343471;
      2110: inst = 32'd203472277;
      2111: inst = 32'd136314880;
      2112: inst = 32'd268468224;
      2113: inst = 32'd201343472;
      2114: inst = 32'd203472277;
      2115: inst = 32'd136314880;
      2116: inst = 32'd268468224;
      2117: inst = 32'd201343473;
      2118: inst = 32'd203472277;
      2119: inst = 32'd136314880;
      2120: inst = 32'd268468224;
      2121: inst = 32'd201343474;
      2122: inst = 32'd203472277;
      2123: inst = 32'd136314880;
      2124: inst = 32'd268468224;
      2125: inst = 32'd201343475;
      2126: inst = 32'd203472277;
      2127: inst = 32'd136314880;
      2128: inst = 32'd268468224;
      2129: inst = 32'd201343476;
      2130: inst = 32'd203472277;
      2131: inst = 32'd136314880;
      2132: inst = 32'd268468224;
      2133: inst = 32'd201343477;
      2134: inst = 32'd203472277;
      2135: inst = 32'd136314880;
      2136: inst = 32'd268468224;
      2137: inst = 32'd201343478;
      2138: inst = 32'd203472277;
      2139: inst = 32'd136314880;
      2140: inst = 32'd268468224;
      2141: inst = 32'd201343479;
      2142: inst = 32'd203472277;
      2143: inst = 32'd136314880;
      2144: inst = 32'd268468224;
      2145: inst = 32'd201343480;
      2146: inst = 32'd203472277;
      2147: inst = 32'd136314880;
      2148: inst = 32'd268468224;
      2149: inst = 32'd201343481;
      2150: inst = 32'd203472277;
      2151: inst = 32'd136314880;
      2152: inst = 32'd268468224;
      2153: inst = 32'd201343482;
      2154: inst = 32'd203472277;
      2155: inst = 32'd136314880;
      2156: inst = 32'd268468224;
      2157: inst = 32'd201343483;
      2158: inst = 32'd203472277;
      2159: inst = 32'd136314880;
      2160: inst = 32'd268468224;
      2161: inst = 32'd201343484;
      2162: inst = 32'd203472277;
      2163: inst = 32'd136314880;
      2164: inst = 32'd268468224;
      2165: inst = 32'd201343485;
      2166: inst = 32'd203472277;
      2167: inst = 32'd136314880;
      2168: inst = 32'd268468224;
      2169: inst = 32'd201343486;
      2170: inst = 32'd203472277;
      2171: inst = 32'd136314880;
      2172: inst = 32'd268468224;
      2173: inst = 32'd201343487;
      2174: inst = 32'd203472277;
      2175: inst = 32'd136314880;
      2176: inst = 32'd268468224;
      2177: inst = 32'd201343488;
      2178: inst = 32'd203472277;
      2179: inst = 32'd136314880;
      2180: inst = 32'd268468224;
      2181: inst = 32'd201343489;
      2182: inst = 32'd203470196;
      2183: inst = 32'd136314880;
      2184: inst = 32'd268468224;
      2185: inst = 32'd201343490;
      2186: inst = 32'd203472276;
      2187: inst = 32'd136314880;
      2188: inst = 32'd268468224;
      2189: inst = 32'd201343491;
      2190: inst = 32'd203472275;
      2191: inst = 32'd136314880;
      2192: inst = 32'd268468224;
      2193: inst = 32'd201343492;
      2194: inst = 32'd203474290;
      2195: inst = 32'd136314880;
      2196: inst = 32'd268468224;
      2197: inst = 32'd201343493;
      2198: inst = 32'd203476435;
      2199: inst = 32'd136314880;
      2200: inst = 32'd268468224;
      2201: inst = 32'd201343494;
      2202: inst = 32'd203484822;
      2203: inst = 32'd136314880;
      2204: inst = 32'd268468224;
      2205: inst = 32'd201343495;
      2206: inst = 32'd203486935;
      2207: inst = 32'd136314880;
      2208: inst = 32'd268468224;
      2209: inst = 32'd201343496;
      2210: inst = 32'd203484854;
      2211: inst = 32'd136314880;
      2212: inst = 32'd268468224;
      2213: inst = 32'd201343497;
      2214: inst = 32'd203484854;
      2215: inst = 32'd136314880;
      2216: inst = 32'd268468224;
      2217: inst = 32'd201343498;
      2218: inst = 32'd203484854;
      2219: inst = 32'd136314880;
      2220: inst = 32'd268468224;
      2221: inst = 32'd201343499;
      2222: inst = 32'd203484854;
      2223: inst = 32'd136314880;
      2224: inst = 32'd268468224;
      2225: inst = 32'd201343500;
      2226: inst = 32'd203484854;
      2227: inst = 32'd136314880;
      2228: inst = 32'd268468224;
      2229: inst = 32'd201343501;
      2230: inst = 32'd203484854;
      2231: inst = 32'd136314880;
      2232: inst = 32'd268468224;
      2233: inst = 32'd201343502;
      2234: inst = 32'd203484854;
      2235: inst = 32'd136314880;
      2236: inst = 32'd268468224;
      2237: inst = 32'd201343503;
      2238: inst = 32'd203484854;
      2239: inst = 32'd136314880;
      2240: inst = 32'd268468224;
      2241: inst = 32'd201343504;
      2242: inst = 32'd203484854;
      2243: inst = 32'd136314880;
      2244: inst = 32'd268468224;
      2245: inst = 32'd201343505;
      2246: inst = 32'd203484854;
      2247: inst = 32'd136314880;
      2248: inst = 32'd268468224;
      2249: inst = 32'd201343506;
      2250: inst = 32'd203484854;
      2251: inst = 32'd136314880;
      2252: inst = 32'd268468224;
      2253: inst = 32'd201343507;
      2254: inst = 32'd203484854;
      2255: inst = 32'd136314880;
      2256: inst = 32'd268468224;
      2257: inst = 32'd201343508;
      2258: inst = 32'd203484854;
      2259: inst = 32'd136314880;
      2260: inst = 32'd268468224;
      2261: inst = 32'd201343509;
      2262: inst = 32'd203484854;
      2263: inst = 32'd136314880;
      2264: inst = 32'd268468224;
      2265: inst = 32'd201343510;
      2266: inst = 32'd203484854;
      2267: inst = 32'd136314880;
      2268: inst = 32'd268468224;
      2269: inst = 32'd201343511;
      2270: inst = 32'd203484854;
      2271: inst = 32'd136314880;
      2272: inst = 32'd268468224;
      2273: inst = 32'd201343512;
      2274: inst = 32'd203484854;
      2275: inst = 32'd136314880;
      2276: inst = 32'd268468224;
      2277: inst = 32'd201343513;
      2278: inst = 32'd203484854;
      2279: inst = 32'd136314880;
      2280: inst = 32'd268468224;
      2281: inst = 32'd201343514;
      2282: inst = 32'd203484854;
      2283: inst = 32'd136314880;
      2284: inst = 32'd268468224;
      2285: inst = 32'd201343515;
      2286: inst = 32'd203484854;
      2287: inst = 32'd136314880;
      2288: inst = 32'd268468224;
      2289: inst = 32'd201343516;
      2290: inst = 32'd203484854;
      2291: inst = 32'd136314880;
      2292: inst = 32'd268468224;
      2293: inst = 32'd201343517;
      2294: inst = 32'd203484854;
      2295: inst = 32'd136314880;
      2296: inst = 32'd268468224;
      2297: inst = 32'd201343518;
      2298: inst = 32'd203484854;
      2299: inst = 32'd136314880;
      2300: inst = 32'd268468224;
      2301: inst = 32'd201343519;
      2302: inst = 32'd203484854;
      2303: inst = 32'd136314880;
      2304: inst = 32'd268468224;
      2305: inst = 32'd201343520;
      2306: inst = 32'd203482839;
      2307: inst = 32'd136314880;
      2308: inst = 32'd268468224;
      2309: inst = 32'd201343521;
      2310: inst = 32'd203484855;
      2311: inst = 32'd136314880;
      2312: inst = 32'd268468224;
      2313: inst = 32'd201343522;
      2314: inst = 32'd203484854;
      2315: inst = 32'd136314880;
      2316: inst = 32'd268468224;
      2317: inst = 32'd201343523;
      2318: inst = 32'd203484854;
      2319: inst = 32'd136314880;
      2320: inst = 32'd268468224;
      2321: inst = 32'd201343524;
      2322: inst = 32'd203486870;
      2323: inst = 32'd136314880;
      2324: inst = 32'd268468224;
      2325: inst = 32'd201343525;
      2326: inst = 32'd203486870;
      2327: inst = 32'd136314880;
      2328: inst = 32'd268468224;
      2329: inst = 32'd201343526;
      2330: inst = 32'd203486870;
      2331: inst = 32'd136314880;
      2332: inst = 32'd268468224;
      2333: inst = 32'd201343527;
      2334: inst = 32'd203484854;
      2335: inst = 32'd136314880;
      2336: inst = 32'd268468224;
      2337: inst = 32'd201343528;
      2338: inst = 32'd203484855;
      2339: inst = 32'd136314880;
      2340: inst = 32'd268468224;
      2341: inst = 32'd201343529;
      2342: inst = 32'd203482807;
      2343: inst = 32'd136314880;
      2344: inst = 32'd268468224;
      2345: inst = 32'd201343530;
      2346: inst = 32'd203484887;
      2347: inst = 32'd136314880;
      2348: inst = 32'd268468224;
      2349: inst = 32'd201343531;
      2350: inst = 32'd203465871;
      2351: inst = 32'd136314880;
      2352: inst = 32'd268468224;
      2353: inst = 32'd201343532;
      2354: inst = 32'd203484855;
      2355: inst = 32'd136314880;
      2356: inst = 32'd268468224;
      2357: inst = 32'd201343533;
      2358: inst = 32'd203484855;
      2359: inst = 32'd136314880;
      2360: inst = 32'd268468224;
      2361: inst = 32'd201343534;
      2362: inst = 32'd203484823;
      2363: inst = 32'd136314880;
      2364: inst = 32'd268468224;
      2365: inst = 32'd201343535;
      2366: inst = 32'd203486871;
      2367: inst = 32'd136314880;
      2368: inst = 32'd268468224;
      2369: inst = 32'd201343536;
      2370: inst = 32'd203486902;
      2371: inst = 32'd136314880;
      2372: inst = 32'd268468224;
      2373: inst = 32'd201343537;
      2374: inst = 32'd203486902;
      2375: inst = 32'd136314880;
      2376: inst = 32'd268468224;
      2377: inst = 32'd201343538;
      2378: inst = 32'd203484854;
      2379: inst = 32'd136314880;
      2380: inst = 32'd268468224;
      2381: inst = 32'd201343539;
      2382: inst = 32'd203484854;
      2383: inst = 32'd136314880;
      2384: inst = 32'd268468224;
      2385: inst = 32'd201343540;
      2386: inst = 32'd203484854;
      2387: inst = 32'd136314880;
      2388: inst = 32'd268468224;
      2389: inst = 32'd201343541;
      2390: inst = 32'd203484854;
      2391: inst = 32'd136314880;
      2392: inst = 32'd268468224;
      2393: inst = 32'd201343542;
      2394: inst = 32'd203484854;
      2395: inst = 32'd136314880;
      2396: inst = 32'd268468224;
      2397: inst = 32'd201343543;
      2398: inst = 32'd203484854;
      2399: inst = 32'd136314880;
      2400: inst = 32'd268468224;
      2401: inst = 32'd201343544;
      2402: inst = 32'd203482774;
      2403: inst = 32'd136314880;
      2404: inst = 32'd268468224;
      2405: inst = 32'd201343545;
      2406: inst = 32'd203484855;
      2407: inst = 32'd136314880;
      2408: inst = 32'd268468224;
      2409: inst = 32'd201343546;
      2410: inst = 32'd203482775;
      2411: inst = 32'd136314880;
      2412: inst = 32'd268468224;
      2413: inst = 32'd201343547;
      2414: inst = 32'd203484888;
      2415: inst = 32'd136314880;
      2416: inst = 32'd268468224;
      2417: inst = 32'd201343548;
      2418: inst = 32'd203489212;
      2419: inst = 32'd136314880;
      2420: inst = 32'd268468224;
      2421: inst = 32'd201343549;
      2422: inst = 32'd203489278;
      2423: inst = 32'd136314880;
      2424: inst = 32'd268468224;
      2425: inst = 32'd201343550;
      2426: inst = 32'd203489279;
      2427: inst = 32'd136314880;
      2428: inst = 32'd268468224;
      2429: inst = 32'd201343551;
      2430: inst = 32'd203489279;
      2431: inst = 32'd136314880;
      2432: inst = 32'd268468224;
      2433: inst = 32'd201343552;
      2434: inst = 32'd203489279;
      2435: inst = 32'd136314880;
      2436: inst = 32'd268468224;
      2437: inst = 32'd201343553;
      2438: inst = 32'd203489279;
      2439: inst = 32'd136314880;
      2440: inst = 32'd268468224;
      2441: inst = 32'd201343554;
      2442: inst = 32'd203489279;
      2443: inst = 32'd136314880;
      2444: inst = 32'd268468224;
      2445: inst = 32'd201343555;
      2446: inst = 32'd203489279;
      2447: inst = 32'd136314880;
      2448: inst = 32'd268468224;
      2449: inst = 32'd201343556;
      2450: inst = 32'd203489279;
      2451: inst = 32'd136314880;
      2452: inst = 32'd268468224;
      2453: inst = 32'd201343557;
      2454: inst = 32'd203489279;
      2455: inst = 32'd136314880;
      2456: inst = 32'd268468224;
      2457: inst = 32'd201343558;
      2458: inst = 32'd203489279;
      2459: inst = 32'd136314880;
      2460: inst = 32'd268468224;
      2461: inst = 32'd201343559;
      2462: inst = 32'd203489279;
      2463: inst = 32'd136314880;
      2464: inst = 32'd268468224;
      2465: inst = 32'd201343560;
      2466: inst = 32'd203489279;
      2467: inst = 32'd136314880;
      2468: inst = 32'd268468224;
      2469: inst = 32'd201343561;
      2470: inst = 32'd203489279;
      2471: inst = 32'd136314880;
      2472: inst = 32'd268468224;
      2473: inst = 32'd201343562;
      2474: inst = 32'd203489279;
      2475: inst = 32'd136314880;
      2476: inst = 32'd268468224;
      2477: inst = 32'd201343563;
      2478: inst = 32'd203489279;
      2479: inst = 32'd136314880;
      2480: inst = 32'd268468224;
      2481: inst = 32'd201343564;
      2482: inst = 32'd203489279;
      2483: inst = 32'd136314880;
      2484: inst = 32'd268468224;
      2485: inst = 32'd201343565;
      2486: inst = 32'd203489279;
      2487: inst = 32'd136314880;
      2488: inst = 32'd268468224;
      2489: inst = 32'd201343566;
      2490: inst = 32'd203489279;
      2491: inst = 32'd136314880;
      2492: inst = 32'd268468224;
      2493: inst = 32'd201343567;
      2494: inst = 32'd203489279;
      2495: inst = 32'd136314880;
      2496: inst = 32'd268468224;
      2497: inst = 32'd201343568;
      2498: inst = 32'd203489279;
      2499: inst = 32'd136314880;
      2500: inst = 32'd268468224;
      2501: inst = 32'd201343569;
      2502: inst = 32'd203489279;
      2503: inst = 32'd136314880;
      2504: inst = 32'd268468224;
      2505: inst = 32'd201343570;
      2506: inst = 32'd203489279;
      2507: inst = 32'd136314880;
      2508: inst = 32'd268468224;
      2509: inst = 32'd201343571;
      2510: inst = 32'd203489279;
      2511: inst = 32'd136314880;
      2512: inst = 32'd268468224;
      2513: inst = 32'd201343572;
      2514: inst = 32'd203489279;
      2515: inst = 32'd136314880;
      2516: inst = 32'd268468224;
      2517: inst = 32'd201343573;
      2518: inst = 32'd203489279;
      2519: inst = 32'd136314880;
      2520: inst = 32'd268468224;
      2521: inst = 32'd201343574;
      2522: inst = 32'd203489279;
      2523: inst = 32'd136314880;
      2524: inst = 32'd268468224;
      2525: inst = 32'd201343575;
      2526: inst = 32'd203489279;
      2527: inst = 32'd136314880;
      2528: inst = 32'd268468224;
      2529: inst = 32'd201343576;
      2530: inst = 32'd203489279;
      2531: inst = 32'd136314880;
      2532: inst = 32'd268468224;
      2533: inst = 32'd201343577;
      2534: inst = 32'd203489279;
      2535: inst = 32'd136314880;
      2536: inst = 32'd268468224;
      2537: inst = 32'd201343578;
      2538: inst = 32'd203489279;
      2539: inst = 32'd136314880;
      2540: inst = 32'd268468224;
      2541: inst = 32'd201343579;
      2542: inst = 32'd203489279;
      2543: inst = 32'd136314880;
      2544: inst = 32'd268468224;
      2545: inst = 32'd201343580;
      2546: inst = 32'd203489279;
      2547: inst = 32'd136314880;
      2548: inst = 32'd268468224;
      2549: inst = 32'd201343581;
      2550: inst = 32'd203489279;
      2551: inst = 32'd136314880;
      2552: inst = 32'd268468224;
      2553: inst = 32'd201343582;
      2554: inst = 32'd203489279;
      2555: inst = 32'd136314880;
      2556: inst = 32'd268468224;
      2557: inst = 32'd201343583;
      2558: inst = 32'd203489279;
      2559: inst = 32'd136314880;
      2560: inst = 32'd268468224;
      2561: inst = 32'd201343584;
      2562: inst = 32'd203489279;
      2563: inst = 32'd136314880;
      2564: inst = 32'd268468224;
      2565: inst = 32'd201343585;
      2566: inst = 32'd203489279;
      2567: inst = 32'd136314880;
      2568: inst = 32'd268468224;
      2569: inst = 32'd201343586;
      2570: inst = 32'd203489278;
      2571: inst = 32'd136314880;
      2572: inst = 32'd268468224;
      2573: inst = 32'd201343587;
      2574: inst = 32'd203489212;
      2575: inst = 32'd136314880;
      2576: inst = 32'd268468224;
      2577: inst = 32'd201343588;
      2578: inst = 32'd203484888;
      2579: inst = 32'd136314880;
      2580: inst = 32'd268468224;
      2581: inst = 32'd201343589;
      2582: inst = 32'd203482775;
      2583: inst = 32'd136314880;
      2584: inst = 32'd268468224;
      2585: inst = 32'd201343590;
      2586: inst = 32'd203484855;
      2587: inst = 32'd136314880;
      2588: inst = 32'd268468224;
      2589: inst = 32'd201343591;
      2590: inst = 32'd203484822;
      2591: inst = 32'd136314880;
      2592: inst = 32'd268468224;
      2593: inst = 32'd201343592;
      2594: inst = 32'd203484854;
      2595: inst = 32'd136314880;
      2596: inst = 32'd268468224;
      2597: inst = 32'd201343593;
      2598: inst = 32'd203484854;
      2599: inst = 32'd136314880;
      2600: inst = 32'd268468224;
      2601: inst = 32'd201343594;
      2602: inst = 32'd203484854;
      2603: inst = 32'd136314880;
      2604: inst = 32'd268468224;
      2605: inst = 32'd201343595;
      2606: inst = 32'd203484854;
      2607: inst = 32'd136314880;
      2608: inst = 32'd268468224;
      2609: inst = 32'd201343596;
      2610: inst = 32'd203484854;
      2611: inst = 32'd136314880;
      2612: inst = 32'd268468224;
      2613: inst = 32'd201343597;
      2614: inst = 32'd203484854;
      2615: inst = 32'd136314880;
      2616: inst = 32'd268468224;
      2617: inst = 32'd201343598;
      2618: inst = 32'd203484854;
      2619: inst = 32'd136314880;
      2620: inst = 32'd268468224;
      2621: inst = 32'd201343599;
      2622: inst = 32'd203484854;
      2623: inst = 32'd136314880;
      2624: inst = 32'd268468224;
      2625: inst = 32'd201343600;
      2626: inst = 32'd203484854;
      2627: inst = 32'd136314880;
      2628: inst = 32'd268468224;
      2629: inst = 32'd201343601;
      2630: inst = 32'd203484854;
      2631: inst = 32'd136314880;
      2632: inst = 32'd268468224;
      2633: inst = 32'd201343602;
      2634: inst = 32'd203484854;
      2635: inst = 32'd136314880;
      2636: inst = 32'd268468224;
      2637: inst = 32'd201343603;
      2638: inst = 32'd203484854;
      2639: inst = 32'd136314880;
      2640: inst = 32'd268468224;
      2641: inst = 32'd201343604;
      2642: inst = 32'd203484854;
      2643: inst = 32'd136314880;
      2644: inst = 32'd268468224;
      2645: inst = 32'd201343605;
      2646: inst = 32'd203484854;
      2647: inst = 32'd136314880;
      2648: inst = 32'd268468224;
      2649: inst = 32'd201343606;
      2650: inst = 32'd203484854;
      2651: inst = 32'd136314880;
      2652: inst = 32'd268468224;
      2653: inst = 32'd201343607;
      2654: inst = 32'd203484854;
      2655: inst = 32'd136314880;
      2656: inst = 32'd268468224;
      2657: inst = 32'd201343608;
      2658: inst = 32'd203484854;
      2659: inst = 32'd136314880;
      2660: inst = 32'd268468224;
      2661: inst = 32'd201343609;
      2662: inst = 32'd203484854;
      2663: inst = 32'd136314880;
      2664: inst = 32'd268468224;
      2665: inst = 32'd201343610;
      2666: inst = 32'd203484854;
      2667: inst = 32'd136314880;
      2668: inst = 32'd268468224;
      2669: inst = 32'd201343611;
      2670: inst = 32'd203484854;
      2671: inst = 32'd136314880;
      2672: inst = 32'd268468224;
      2673: inst = 32'd201343612;
      2674: inst = 32'd203484854;
      2675: inst = 32'd136314880;
      2676: inst = 32'd268468224;
      2677: inst = 32'd201343613;
      2678: inst = 32'd203484854;
      2679: inst = 32'd136314880;
      2680: inst = 32'd268468224;
      2681: inst = 32'd201343614;
      2682: inst = 32'd203484854;
      2683: inst = 32'd136314880;
      2684: inst = 32'd268468224;
      2685: inst = 32'd201343615;
      2686: inst = 32'd203484854;
      2687: inst = 32'd136314880;
      2688: inst = 32'd268468224;
      2689: inst = 32'd201343616;
      2690: inst = 32'd203484854;
      2691: inst = 32'd136314880;
      2692: inst = 32'd268468224;
      2693: inst = 32'd201343617;
      2694: inst = 32'd203484854;
      2695: inst = 32'd136314880;
      2696: inst = 32'd268468224;
      2697: inst = 32'd201343618;
      2698: inst = 32'd203484854;
      2699: inst = 32'd136314880;
      2700: inst = 32'd268468224;
      2701: inst = 32'd201343619;
      2702: inst = 32'd203484854;
      2703: inst = 32'd136314880;
      2704: inst = 32'd268468224;
      2705: inst = 32'd201343620;
      2706: inst = 32'd203484854;
      2707: inst = 32'd136314880;
      2708: inst = 32'd268468224;
      2709: inst = 32'd201343621;
      2710: inst = 32'd203484854;
      2711: inst = 32'd136314880;
      2712: inst = 32'd268468224;
      2713: inst = 32'd201343622;
      2714: inst = 32'd203484854;
      2715: inst = 32'd136314880;
      2716: inst = 32'd268468224;
      2717: inst = 32'd201343623;
      2718: inst = 32'd203484886;
      2719: inst = 32'd136314880;
      2720: inst = 32'd268468224;
      2721: inst = 32'd201343624;
      2722: inst = 32'd203484886;
      2723: inst = 32'd136314880;
      2724: inst = 32'd268468224;
      2725: inst = 32'd201343625;
      2726: inst = 32'd203482838;
      2727: inst = 32'd136314880;
      2728: inst = 32'd268468224;
      2729: inst = 32'd201343626;
      2730: inst = 32'd203482838;
      2731: inst = 32'd136314880;
      2732: inst = 32'd268468224;
      2733: inst = 32'd201343627;
      2734: inst = 32'd203465901;
      2735: inst = 32'd136314880;
      2736: inst = 32'd268468224;
      2737: inst = 32'd201343628;
      2738: inst = 32'd203482838;
      2739: inst = 32'd136314880;
      2740: inst = 32'd268468224;
      2741: inst = 32'd201343629;
      2742: inst = 32'd203482837;
      2743: inst = 32'd136314880;
      2744: inst = 32'd268468224;
      2745: inst = 32'd201343630;
      2746: inst = 32'd203482837;
      2747: inst = 32'd136314880;
      2748: inst = 32'd268468224;
      2749: inst = 32'd201343631;
      2750: inst = 32'd203482870;
      2751: inst = 32'd136314880;
      2752: inst = 32'd268468224;
      2753: inst = 32'd201343632;
      2754: inst = 32'd203486902;
      2755: inst = 32'd136314880;
      2756: inst = 32'd268468224;
      2757: inst = 32'd201343633;
      2758: inst = 32'd203486902;
      2759: inst = 32'd136314880;
      2760: inst = 32'd268468224;
      2761: inst = 32'd201343634;
      2762: inst = 32'd203484854;
      2763: inst = 32'd136314880;
      2764: inst = 32'd268468224;
      2765: inst = 32'd201343635;
      2766: inst = 32'd203484854;
      2767: inst = 32'd136314880;
      2768: inst = 32'd268468224;
      2769: inst = 32'd201343636;
      2770: inst = 32'd203484854;
      2771: inst = 32'd136314880;
      2772: inst = 32'd268468224;
      2773: inst = 32'd201343637;
      2774: inst = 32'd203484854;
      2775: inst = 32'd136314880;
      2776: inst = 32'd268468224;
      2777: inst = 32'd201343638;
      2778: inst = 32'd203484854;
      2779: inst = 32'd136314880;
      2780: inst = 32'd268468224;
      2781: inst = 32'd201343639;
      2782: inst = 32'd203484854;
      2783: inst = 32'd136314880;
      2784: inst = 32'd268468224;
      2785: inst = 32'd201343640;
      2786: inst = 32'd203484887;
      2787: inst = 32'd136314880;
      2788: inst = 32'd268468224;
      2789: inst = 32'd201343641;
      2790: inst = 32'd203484887;
      2791: inst = 32'd136314880;
      2792: inst = 32'd268468224;
      2793: inst = 32'd201343642;
      2794: inst = 32'd203482807;
      2795: inst = 32'd136314880;
      2796: inst = 32'd268468224;
      2797: inst = 32'd201343643;
      2798: inst = 32'd203484888;
      2799: inst = 32'd136314880;
      2800: inst = 32'd268468224;
      2801: inst = 32'd201343644;
      2802: inst = 32'd203489278;
      2803: inst = 32'd136314880;
      2804: inst = 32'd268468224;
      2805: inst = 32'd201343645;
      2806: inst = 32'd203489279;
      2807: inst = 32'd136314880;
      2808: inst = 32'd268468224;
      2809: inst = 32'd201343646;
      2810: inst = 32'd203489279;
      2811: inst = 32'd136314880;
      2812: inst = 32'd268468224;
      2813: inst = 32'd201343647;
      2814: inst = 32'd203489279;
      2815: inst = 32'd136314880;
      2816: inst = 32'd268468224;
      2817: inst = 32'd201343648;
      2818: inst = 32'd203489279;
      2819: inst = 32'd136314880;
      2820: inst = 32'd268468224;
      2821: inst = 32'd201343649;
      2822: inst = 32'd203489279;
      2823: inst = 32'd136314880;
      2824: inst = 32'd268468224;
      2825: inst = 32'd201343650;
      2826: inst = 32'd203489279;
      2827: inst = 32'd136314880;
      2828: inst = 32'd268468224;
      2829: inst = 32'd201343651;
      2830: inst = 32'd203489279;
      2831: inst = 32'd136314880;
      2832: inst = 32'd268468224;
      2833: inst = 32'd201343652;
      2834: inst = 32'd203489279;
      2835: inst = 32'd136314880;
      2836: inst = 32'd268468224;
      2837: inst = 32'd201343653;
      2838: inst = 32'd203489279;
      2839: inst = 32'd136314880;
      2840: inst = 32'd268468224;
      2841: inst = 32'd201343654;
      2842: inst = 32'd203489279;
      2843: inst = 32'd136314880;
      2844: inst = 32'd268468224;
      2845: inst = 32'd201343655;
      2846: inst = 32'd203489279;
      2847: inst = 32'd136314880;
      2848: inst = 32'd268468224;
      2849: inst = 32'd201343656;
      2850: inst = 32'd203489279;
      2851: inst = 32'd136314880;
      2852: inst = 32'd268468224;
      2853: inst = 32'd201343657;
      2854: inst = 32'd203489279;
      2855: inst = 32'd136314880;
      2856: inst = 32'd268468224;
      2857: inst = 32'd201343658;
      2858: inst = 32'd203489279;
      2859: inst = 32'd136314880;
      2860: inst = 32'd268468224;
      2861: inst = 32'd201343659;
      2862: inst = 32'd203489279;
      2863: inst = 32'd136314880;
      2864: inst = 32'd268468224;
      2865: inst = 32'd201343660;
      2866: inst = 32'd203489279;
      2867: inst = 32'd136314880;
      2868: inst = 32'd268468224;
      2869: inst = 32'd201343661;
      2870: inst = 32'd203489279;
      2871: inst = 32'd136314880;
      2872: inst = 32'd268468224;
      2873: inst = 32'd201343662;
      2874: inst = 32'd203489279;
      2875: inst = 32'd136314880;
      2876: inst = 32'd268468224;
      2877: inst = 32'd201343663;
      2878: inst = 32'd203489279;
      2879: inst = 32'd136314880;
      2880: inst = 32'd268468224;
      2881: inst = 32'd201343664;
      2882: inst = 32'd203489279;
      2883: inst = 32'd136314880;
      2884: inst = 32'd268468224;
      2885: inst = 32'd201343665;
      2886: inst = 32'd203489279;
      2887: inst = 32'd136314880;
      2888: inst = 32'd268468224;
      2889: inst = 32'd201343666;
      2890: inst = 32'd203489279;
      2891: inst = 32'd136314880;
      2892: inst = 32'd268468224;
      2893: inst = 32'd201343667;
      2894: inst = 32'd203489279;
      2895: inst = 32'd136314880;
      2896: inst = 32'd268468224;
      2897: inst = 32'd201343668;
      2898: inst = 32'd203489279;
      2899: inst = 32'd136314880;
      2900: inst = 32'd268468224;
      2901: inst = 32'd201343669;
      2902: inst = 32'd203489279;
      2903: inst = 32'd136314880;
      2904: inst = 32'd268468224;
      2905: inst = 32'd201343670;
      2906: inst = 32'd203489279;
      2907: inst = 32'd136314880;
      2908: inst = 32'd268468224;
      2909: inst = 32'd201343671;
      2910: inst = 32'd203489279;
      2911: inst = 32'd136314880;
      2912: inst = 32'd268468224;
      2913: inst = 32'd201343672;
      2914: inst = 32'd203489279;
      2915: inst = 32'd136314880;
      2916: inst = 32'd268468224;
      2917: inst = 32'd201343673;
      2918: inst = 32'd203489279;
      2919: inst = 32'd136314880;
      2920: inst = 32'd268468224;
      2921: inst = 32'd201343674;
      2922: inst = 32'd203489279;
      2923: inst = 32'd136314880;
      2924: inst = 32'd268468224;
      2925: inst = 32'd201343675;
      2926: inst = 32'd203489279;
      2927: inst = 32'd136314880;
      2928: inst = 32'd268468224;
      2929: inst = 32'd201343676;
      2930: inst = 32'd203489279;
      2931: inst = 32'd136314880;
      2932: inst = 32'd268468224;
      2933: inst = 32'd201343677;
      2934: inst = 32'd203489279;
      2935: inst = 32'd136314880;
      2936: inst = 32'd268468224;
      2937: inst = 32'd201343678;
      2938: inst = 32'd203489279;
      2939: inst = 32'd136314880;
      2940: inst = 32'd268468224;
      2941: inst = 32'd201343679;
      2942: inst = 32'd203489279;
      2943: inst = 32'd136314880;
      2944: inst = 32'd268468224;
      2945: inst = 32'd201343680;
      2946: inst = 32'd203489279;
      2947: inst = 32'd136314880;
      2948: inst = 32'd268468224;
      2949: inst = 32'd201343681;
      2950: inst = 32'd203489279;
      2951: inst = 32'd136314880;
      2952: inst = 32'd268468224;
      2953: inst = 32'd201343682;
      2954: inst = 32'd203489279;
      2955: inst = 32'd136314880;
      2956: inst = 32'd268468224;
      2957: inst = 32'd201343683;
      2958: inst = 32'd203489278;
      2959: inst = 32'd136314880;
      2960: inst = 32'd268468224;
      2961: inst = 32'd201343684;
      2962: inst = 32'd203484888;
      2963: inst = 32'd136314880;
      2964: inst = 32'd268468224;
      2965: inst = 32'd201343685;
      2966: inst = 32'd203484855;
      2967: inst = 32'd136314880;
      2968: inst = 32'd268468224;
      2969: inst = 32'd201343686;
      2970: inst = 32'd203484887;
      2971: inst = 32'd136314880;
      2972: inst = 32'd268468224;
      2973: inst = 32'd201343687;
      2974: inst = 32'd203484855;
      2975: inst = 32'd136314880;
      2976: inst = 32'd268468224;
      2977: inst = 32'd201343688;
      2978: inst = 32'd203484854;
      2979: inst = 32'd136314880;
      2980: inst = 32'd268468224;
      2981: inst = 32'd201343689;
      2982: inst = 32'd203484854;
      2983: inst = 32'd136314880;
      2984: inst = 32'd268468224;
      2985: inst = 32'd201343690;
      2986: inst = 32'd203484854;
      2987: inst = 32'd136314880;
      2988: inst = 32'd268468224;
      2989: inst = 32'd201343691;
      2990: inst = 32'd203484854;
      2991: inst = 32'd136314880;
      2992: inst = 32'd268468224;
      2993: inst = 32'd201343692;
      2994: inst = 32'd203484854;
      2995: inst = 32'd136314880;
      2996: inst = 32'd268468224;
      2997: inst = 32'd201343693;
      2998: inst = 32'd203484854;
      2999: inst = 32'd136314880;
      3000: inst = 32'd268468224;
      3001: inst = 32'd201343694;
      3002: inst = 32'd203484854;
      3003: inst = 32'd136314880;
      3004: inst = 32'd268468224;
      3005: inst = 32'd201343695;
      3006: inst = 32'd203484854;
      3007: inst = 32'd136314880;
      3008: inst = 32'd268468224;
      3009: inst = 32'd201343696;
      3010: inst = 32'd203484854;
      3011: inst = 32'd136314880;
      3012: inst = 32'd268468224;
      3013: inst = 32'd201343697;
      3014: inst = 32'd203484854;
      3015: inst = 32'd136314880;
      3016: inst = 32'd268468224;
      3017: inst = 32'd201343698;
      3018: inst = 32'd203484854;
      3019: inst = 32'd136314880;
      3020: inst = 32'd268468224;
      3021: inst = 32'd201343699;
      3022: inst = 32'd203484854;
      3023: inst = 32'd136314880;
      3024: inst = 32'd268468224;
      3025: inst = 32'd201343700;
      3026: inst = 32'd203484854;
      3027: inst = 32'd136314880;
      3028: inst = 32'd268468224;
      3029: inst = 32'd201343701;
      3030: inst = 32'd203484854;
      3031: inst = 32'd136314880;
      3032: inst = 32'd268468224;
      3033: inst = 32'd201343702;
      3034: inst = 32'd203484854;
      3035: inst = 32'd136314880;
      3036: inst = 32'd268468224;
      3037: inst = 32'd201343703;
      3038: inst = 32'd203484854;
      3039: inst = 32'd136314880;
      3040: inst = 32'd268468224;
      3041: inst = 32'd201343704;
      3042: inst = 32'd203484854;
      3043: inst = 32'd136314880;
      3044: inst = 32'd268468224;
      3045: inst = 32'd201343705;
      3046: inst = 32'd203484854;
      3047: inst = 32'd136314880;
      3048: inst = 32'd268468224;
      3049: inst = 32'd201343706;
      3050: inst = 32'd203484854;
      3051: inst = 32'd136314880;
      3052: inst = 32'd268468224;
      3053: inst = 32'd201343707;
      3054: inst = 32'd203484854;
      3055: inst = 32'd136314880;
      3056: inst = 32'd268468224;
      3057: inst = 32'd201343708;
      3058: inst = 32'd203484854;
      3059: inst = 32'd136314880;
      3060: inst = 32'd268468224;
      3061: inst = 32'd201343709;
      3062: inst = 32'd203484854;
      3063: inst = 32'd136314880;
      3064: inst = 32'd268468224;
      3065: inst = 32'd201343710;
      3066: inst = 32'd203484854;
      3067: inst = 32'd136314880;
      3068: inst = 32'd268468224;
      3069: inst = 32'd201343711;
      3070: inst = 32'd203484854;
      3071: inst = 32'd136314880;
      3072: inst = 32'd268468224;
      3073: inst = 32'd201343712;
      3074: inst = 32'd203486903;
      3075: inst = 32'd136314880;
      3076: inst = 32'd268468224;
      3077: inst = 32'd201343713;
      3078: inst = 32'd203484790;
      3079: inst = 32'd136314880;
      3080: inst = 32'd268468224;
      3081: inst = 32'd201343714;
      3082: inst = 32'd203484822;
      3083: inst = 32'd136314880;
      3084: inst = 32'd268468224;
      3085: inst = 32'd201343715;
      3086: inst = 32'd203484887;
      3087: inst = 32'd136314880;
      3088: inst = 32'd268468224;
      3089: inst = 32'd201343716;
      3090: inst = 32'd203484919;
      3091: inst = 32'd136314880;
      3092: inst = 32'd268468224;
      3093: inst = 32'd201343717;
      3094: inst = 32'd203482806;
      3095: inst = 32'd136314880;
      3096: inst = 32'd268468224;
      3097: inst = 32'd201343718;
      3098: inst = 32'd203482805;
      3099: inst = 32'd136314880;
      3100: inst = 32'd268468224;
      3101: inst = 32'd201343719;
      3102: inst = 32'd203484885;
      3103: inst = 32'd136314880;
      3104: inst = 32'd268468224;
      3105: inst = 32'd201343720;
      3106: inst = 32'd203484821;
      3107: inst = 32'd136314880;
      3108: inst = 32'd268468224;
      3109: inst = 32'd201343721;
      3110: inst = 32'd203488982;
      3111: inst = 32'd136314880;
      3112: inst = 32'd268468224;
      3113: inst = 32'd201343722;
      3114: inst = 32'd203484723;
      3115: inst = 32'd136314880;
      3116: inst = 32'd268468224;
      3117: inst = 32'd201343723;
      3118: inst = 32'd203469964;
      3119: inst = 32'd136314880;
      3120: inst = 32'd268468224;
      3121: inst = 32'd201343724;
      3122: inst = 32'd203469964;
      3123: inst = 32'd136314880;
      3124: inst = 32'd268468224;
      3125: inst = 32'd201343725;
      3126: inst = 32'd203482707;
      3127: inst = 32'd136314880;
      3128: inst = 32'd268468224;
      3129: inst = 32'd201343726;
      3130: inst = 32'd203486965;
      3131: inst = 32'd136314880;
      3132: inst = 32'd268468224;
      3133: inst = 32'd201343727;
      3134: inst = 32'd203484852;
      3135: inst = 32'd136314880;
      3136: inst = 32'd268468224;
      3137: inst = 32'd201343728;
      3138: inst = 32'd203486902;
      3139: inst = 32'd136314880;
      3140: inst = 32'd268468224;
      3141: inst = 32'd201343729;
      3142: inst = 32'd203484822;
      3143: inst = 32'd136314880;
      3144: inst = 32'd268468224;
      3145: inst = 32'd201343730;
      3146: inst = 32'd203484854;
      3147: inst = 32'd136314880;
      3148: inst = 32'd268468224;
      3149: inst = 32'd201343731;
      3150: inst = 32'd203486935;
      3151: inst = 32'd136314880;
      3152: inst = 32'd268468224;
      3153: inst = 32'd201343732;
      3154: inst = 32'd203484887;
      3155: inst = 32'd136314880;
      3156: inst = 32'd268468224;
      3157: inst = 32'd201343733;
      3158: inst = 32'd203482774;
      3159: inst = 32'd136314880;
      3160: inst = 32'd268468224;
      3161: inst = 32'd201343734;
      3162: inst = 32'd203482774;
      3163: inst = 32'd136314880;
      3164: inst = 32'd268468224;
      3165: inst = 32'd201343735;
      3166: inst = 32'd203484887;
      3167: inst = 32'd136314880;
      3168: inst = 32'd268468224;
      3169: inst = 32'd201343736;
      3170: inst = 32'd203484855;
      3171: inst = 32'd136314880;
      3172: inst = 32'd268468224;
      3173: inst = 32'd201343737;
      3174: inst = 32'd203484855;
      3175: inst = 32'd136314880;
      3176: inst = 32'd268468224;
      3177: inst = 32'd201343738;
      3178: inst = 32'd203484888;
      3179: inst = 32'd136314880;
      3180: inst = 32'd268468224;
      3181: inst = 32'd201343739;
      3182: inst = 32'd203482808;
      3183: inst = 32'd136314880;
      3184: inst = 32'd268468224;
      3185: inst = 32'd201343740;
      3186: inst = 32'd203489278;
      3187: inst = 32'd136314880;
      3188: inst = 32'd268468224;
      3189: inst = 32'd201343741;
      3190: inst = 32'd203489279;
      3191: inst = 32'd136314880;
      3192: inst = 32'd268468224;
      3193: inst = 32'd201343742;
      3194: inst = 32'd203489279;
      3195: inst = 32'd136314880;
      3196: inst = 32'd268468224;
      3197: inst = 32'd201343743;
      3198: inst = 32'd203489279;
      3199: inst = 32'd136314880;
      3200: inst = 32'd268468224;
      3201: inst = 32'd201343744;
      3202: inst = 32'd203489279;
      3203: inst = 32'd136314880;
      3204: inst = 32'd268468224;
      3205: inst = 32'd201343745;
      3206: inst = 32'd203489279;
      3207: inst = 32'd136314880;
      3208: inst = 32'd268468224;
      3209: inst = 32'd201343746;
      3210: inst = 32'd203489279;
      3211: inst = 32'd136314880;
      3212: inst = 32'd268468224;
      3213: inst = 32'd201343747;
      3214: inst = 32'd203489279;
      3215: inst = 32'd136314880;
      3216: inst = 32'd268468224;
      3217: inst = 32'd201343748;
      3218: inst = 32'd203489279;
      3219: inst = 32'd136314880;
      3220: inst = 32'd268468224;
      3221: inst = 32'd201343749;
      3222: inst = 32'd203489279;
      3223: inst = 32'd136314880;
      3224: inst = 32'd268468224;
      3225: inst = 32'd201343750;
      3226: inst = 32'd203489279;
      3227: inst = 32'd136314880;
      3228: inst = 32'd268468224;
      3229: inst = 32'd201343751;
      3230: inst = 32'd203489279;
      3231: inst = 32'd136314880;
      3232: inst = 32'd268468224;
      3233: inst = 32'd201343752;
      3234: inst = 32'd203489279;
      3235: inst = 32'd136314880;
      3236: inst = 32'd268468224;
      3237: inst = 32'd201343753;
      3238: inst = 32'd203489279;
      3239: inst = 32'd136314880;
      3240: inst = 32'd268468224;
      3241: inst = 32'd201343754;
      3242: inst = 32'd203489279;
      3243: inst = 32'd136314880;
      3244: inst = 32'd268468224;
      3245: inst = 32'd201343755;
      3246: inst = 32'd203489279;
      3247: inst = 32'd136314880;
      3248: inst = 32'd268468224;
      3249: inst = 32'd201343756;
      3250: inst = 32'd203489279;
      3251: inst = 32'd136314880;
      3252: inst = 32'd268468224;
      3253: inst = 32'd201343757;
      3254: inst = 32'd203489279;
      3255: inst = 32'd136314880;
      3256: inst = 32'd268468224;
      3257: inst = 32'd201343758;
      3258: inst = 32'd203489279;
      3259: inst = 32'd136314880;
      3260: inst = 32'd268468224;
      3261: inst = 32'd201343759;
      3262: inst = 32'd203489279;
      3263: inst = 32'd136314880;
      3264: inst = 32'd268468224;
      3265: inst = 32'd201343760;
      3266: inst = 32'd203489279;
      3267: inst = 32'd136314880;
      3268: inst = 32'd268468224;
      3269: inst = 32'd201343761;
      3270: inst = 32'd203489279;
      3271: inst = 32'd136314880;
      3272: inst = 32'd268468224;
      3273: inst = 32'd201343762;
      3274: inst = 32'd203489279;
      3275: inst = 32'd136314880;
      3276: inst = 32'd268468224;
      3277: inst = 32'd201343763;
      3278: inst = 32'd203489279;
      3279: inst = 32'd136314880;
      3280: inst = 32'd268468224;
      3281: inst = 32'd201343764;
      3282: inst = 32'd203489279;
      3283: inst = 32'd136314880;
      3284: inst = 32'd268468224;
      3285: inst = 32'd201343765;
      3286: inst = 32'd203489279;
      3287: inst = 32'd136314880;
      3288: inst = 32'd268468224;
      3289: inst = 32'd201343766;
      3290: inst = 32'd203489279;
      3291: inst = 32'd136314880;
      3292: inst = 32'd268468224;
      3293: inst = 32'd201343767;
      3294: inst = 32'd203489279;
      3295: inst = 32'd136314880;
      3296: inst = 32'd268468224;
      3297: inst = 32'd201343768;
      3298: inst = 32'd203489279;
      3299: inst = 32'd136314880;
      3300: inst = 32'd268468224;
      3301: inst = 32'd201343769;
      3302: inst = 32'd203489279;
      3303: inst = 32'd136314880;
      3304: inst = 32'd268468224;
      3305: inst = 32'd201343770;
      3306: inst = 32'd203489279;
      3307: inst = 32'd136314880;
      3308: inst = 32'd268468224;
      3309: inst = 32'd201343771;
      3310: inst = 32'd203489279;
      3311: inst = 32'd136314880;
      3312: inst = 32'd268468224;
      3313: inst = 32'd201343772;
      3314: inst = 32'd203489279;
      3315: inst = 32'd136314880;
      3316: inst = 32'd268468224;
      3317: inst = 32'd201343773;
      3318: inst = 32'd203489279;
      3319: inst = 32'd136314880;
      3320: inst = 32'd268468224;
      3321: inst = 32'd201343774;
      3322: inst = 32'd203489279;
      3323: inst = 32'd136314880;
      3324: inst = 32'd268468224;
      3325: inst = 32'd201343775;
      3326: inst = 32'd203489279;
      3327: inst = 32'd136314880;
      3328: inst = 32'd268468224;
      3329: inst = 32'd201343776;
      3330: inst = 32'd203489279;
      3331: inst = 32'd136314880;
      3332: inst = 32'd268468224;
      3333: inst = 32'd201343777;
      3334: inst = 32'd203489279;
      3335: inst = 32'd136314880;
      3336: inst = 32'd268468224;
      3337: inst = 32'd201343778;
      3338: inst = 32'd203489279;
      3339: inst = 32'd136314880;
      3340: inst = 32'd268468224;
      3341: inst = 32'd201343779;
      3342: inst = 32'd203489278;
      3343: inst = 32'd136314880;
      3344: inst = 32'd268468224;
      3345: inst = 32'd201343780;
      3346: inst = 32'd203482808;
      3347: inst = 32'd136314880;
      3348: inst = 32'd268468224;
      3349: inst = 32'd201343781;
      3350: inst = 32'd203484856;
      3351: inst = 32'd136314880;
      3352: inst = 32'd268468224;
      3353: inst = 32'd201343782;
      3354: inst = 32'd203484855;
      3355: inst = 32'd136314880;
      3356: inst = 32'd268468224;
      3357: inst = 32'd201343783;
      3358: inst = 32'd203484855;
      3359: inst = 32'd136314880;
      3360: inst = 32'd268468224;
      3361: inst = 32'd201343784;
      3362: inst = 32'd203484854;
      3363: inst = 32'd136314880;
      3364: inst = 32'd268468224;
      3365: inst = 32'd201343785;
      3366: inst = 32'd203484854;
      3367: inst = 32'd136314880;
      3368: inst = 32'd268468224;
      3369: inst = 32'd201343786;
      3370: inst = 32'd203484854;
      3371: inst = 32'd136314880;
      3372: inst = 32'd268468224;
      3373: inst = 32'd201343787;
      3374: inst = 32'd203484854;
      3375: inst = 32'd136314880;
      3376: inst = 32'd268468224;
      3377: inst = 32'd201343788;
      3378: inst = 32'd203484854;
      3379: inst = 32'd136314880;
      3380: inst = 32'd268468224;
      3381: inst = 32'd201343789;
      3382: inst = 32'd203484854;
      3383: inst = 32'd136314880;
      3384: inst = 32'd268468224;
      3385: inst = 32'd201343790;
      3386: inst = 32'd203484854;
      3387: inst = 32'd136314880;
      3388: inst = 32'd268468224;
      3389: inst = 32'd201343791;
      3390: inst = 32'd203484854;
      3391: inst = 32'd136314880;
      3392: inst = 32'd268468224;
      3393: inst = 32'd201343792;
      3394: inst = 32'd203484854;
      3395: inst = 32'd136314880;
      3396: inst = 32'd268468224;
      3397: inst = 32'd201343793;
      3398: inst = 32'd203484854;
      3399: inst = 32'd136314880;
      3400: inst = 32'd268468224;
      3401: inst = 32'd201343794;
      3402: inst = 32'd203484854;
      3403: inst = 32'd136314880;
      3404: inst = 32'd268468224;
      3405: inst = 32'd201343795;
      3406: inst = 32'd203484854;
      3407: inst = 32'd136314880;
      3408: inst = 32'd268468224;
      3409: inst = 32'd201343796;
      3410: inst = 32'd203484854;
      3411: inst = 32'd136314880;
      3412: inst = 32'd268468224;
      3413: inst = 32'd201343797;
      3414: inst = 32'd203484854;
      3415: inst = 32'd136314880;
      3416: inst = 32'd268468224;
      3417: inst = 32'd201343798;
      3418: inst = 32'd203484854;
      3419: inst = 32'd136314880;
      3420: inst = 32'd268468224;
      3421: inst = 32'd201343799;
      3422: inst = 32'd203484854;
      3423: inst = 32'd136314880;
      3424: inst = 32'd268468224;
      3425: inst = 32'd201343800;
      3426: inst = 32'd203484854;
      3427: inst = 32'd136314880;
      3428: inst = 32'd268468224;
      3429: inst = 32'd201343801;
      3430: inst = 32'd203484854;
      3431: inst = 32'd136314880;
      3432: inst = 32'd268468224;
      3433: inst = 32'd201343802;
      3434: inst = 32'd203484854;
      3435: inst = 32'd136314880;
      3436: inst = 32'd268468224;
      3437: inst = 32'd201343803;
      3438: inst = 32'd203484854;
      3439: inst = 32'd136314880;
      3440: inst = 32'd268468224;
      3441: inst = 32'd201343804;
      3442: inst = 32'd203484854;
      3443: inst = 32'd136314880;
      3444: inst = 32'd268468224;
      3445: inst = 32'd201343805;
      3446: inst = 32'd203484854;
      3447: inst = 32'd136314880;
      3448: inst = 32'd268468224;
      3449: inst = 32'd201343806;
      3450: inst = 32'd203484854;
      3451: inst = 32'd136314880;
      3452: inst = 32'd268468224;
      3453: inst = 32'd201343807;
      3454: inst = 32'd203484854;
      3455: inst = 32'd136314880;
      3456: inst = 32'd268468224;
      3457: inst = 32'd201343808;
      3458: inst = 32'd203486870;
      3459: inst = 32'd136314880;
      3460: inst = 32'd268468224;
      3461: inst = 32'd201343809;
      3462: inst = 32'd203486902;
      3463: inst = 32'd136314880;
      3464: inst = 32'd268468224;
      3465: inst = 32'd201343810;
      3466: inst = 32'd203484886;
      3467: inst = 32'd136314880;
      3468: inst = 32'd268468224;
      3469: inst = 32'd201343811;
      3470: inst = 32'd203482806;
      3471: inst = 32'd136314880;
      3472: inst = 32'd268468224;
      3473: inst = 32'd201343812;
      3474: inst = 32'd203482806;
      3475: inst = 32'd136314880;
      3476: inst = 32'd268468224;
      3477: inst = 32'd201343813;
      3478: inst = 32'd203482805;
      3479: inst = 32'd136314880;
      3480: inst = 32'd268468224;
      3481: inst = 32'd201343814;
      3482: inst = 32'd203484853;
      3483: inst = 32'd136314880;
      3484: inst = 32'd268468224;
      3485: inst = 32'd201343815;
      3486: inst = 32'd203488917;
      3487: inst = 32'd136314880;
      3488: inst = 32'd268468224;
      3489: inst = 32'd201343816;
      3490: inst = 32'd203488852;
      3491: inst = 32'd136314880;
      3492: inst = 32'd268468224;
      3493: inst = 32'd201343817;
      3494: inst = 32'd203484496;
      3495: inst = 32'd136314880;
      3496: inst = 32'd268468224;
      3497: inst = 32'd201343818;
      3498: inst = 32'd203471721;
      3499: inst = 32'd136314880;
      3500: inst = 32'd268468224;
      3501: inst = 32'd201343819;
      3502: inst = 32'd203471656;
      3503: inst = 32'd136314880;
      3504: inst = 32'd268468224;
      3505: inst = 32'd201343820;
      3506: inst = 32'd203469608;
      3507: inst = 32'd136314880;
      3508: inst = 32'd268468224;
      3509: inst = 32'd201343821;
      3510: inst = 32'd203471753;
      3511: inst = 32'd136314880;
      3512: inst = 32'd268468224;
      3513: inst = 32'd201343822;
      3514: inst = 32'd203484495;
      3515: inst = 32'd136314880;
      3516: inst = 32'd268468224;
      3517: inst = 32'd201343823;
      3518: inst = 32'd203488851;
      3519: inst = 32'd136314880;
      3520: inst = 32'd268468224;
      3521: inst = 32'd201343824;
      3522: inst = 32'd203486902;
      3523: inst = 32'd136314880;
      3524: inst = 32'd268468224;
      3525: inst = 32'd201343825;
      3526: inst = 32'd203486870;
      3527: inst = 32'd136314880;
      3528: inst = 32'd268468224;
      3529: inst = 32'd201343826;
      3530: inst = 32'd203484822;
      3531: inst = 32'd136314880;
      3532: inst = 32'd268468224;
      3533: inst = 32'd201343827;
      3534: inst = 32'd203484822;
      3535: inst = 32'd136314880;
      3536: inst = 32'd268468224;
      3537: inst = 32'd201343828;
      3538: inst = 32'd203484854;
      3539: inst = 32'd136314880;
      3540: inst = 32'd268468224;
      3541: inst = 32'd201343829;
      3542: inst = 32'd203484886;
      3543: inst = 32'd136314880;
      3544: inst = 32'd268468224;
      3545: inst = 32'd201343830;
      3546: inst = 32'd203484886;
      3547: inst = 32'd136314880;
      3548: inst = 32'd268468224;
      3549: inst = 32'd201343831;
      3550: inst = 32'd203484854;
      3551: inst = 32'd136314880;
      3552: inst = 32'd268468224;
      3553: inst = 32'd201343832;
      3554: inst = 32'd203484854;
      3555: inst = 32'd136314880;
      3556: inst = 32'd268468224;
      3557: inst = 32'd201343833;
      3558: inst = 32'd203484855;
      3559: inst = 32'd136314880;
      3560: inst = 32'd268468224;
      3561: inst = 32'd201343834;
      3562: inst = 32'd203484888;
      3563: inst = 32'd136314880;
      3564: inst = 32'd268468224;
      3565: inst = 32'd201343835;
      3566: inst = 32'd203482808;
      3567: inst = 32'd136314880;
      3568: inst = 32'd268468224;
      3569: inst = 32'd201343836;
      3570: inst = 32'd203489278;
      3571: inst = 32'd136314880;
      3572: inst = 32'd268468224;
      3573: inst = 32'd201343837;
      3574: inst = 32'd203489279;
      3575: inst = 32'd136314880;
      3576: inst = 32'd268468224;
      3577: inst = 32'd201343838;
      3578: inst = 32'd203489279;
      3579: inst = 32'd136314880;
      3580: inst = 32'd268468224;
      3581: inst = 32'd201343839;
      3582: inst = 32'd203489279;
      3583: inst = 32'd136314880;
      3584: inst = 32'd268468224;
      3585: inst = 32'd201343840;
      3586: inst = 32'd203489279;
      3587: inst = 32'd136314880;
      3588: inst = 32'd268468224;
      3589: inst = 32'd201343841;
      3590: inst = 32'd203489279;
      3591: inst = 32'd136314880;
      3592: inst = 32'd268468224;
      3593: inst = 32'd201343842;
      3594: inst = 32'd203489279;
      3595: inst = 32'd136314880;
      3596: inst = 32'd268468224;
      3597: inst = 32'd201343843;
      3598: inst = 32'd203489279;
      3599: inst = 32'd136314880;
      3600: inst = 32'd268468224;
      3601: inst = 32'd201343844;
      3602: inst = 32'd203489279;
      3603: inst = 32'd136314880;
      3604: inst = 32'd268468224;
      3605: inst = 32'd201343845;
      3606: inst = 32'd203489279;
      3607: inst = 32'd136314880;
      3608: inst = 32'd268468224;
      3609: inst = 32'd201343846;
      3610: inst = 32'd203489279;
      3611: inst = 32'd136314880;
      3612: inst = 32'd268468224;
      3613: inst = 32'd201343847;
      3614: inst = 32'd203489279;
      3615: inst = 32'd136314880;
      3616: inst = 32'd268468224;
      3617: inst = 32'd201343848;
      3618: inst = 32'd203489279;
      3619: inst = 32'd136314880;
      3620: inst = 32'd268468224;
      3621: inst = 32'd201343849;
      3622: inst = 32'd203489279;
      3623: inst = 32'd136314880;
      3624: inst = 32'd268468224;
      3625: inst = 32'd201343850;
      3626: inst = 32'd203489279;
      3627: inst = 32'd136314880;
      3628: inst = 32'd268468224;
      3629: inst = 32'd201343851;
      3630: inst = 32'd203489279;
      3631: inst = 32'd136314880;
      3632: inst = 32'd268468224;
      3633: inst = 32'd201343852;
      3634: inst = 32'd203489279;
      3635: inst = 32'd136314880;
      3636: inst = 32'd268468224;
      3637: inst = 32'd201343853;
      3638: inst = 32'd203489279;
      3639: inst = 32'd136314880;
      3640: inst = 32'd268468224;
      3641: inst = 32'd201343854;
      3642: inst = 32'd203489279;
      3643: inst = 32'd136314880;
      3644: inst = 32'd268468224;
      3645: inst = 32'd201343855;
      3646: inst = 32'd203489279;
      3647: inst = 32'd136314880;
      3648: inst = 32'd268468224;
      3649: inst = 32'd201343856;
      3650: inst = 32'd203489279;
      3651: inst = 32'd136314880;
      3652: inst = 32'd268468224;
      3653: inst = 32'd201343857;
      3654: inst = 32'd203489279;
      3655: inst = 32'd136314880;
      3656: inst = 32'd268468224;
      3657: inst = 32'd201343858;
      3658: inst = 32'd203489279;
      3659: inst = 32'd136314880;
      3660: inst = 32'd268468224;
      3661: inst = 32'd201343859;
      3662: inst = 32'd203489279;
      3663: inst = 32'd136314880;
      3664: inst = 32'd268468224;
      3665: inst = 32'd201343860;
      3666: inst = 32'd203489279;
      3667: inst = 32'd136314880;
      3668: inst = 32'd268468224;
      3669: inst = 32'd201343861;
      3670: inst = 32'd203489279;
      3671: inst = 32'd136314880;
      3672: inst = 32'd268468224;
      3673: inst = 32'd201343862;
      3674: inst = 32'd203489279;
      3675: inst = 32'd136314880;
      3676: inst = 32'd268468224;
      3677: inst = 32'd201343863;
      3678: inst = 32'd203489279;
      3679: inst = 32'd136314880;
      3680: inst = 32'd268468224;
      3681: inst = 32'd201343864;
      3682: inst = 32'd203489279;
      3683: inst = 32'd136314880;
      3684: inst = 32'd268468224;
      3685: inst = 32'd201343865;
      3686: inst = 32'd203489279;
      3687: inst = 32'd136314880;
      3688: inst = 32'd268468224;
      3689: inst = 32'd201343866;
      3690: inst = 32'd203489279;
      3691: inst = 32'd136314880;
      3692: inst = 32'd268468224;
      3693: inst = 32'd201343867;
      3694: inst = 32'd203489279;
      3695: inst = 32'd136314880;
      3696: inst = 32'd268468224;
      3697: inst = 32'd201343868;
      3698: inst = 32'd203489279;
      3699: inst = 32'd136314880;
      3700: inst = 32'd268468224;
      3701: inst = 32'd201343869;
      3702: inst = 32'd203489279;
      3703: inst = 32'd136314880;
      3704: inst = 32'd268468224;
      3705: inst = 32'd201343870;
      3706: inst = 32'd203489279;
      3707: inst = 32'd136314880;
      3708: inst = 32'd268468224;
      3709: inst = 32'd201343871;
      3710: inst = 32'd203489279;
      3711: inst = 32'd136314880;
      3712: inst = 32'd268468224;
      3713: inst = 32'd201343872;
      3714: inst = 32'd203489279;
      3715: inst = 32'd136314880;
      3716: inst = 32'd268468224;
      3717: inst = 32'd201343873;
      3718: inst = 32'd203489279;
      3719: inst = 32'd136314880;
      3720: inst = 32'd268468224;
      3721: inst = 32'd201343874;
      3722: inst = 32'd203489279;
      3723: inst = 32'd136314880;
      3724: inst = 32'd268468224;
      3725: inst = 32'd201343875;
      3726: inst = 32'd203489278;
      3727: inst = 32'd136314880;
      3728: inst = 32'd268468224;
      3729: inst = 32'd201343876;
      3730: inst = 32'd203482808;
      3731: inst = 32'd136314880;
      3732: inst = 32'd268468224;
      3733: inst = 32'd201343877;
      3734: inst = 32'd203484856;
      3735: inst = 32'd136314880;
      3736: inst = 32'd268468224;
      3737: inst = 32'd201343878;
      3738: inst = 32'd203484855;
      3739: inst = 32'd136314880;
      3740: inst = 32'd268468224;
      3741: inst = 32'd201343879;
      3742: inst = 32'd203484854;
      3743: inst = 32'd136314880;
      3744: inst = 32'd268468224;
      3745: inst = 32'd201343880;
      3746: inst = 32'd203484854;
      3747: inst = 32'd136314880;
      3748: inst = 32'd268468224;
      3749: inst = 32'd201343881;
      3750: inst = 32'd203484854;
      3751: inst = 32'd136314880;
      3752: inst = 32'd268468224;
      3753: inst = 32'd201343882;
      3754: inst = 32'd203484854;
      3755: inst = 32'd136314880;
      3756: inst = 32'd268468224;
      3757: inst = 32'd201343883;
      3758: inst = 32'd203484854;
      3759: inst = 32'd136314880;
      3760: inst = 32'd268468224;
      3761: inst = 32'd201343884;
      3762: inst = 32'd203484854;
      3763: inst = 32'd136314880;
      3764: inst = 32'd268468224;
      3765: inst = 32'd201343885;
      3766: inst = 32'd203484854;
      3767: inst = 32'd136314880;
      3768: inst = 32'd268468224;
      3769: inst = 32'd201343886;
      3770: inst = 32'd203484854;
      3771: inst = 32'd136314880;
      3772: inst = 32'd268468224;
      3773: inst = 32'd201343887;
      3774: inst = 32'd203484854;
      3775: inst = 32'd136314880;
      3776: inst = 32'd268468224;
      3777: inst = 32'd201343888;
      3778: inst = 32'd203486934;
      3779: inst = 32'd136314880;
      3780: inst = 32'd268468224;
      3781: inst = 32'd201343889;
      3782: inst = 32'd203484886;
      3783: inst = 32'd136314880;
      3784: inst = 32'd268468224;
      3785: inst = 32'd201343890;
      3786: inst = 32'd203484886;
      3787: inst = 32'd136314880;
      3788: inst = 32'd268468224;
      3789: inst = 32'd201343891;
      3790: inst = 32'd203484886;
      3791: inst = 32'd136314880;
      3792: inst = 32'd268468224;
      3793: inst = 32'd201343892;
      3794: inst = 32'd203484886;
      3795: inst = 32'd136314880;
      3796: inst = 32'd268468224;
      3797: inst = 32'd201343893;
      3798: inst = 32'd203484854;
      3799: inst = 32'd136314880;
      3800: inst = 32'd268468224;
      3801: inst = 32'd201343894;
      3802: inst = 32'd203484886;
      3803: inst = 32'd136314880;
      3804: inst = 32'd268468224;
      3805: inst = 32'd201343895;
      3806: inst = 32'd203486934;
      3807: inst = 32'd136314880;
      3808: inst = 32'd268468224;
      3809: inst = 32'd201343896;
      3810: inst = 32'd203484854;
      3811: inst = 32'd136314880;
      3812: inst = 32'd268468224;
      3813: inst = 32'd201343897;
      3814: inst = 32'd203484854;
      3815: inst = 32'd136314880;
      3816: inst = 32'd268468224;
      3817: inst = 32'd201343898;
      3818: inst = 32'd203484854;
      3819: inst = 32'd136314880;
      3820: inst = 32'd268468224;
      3821: inst = 32'd201343899;
      3822: inst = 32'd203484854;
      3823: inst = 32'd136314880;
      3824: inst = 32'd268468224;
      3825: inst = 32'd201343900;
      3826: inst = 32'd203484854;
      3827: inst = 32'd136314880;
      3828: inst = 32'd268468224;
      3829: inst = 32'd201343901;
      3830: inst = 32'd203484854;
      3831: inst = 32'd136314880;
      3832: inst = 32'd268468224;
      3833: inst = 32'd201343902;
      3834: inst = 32'd203484854;
      3835: inst = 32'd136314880;
      3836: inst = 32'd268468224;
      3837: inst = 32'd201343903;
      3838: inst = 32'd203484854;
      3839: inst = 32'd136314880;
      3840: inst = 32'd268468224;
      3841: inst = 32'd201343904;
      3842: inst = 32'd203484789;
      3843: inst = 32'd136314880;
      3844: inst = 32'd268468224;
      3845: inst = 32'd201343905;
      3846: inst = 32'd203486935;
      3847: inst = 32'd136314880;
      3848: inst = 32'd268468224;
      3849: inst = 32'd201343906;
      3850: inst = 32'd203484919;
      3851: inst = 32'd136314880;
      3852: inst = 32'd268468224;
      3853: inst = 32'd201343907;
      3854: inst = 32'd203482806;
      3855: inst = 32'd136314880;
      3856: inst = 32'd268468224;
      3857: inst = 32'd201343908;
      3858: inst = 32'd203482838;
      3859: inst = 32'd136314880;
      3860: inst = 32'd268468224;
      3861: inst = 32'd201343909;
      3862: inst = 32'd203484918;
      3863: inst = 32'd136314880;
      3864: inst = 32'd268468224;
      3865: inst = 32'd201343910;
      3866: inst = 32'd203486902;
      3867: inst = 32'd136314880;
      3868: inst = 32'd268468224;
      3869: inst = 32'd201343911;
      3870: inst = 32'd203488852;
      3871: inst = 32'd136314880;
      3872: inst = 32'd268468224;
      3873: inst = 32'd201343912;
      3874: inst = 32'd203478093;
      3875: inst = 32'd136314880;
      3876: inst = 32'd268468224;
      3877: inst = 32'd201343913;
      3878: inst = 32'd203471591;
      3879: inst = 32'd136314880;
      3880: inst = 32'd268468224;
      3881: inst = 32'd201343914;
      3882: inst = 32'd203475655;
      3883: inst = 32'd136314880;
      3884: inst = 32'd268468224;
      3885: inst = 32'd201343915;
      3886: inst = 32'd203475622;
      3887: inst = 32'd136314880;
      3888: inst = 32'd268468224;
      3889: inst = 32'd201343916;
      3890: inst = 32'd203475622;
      3891: inst = 32'd136314880;
      3892: inst = 32'd268468224;
      3893: inst = 32'd201343917;
      3894: inst = 32'd203473607;
      3895: inst = 32'd136314880;
      3896: inst = 32'd268468224;
      3897: inst = 32'd201343918;
      3898: inst = 32'd203473639;
      3899: inst = 32'd136314880;
      3900: inst = 32'd268468224;
      3901: inst = 32'd201343919;
      3902: inst = 32'd203482123;
      3903: inst = 32'd136314880;
      3904: inst = 32'd268468224;
      3905: inst = 32'd201343920;
      3906: inst = 32'd203484822;
      3907: inst = 32'd136314880;
      3908: inst = 32'd268468224;
      3909: inst = 32'd201343921;
      3910: inst = 32'd203486902;
      3911: inst = 32'd136314880;
      3912: inst = 32'd268468224;
      3913: inst = 32'd201343922;
      3914: inst = 32'd203486935;
      3915: inst = 32'd136314880;
      3916: inst = 32'd268468224;
      3917: inst = 32'd201343923;
      3918: inst = 32'd203484822;
      3919: inst = 32'd136314880;
      3920: inst = 32'd268468224;
      3921: inst = 32'd201343924;
      3922: inst = 32'd203484854;
      3923: inst = 32'd136314880;
      3924: inst = 32'd268468224;
      3925: inst = 32'd201343925;
      3926: inst = 32'd203486967;
      3927: inst = 32'd136314880;
      3928: inst = 32'd268468224;
      3929: inst = 32'd201343926;
      3930: inst = 32'd203484887;
      3931: inst = 32'd136314880;
      3932: inst = 32'd268468224;
      3933: inst = 32'd201343927;
      3934: inst = 32'd203482774;
      3935: inst = 32'd136314880;
      3936: inst = 32'd268468224;
      3937: inst = 32'd201343928;
      3938: inst = 32'd203484854;
      3939: inst = 32'd136314880;
      3940: inst = 32'd268468224;
      3941: inst = 32'd201343929;
      3942: inst = 32'd203484855;
      3943: inst = 32'd136314880;
      3944: inst = 32'd268468224;
      3945: inst = 32'd201343930;
      3946: inst = 32'd203484887;
      3947: inst = 32'd136314880;
      3948: inst = 32'd268468224;
      3949: inst = 32'd201343931;
      3950: inst = 32'd203482808;
      3951: inst = 32'd136314880;
      3952: inst = 32'd268468224;
      3953: inst = 32'd201343932;
      3954: inst = 32'd203489278;
      3955: inst = 32'd136314880;
      3956: inst = 32'd268468224;
      3957: inst = 32'd201343933;
      3958: inst = 32'd203489279;
      3959: inst = 32'd136314880;
      3960: inst = 32'd268468224;
      3961: inst = 32'd201343934;
      3962: inst = 32'd203489279;
      3963: inst = 32'd136314880;
      3964: inst = 32'd268468224;
      3965: inst = 32'd201343935;
      3966: inst = 32'd203489279;
      3967: inst = 32'd136314880;
      3968: inst = 32'd268468224;
      3969: inst = 32'd201343936;
      3970: inst = 32'd203489279;
      3971: inst = 32'd136314880;
      3972: inst = 32'd268468224;
      3973: inst = 32'd201343937;
      3974: inst = 32'd203489279;
      3975: inst = 32'd136314880;
      3976: inst = 32'd268468224;
      3977: inst = 32'd201343938;
      3978: inst = 32'd203489279;
      3979: inst = 32'd136314880;
      3980: inst = 32'd268468224;
      3981: inst = 32'd201343939;
      3982: inst = 32'd203489279;
      3983: inst = 32'd136314880;
      3984: inst = 32'd268468224;
      3985: inst = 32'd201343940;
      3986: inst = 32'd203489279;
      3987: inst = 32'd136314880;
      3988: inst = 32'd268468224;
      3989: inst = 32'd201343941;
      3990: inst = 32'd203489279;
      3991: inst = 32'd136314880;
      3992: inst = 32'd268468224;
      3993: inst = 32'd201343942;
      3994: inst = 32'd203489279;
      3995: inst = 32'd136314880;
      3996: inst = 32'd268468224;
      3997: inst = 32'd201343943;
      3998: inst = 32'd203489279;
      3999: inst = 32'd136314880;
      4000: inst = 32'd268468224;
      4001: inst = 32'd201343944;
      4002: inst = 32'd203489279;
      4003: inst = 32'd136314880;
      4004: inst = 32'd268468224;
      4005: inst = 32'd201343945;
      4006: inst = 32'd203489279;
      4007: inst = 32'd136314880;
      4008: inst = 32'd268468224;
      4009: inst = 32'd201343946;
      4010: inst = 32'd203489279;
      4011: inst = 32'd136314880;
      4012: inst = 32'd268468224;
      4013: inst = 32'd201343947;
      4014: inst = 32'd203489279;
      4015: inst = 32'd136314880;
      4016: inst = 32'd268468224;
      4017: inst = 32'd201343948;
      4018: inst = 32'd203489279;
      4019: inst = 32'd136314880;
      4020: inst = 32'd268468224;
      4021: inst = 32'd201343949;
      4022: inst = 32'd203489279;
      4023: inst = 32'd136314880;
      4024: inst = 32'd268468224;
      4025: inst = 32'd201343950;
      4026: inst = 32'd203489279;
      4027: inst = 32'd136314880;
      4028: inst = 32'd268468224;
      4029: inst = 32'd201343951;
      4030: inst = 32'd203489279;
      4031: inst = 32'd136314880;
      4032: inst = 32'd268468224;
      4033: inst = 32'd201343952;
      4034: inst = 32'd203489279;
      4035: inst = 32'd136314880;
      4036: inst = 32'd268468224;
      4037: inst = 32'd201343953;
      4038: inst = 32'd203489279;
      4039: inst = 32'd136314880;
      4040: inst = 32'd268468224;
      4041: inst = 32'd201343954;
      4042: inst = 32'd203489279;
      4043: inst = 32'd136314880;
      4044: inst = 32'd268468224;
      4045: inst = 32'd201343955;
      4046: inst = 32'd203489279;
      4047: inst = 32'd136314880;
      4048: inst = 32'd268468224;
      4049: inst = 32'd201343956;
      4050: inst = 32'd203489279;
      4051: inst = 32'd136314880;
      4052: inst = 32'd268468224;
      4053: inst = 32'd201343957;
      4054: inst = 32'd203489279;
      4055: inst = 32'd136314880;
      4056: inst = 32'd268468224;
      4057: inst = 32'd201343958;
      4058: inst = 32'd203489279;
      4059: inst = 32'd136314880;
      4060: inst = 32'd268468224;
      4061: inst = 32'd201343959;
      4062: inst = 32'd203489279;
      4063: inst = 32'd136314880;
      4064: inst = 32'd268468224;
      4065: inst = 32'd201343960;
      4066: inst = 32'd203489279;
      4067: inst = 32'd136314880;
      4068: inst = 32'd268468224;
      4069: inst = 32'd201343961;
      4070: inst = 32'd203489279;
      4071: inst = 32'd136314880;
      4072: inst = 32'd268468224;
      4073: inst = 32'd201343962;
      4074: inst = 32'd203489279;
      4075: inst = 32'd136314880;
      4076: inst = 32'd268468224;
      4077: inst = 32'd201343963;
      4078: inst = 32'd203489279;
      4079: inst = 32'd136314880;
      4080: inst = 32'd268468224;
      4081: inst = 32'd201343964;
      4082: inst = 32'd203489279;
      4083: inst = 32'd136314880;
      4084: inst = 32'd268468224;
      4085: inst = 32'd201343965;
      4086: inst = 32'd203489279;
      4087: inst = 32'd136314880;
      4088: inst = 32'd268468224;
      4089: inst = 32'd201343966;
      4090: inst = 32'd203489279;
      4091: inst = 32'd136314880;
      4092: inst = 32'd268468224;
      4093: inst = 32'd201343967;
      4094: inst = 32'd203489279;
      4095: inst = 32'd136314880;
      4096: inst = 32'd268468224;
      4097: inst = 32'd201343968;
      4098: inst = 32'd203489279;
      4099: inst = 32'd136314880;
      4100: inst = 32'd268468224;
      4101: inst = 32'd201343969;
      4102: inst = 32'd203489279;
      4103: inst = 32'd136314880;
      4104: inst = 32'd268468224;
      4105: inst = 32'd201343970;
      4106: inst = 32'd203489279;
      4107: inst = 32'd136314880;
      4108: inst = 32'd268468224;
      4109: inst = 32'd201343971;
      4110: inst = 32'd203489278;
      4111: inst = 32'd136314880;
      4112: inst = 32'd268468224;
      4113: inst = 32'd201343972;
      4114: inst = 32'd203482808;
      4115: inst = 32'd136314880;
      4116: inst = 32'd268468224;
      4117: inst = 32'd201343973;
      4118: inst = 32'd203484855;
      4119: inst = 32'd136314880;
      4120: inst = 32'd268468224;
      4121: inst = 32'd201343974;
      4122: inst = 32'd203484855;
      4123: inst = 32'd136314880;
      4124: inst = 32'd268468224;
      4125: inst = 32'd201343975;
      4126: inst = 32'd203484854;
      4127: inst = 32'd136314880;
      4128: inst = 32'd268468224;
      4129: inst = 32'd201343976;
      4130: inst = 32'd203484854;
      4131: inst = 32'd136314880;
      4132: inst = 32'd268468224;
      4133: inst = 32'd201343977;
      4134: inst = 32'd203484854;
      4135: inst = 32'd136314880;
      4136: inst = 32'd268468224;
      4137: inst = 32'd201343978;
      4138: inst = 32'd203484854;
      4139: inst = 32'd136314880;
      4140: inst = 32'd268468224;
      4141: inst = 32'd201343979;
      4142: inst = 32'd203484854;
      4143: inst = 32'd136314880;
      4144: inst = 32'd268468224;
      4145: inst = 32'd201343980;
      4146: inst = 32'd203484854;
      4147: inst = 32'd136314880;
      4148: inst = 32'd268468224;
      4149: inst = 32'd201343981;
      4150: inst = 32'd203484854;
      4151: inst = 32'd136314880;
      4152: inst = 32'd268468224;
      4153: inst = 32'd201343982;
      4154: inst = 32'd203484854;
      4155: inst = 32'd136314880;
      4156: inst = 32'd268468224;
      4157: inst = 32'd201343983;
      4158: inst = 32'd203484854;
      4159: inst = 32'd136314880;
      4160: inst = 32'd268468224;
      4161: inst = 32'd201343984;
      4162: inst = 32'd203484853;
      4163: inst = 32'd136314880;
      4164: inst = 32'd268468224;
      4165: inst = 32'd201343985;
      4166: inst = 32'd203484854;
      4167: inst = 32'd136314880;
      4168: inst = 32'd268468224;
      4169: inst = 32'd201343986;
      4170: inst = 32'd203484854;
      4171: inst = 32'd136314880;
      4172: inst = 32'd268468224;
      4173: inst = 32'd201343987;
      4174: inst = 32'd203484854;
      4175: inst = 32'd136314880;
      4176: inst = 32'd268468224;
      4177: inst = 32'd201343988;
      4178: inst = 32'd203484854;
      4179: inst = 32'd136314880;
      4180: inst = 32'd268468224;
      4181: inst = 32'd201343989;
      4182: inst = 32'd203484854;
      4183: inst = 32'd136314880;
      4184: inst = 32'd268468224;
      4185: inst = 32'd201343990;
      4186: inst = 32'd203484854;
      4187: inst = 32'd136314880;
      4188: inst = 32'd268468224;
      4189: inst = 32'd201343991;
      4190: inst = 32'd203484822;
      4191: inst = 32'd136314880;
      4192: inst = 32'd268468224;
      4193: inst = 32'd201343992;
      4194: inst = 32'd203484854;
      4195: inst = 32'd136314880;
      4196: inst = 32'd268468224;
      4197: inst = 32'd201343993;
      4198: inst = 32'd203484854;
      4199: inst = 32'd136314880;
      4200: inst = 32'd268468224;
      4201: inst = 32'd201343994;
      4202: inst = 32'd203484854;
      4203: inst = 32'd136314880;
      4204: inst = 32'd268468224;
      4205: inst = 32'd201343995;
      4206: inst = 32'd203484854;
      4207: inst = 32'd136314880;
      4208: inst = 32'd268468224;
      4209: inst = 32'd201343996;
      4210: inst = 32'd203484854;
      4211: inst = 32'd136314880;
      4212: inst = 32'd268468224;
      4213: inst = 32'd201343997;
      4214: inst = 32'd203484854;
      4215: inst = 32'd136314880;
      4216: inst = 32'd268468224;
      4217: inst = 32'd201343998;
      4218: inst = 32'd203484854;
      4219: inst = 32'd136314880;
      4220: inst = 32'd268468224;
      4221: inst = 32'd201343999;
      4222: inst = 32'd203484854;
      4223: inst = 32'd136314880;
      4224: inst = 32'd268468224;
      4225: inst = 32'd201344000;
      4226: inst = 32'd203486934;
      4227: inst = 32'd136314880;
      4228: inst = 32'd268468224;
      4229: inst = 32'd201344001;
      4230: inst = 32'd203484854;
      4231: inst = 32'd136314880;
      4232: inst = 32'd268468224;
      4233: inst = 32'd201344002;
      4234: inst = 32'd203482773;
      4235: inst = 32'd136314880;
      4236: inst = 32'd268468224;
      4237: inst = 32'd201344003;
      4238: inst = 32'd203482806;
      4239: inst = 32'd136314880;
      4240: inst = 32'd268468224;
      4241: inst = 32'd201344004;
      4242: inst = 32'd203484951;
      4243: inst = 32'd136314880;
      4244: inst = 32'd268468224;
      4245: inst = 32'd201344005;
      4246: inst = 32'd203484886;
      4247: inst = 32'd136314880;
      4248: inst = 32'd268468224;
      4249: inst = 32'd201344006;
      4250: inst = 32'd203476304;
      4251: inst = 32'd136314880;
      4252: inst = 32'd268468224;
      4253: inst = 32'd201344007;
      4254: inst = 32'd203467722;
      4255: inst = 32'd136314880;
      4256: inst = 32'd268468224;
      4257: inst = 32'd201344008;
      4258: inst = 32'd203467527;
      4259: inst = 32'd136314880;
      4260: inst = 32'd268468224;
      4261: inst = 32'd201344009;
      4262: inst = 32'd203473704;
      4263: inst = 32'd136314880;
      4264: inst = 32'd268468224;
      4265: inst = 32'd201344010;
      4266: inst = 32'd203473639;
      4267: inst = 32'd136314880;
      4268: inst = 32'd268468224;
      4269: inst = 32'd201344011;
      4270: inst = 32'd203475655;
      4271: inst = 32'd136314880;
      4272: inst = 32'd268468224;
      4273: inst = 32'd201344012;
      4274: inst = 32'd203473607;
      4275: inst = 32'd136314880;
      4276: inst = 32'd268468224;
      4277: inst = 32'd201344013;
      4278: inst = 32'd203473639;
      4279: inst = 32'd136314880;
      4280: inst = 32'd268468224;
      4281: inst = 32'd201344014;
      4282: inst = 32'd203473672;
      4283: inst = 32'd136314880;
      4284: inst = 32'd268468224;
      4285: inst = 32'd201344015;
      4286: inst = 32'd203469511;
      4287: inst = 32'd136314880;
      4288: inst = 32'd268468224;
      4289: inst = 32'd201344016;
      4290: inst = 32'd203463660;
      4291: inst = 32'd136314880;
      4292: inst = 32'd268468224;
      4293: inst = 32'd201344017;
      4294: inst = 32'd203476305;
      4295: inst = 32'd136314880;
      4296: inst = 32'd268468224;
      4297: inst = 32'd201344018;
      4298: inst = 32'd203486902;
      4299: inst = 32'd136314880;
      4300: inst = 32'd268468224;
      4301: inst = 32'd201344019;
      4302: inst = 32'd203486967;
      4303: inst = 32'd136314880;
      4304: inst = 32'd268468224;
      4305: inst = 32'd201344020;
      4306: inst = 32'd203484822;
      4307: inst = 32'd136314880;
      4308: inst = 32'd268468224;
      4309: inst = 32'd201344021;
      4310: inst = 32'd203482773;
      4311: inst = 32'd136314880;
      4312: inst = 32'd268468224;
      4313: inst = 32'd201344022;
      4314: inst = 32'd203484854;
      4315: inst = 32'd136314880;
      4316: inst = 32'd268468224;
      4317: inst = 32'd201344023;
      4318: inst = 32'd203484887;
      4319: inst = 32'd136314880;
      4320: inst = 32'd268468224;
      4321: inst = 32'd201344024;
      4322: inst = 32'd203484854;
      4323: inst = 32'd136314880;
      4324: inst = 32'd268468224;
      4325: inst = 32'd201344025;
      4326: inst = 32'd203484855;
      4327: inst = 32'd136314880;
      4328: inst = 32'd268468224;
      4329: inst = 32'd201344026;
      4330: inst = 32'd203484887;
      4331: inst = 32'd136314880;
      4332: inst = 32'd268468224;
      4333: inst = 32'd201344027;
      4334: inst = 32'd203482808;
      4335: inst = 32'd136314880;
      4336: inst = 32'd268468224;
      4337: inst = 32'd201344028;
      4338: inst = 32'd203489278;
      4339: inst = 32'd136314880;
      4340: inst = 32'd268468224;
      4341: inst = 32'd201344029;
      4342: inst = 32'd203489279;
      4343: inst = 32'd136314880;
      4344: inst = 32'd268468224;
      4345: inst = 32'd201344030;
      4346: inst = 32'd203489279;
      4347: inst = 32'd136314880;
      4348: inst = 32'd268468224;
      4349: inst = 32'd201344031;
      4350: inst = 32'd203489279;
      4351: inst = 32'd136314880;
      4352: inst = 32'd268468224;
      4353: inst = 32'd201344032;
      4354: inst = 32'd203489279;
      4355: inst = 32'd136314880;
      4356: inst = 32'd268468224;
      4357: inst = 32'd201344033;
      4358: inst = 32'd203489279;
      4359: inst = 32'd136314880;
      4360: inst = 32'd268468224;
      4361: inst = 32'd201344034;
      4362: inst = 32'd203489279;
      4363: inst = 32'd136314880;
      4364: inst = 32'd268468224;
      4365: inst = 32'd201344035;
      4366: inst = 32'd203489279;
      4367: inst = 32'd136314880;
      4368: inst = 32'd268468224;
      4369: inst = 32'd201344036;
      4370: inst = 32'd203489279;
      4371: inst = 32'd136314880;
      4372: inst = 32'd268468224;
      4373: inst = 32'd201344037;
      4374: inst = 32'd203489279;
      4375: inst = 32'd136314880;
      4376: inst = 32'd268468224;
      4377: inst = 32'd201344038;
      4378: inst = 32'd203489279;
      4379: inst = 32'd136314880;
      4380: inst = 32'd268468224;
      4381: inst = 32'd201344039;
      4382: inst = 32'd203489279;
      4383: inst = 32'd136314880;
      4384: inst = 32'd268468224;
      4385: inst = 32'd201344040;
      4386: inst = 32'd203489279;
      4387: inst = 32'd136314880;
      4388: inst = 32'd268468224;
      4389: inst = 32'd201344041;
      4390: inst = 32'd203489279;
      4391: inst = 32'd136314880;
      4392: inst = 32'd268468224;
      4393: inst = 32'd201344042;
      4394: inst = 32'd203489279;
      4395: inst = 32'd136314880;
      4396: inst = 32'd268468224;
      4397: inst = 32'd201344043;
      4398: inst = 32'd203489279;
      4399: inst = 32'd136314880;
      4400: inst = 32'd268468224;
      4401: inst = 32'd201344044;
      4402: inst = 32'd203489279;
      4403: inst = 32'd136314880;
      4404: inst = 32'd268468224;
      4405: inst = 32'd201344045;
      4406: inst = 32'd203489279;
      4407: inst = 32'd136314880;
      4408: inst = 32'd268468224;
      4409: inst = 32'd201344046;
      4410: inst = 32'd203489279;
      4411: inst = 32'd136314880;
      4412: inst = 32'd268468224;
      4413: inst = 32'd201344047;
      4414: inst = 32'd203489279;
      4415: inst = 32'd136314880;
      4416: inst = 32'd268468224;
      4417: inst = 32'd201344048;
      4418: inst = 32'd203489279;
      4419: inst = 32'd136314880;
      4420: inst = 32'd268468224;
      4421: inst = 32'd201344049;
      4422: inst = 32'd203489279;
      4423: inst = 32'd136314880;
      4424: inst = 32'd268468224;
      4425: inst = 32'd201344050;
      4426: inst = 32'd203489279;
      4427: inst = 32'd136314880;
      4428: inst = 32'd268468224;
      4429: inst = 32'd201344051;
      4430: inst = 32'd203489279;
      4431: inst = 32'd136314880;
      4432: inst = 32'd268468224;
      4433: inst = 32'd201344052;
      4434: inst = 32'd203489279;
      4435: inst = 32'd136314880;
      4436: inst = 32'd268468224;
      4437: inst = 32'd201344053;
      4438: inst = 32'd203489279;
      4439: inst = 32'd136314880;
      4440: inst = 32'd268468224;
      4441: inst = 32'd201344054;
      4442: inst = 32'd203489279;
      4443: inst = 32'd136314880;
      4444: inst = 32'd268468224;
      4445: inst = 32'd201344055;
      4446: inst = 32'd203489279;
      4447: inst = 32'd136314880;
      4448: inst = 32'd268468224;
      4449: inst = 32'd201344056;
      4450: inst = 32'd203489279;
      4451: inst = 32'd136314880;
      4452: inst = 32'd268468224;
      4453: inst = 32'd201344057;
      4454: inst = 32'd203489279;
      4455: inst = 32'd136314880;
      4456: inst = 32'd268468224;
      4457: inst = 32'd201344058;
      4458: inst = 32'd203489279;
      4459: inst = 32'd136314880;
      4460: inst = 32'd268468224;
      4461: inst = 32'd201344059;
      4462: inst = 32'd203489279;
      4463: inst = 32'd136314880;
      4464: inst = 32'd268468224;
      4465: inst = 32'd201344060;
      4466: inst = 32'd203489279;
      4467: inst = 32'd136314880;
      4468: inst = 32'd268468224;
      4469: inst = 32'd201344061;
      4470: inst = 32'd203489279;
      4471: inst = 32'd136314880;
      4472: inst = 32'd268468224;
      4473: inst = 32'd201344062;
      4474: inst = 32'd203489279;
      4475: inst = 32'd136314880;
      4476: inst = 32'd268468224;
      4477: inst = 32'd201344063;
      4478: inst = 32'd203489279;
      4479: inst = 32'd136314880;
      4480: inst = 32'd268468224;
      4481: inst = 32'd201344064;
      4482: inst = 32'd203489279;
      4483: inst = 32'd136314880;
      4484: inst = 32'd268468224;
      4485: inst = 32'd201344065;
      4486: inst = 32'd203489279;
      4487: inst = 32'd136314880;
      4488: inst = 32'd268468224;
      4489: inst = 32'd201344066;
      4490: inst = 32'd203489279;
      4491: inst = 32'd136314880;
      4492: inst = 32'd268468224;
      4493: inst = 32'd201344067;
      4494: inst = 32'd203489278;
      4495: inst = 32'd136314880;
      4496: inst = 32'd268468224;
      4497: inst = 32'd201344068;
      4498: inst = 32'd203482808;
      4499: inst = 32'd136314880;
      4500: inst = 32'd268468224;
      4501: inst = 32'd201344069;
      4502: inst = 32'd203484855;
      4503: inst = 32'd136314880;
      4504: inst = 32'd268468224;
      4505: inst = 32'd201344070;
      4506: inst = 32'd203484855;
      4507: inst = 32'd136314880;
      4508: inst = 32'd268468224;
      4509: inst = 32'd201344071;
      4510: inst = 32'd203484854;
      4511: inst = 32'd136314880;
      4512: inst = 32'd268468224;
      4513: inst = 32'd201344072;
      4514: inst = 32'd203484854;
      4515: inst = 32'd136314880;
      4516: inst = 32'd268468224;
      4517: inst = 32'd201344073;
      4518: inst = 32'd203484854;
      4519: inst = 32'd136314880;
      4520: inst = 32'd268468224;
      4521: inst = 32'd201344074;
      4522: inst = 32'd203484854;
      4523: inst = 32'd136314880;
      4524: inst = 32'd268468224;
      4525: inst = 32'd201344075;
      4526: inst = 32'd203484854;
      4527: inst = 32'd136314880;
      4528: inst = 32'd268468224;
      4529: inst = 32'd201344076;
      4530: inst = 32'd203484854;
      4531: inst = 32'd136314880;
      4532: inst = 32'd268468224;
      4533: inst = 32'd201344077;
      4534: inst = 32'd203484854;
      4535: inst = 32'd136314880;
      4536: inst = 32'd268468224;
      4537: inst = 32'd201344078;
      4538: inst = 32'd203484854;
      4539: inst = 32'd136314880;
      4540: inst = 32'd268468224;
      4541: inst = 32'd201344079;
      4542: inst = 32'd203484854;
      4543: inst = 32'd136314880;
      4544: inst = 32'd268468224;
      4545: inst = 32'd201344080;
      4546: inst = 32'd203486934;
      4547: inst = 32'd136314880;
      4548: inst = 32'd268468224;
      4549: inst = 32'd201344081;
      4550: inst = 32'd203486934;
      4551: inst = 32'd136314880;
      4552: inst = 32'd268468224;
      4553: inst = 32'd201344082;
      4554: inst = 32'd203484886;
      4555: inst = 32'd136314880;
      4556: inst = 32'd268468224;
      4557: inst = 32'd201344083;
      4558: inst = 32'd203484854;
      4559: inst = 32'd136314880;
      4560: inst = 32'd268468224;
      4561: inst = 32'd201344084;
      4562: inst = 32'd203484854;
      4563: inst = 32'd136314880;
      4564: inst = 32'd268468224;
      4565: inst = 32'd201344085;
      4566: inst = 32'd203484886;
      4567: inst = 32'd136314880;
      4568: inst = 32'd268468224;
      4569: inst = 32'd201344086;
      4570: inst = 32'd203486934;
      4571: inst = 32'd136314880;
      4572: inst = 32'd268468224;
      4573: inst = 32'd201344087;
      4574: inst = 32'd203486935;
      4575: inst = 32'd136314880;
      4576: inst = 32'd268468224;
      4577: inst = 32'd201344088;
      4578: inst = 32'd203484854;
      4579: inst = 32'd136314880;
      4580: inst = 32'd268468224;
      4581: inst = 32'd201344089;
      4582: inst = 32'd203484854;
      4583: inst = 32'd136314880;
      4584: inst = 32'd268468224;
      4585: inst = 32'd201344090;
      4586: inst = 32'd203484854;
      4587: inst = 32'd136314880;
      4588: inst = 32'd268468224;
      4589: inst = 32'd201344091;
      4590: inst = 32'd203484854;
      4591: inst = 32'd136314880;
      4592: inst = 32'd268468224;
      4593: inst = 32'd201344092;
      4594: inst = 32'd203484854;
      4595: inst = 32'd136314880;
      4596: inst = 32'd268468224;
      4597: inst = 32'd201344093;
      4598: inst = 32'd203484854;
      4599: inst = 32'd136314880;
      4600: inst = 32'd268468224;
      4601: inst = 32'd201344094;
      4602: inst = 32'd203484854;
      4603: inst = 32'd136314880;
      4604: inst = 32'd268468224;
      4605: inst = 32'd201344095;
      4606: inst = 32'd203484854;
      4607: inst = 32'd136314880;
      4608: inst = 32'd268468224;
      4609: inst = 32'd201344096;
      4610: inst = 32'd203486837;
      4611: inst = 32'd136314880;
      4612: inst = 32'd268468224;
      4613: inst = 32'd201344097;
      4614: inst = 32'd203486902;
      4615: inst = 32'd136314880;
      4616: inst = 32'd268468224;
      4617: inst = 32'd201344098;
      4618: inst = 32'd203486934;
      4619: inst = 32'd136314880;
      4620: inst = 32'd268468224;
      4621: inst = 32'd201344099;
      4622: inst = 32'd203484886;
      4623: inst = 32'd136314880;
      4624: inst = 32'd268468224;
      4625: inst = 32'd201344100;
      4626: inst = 32'd203482806;
      4627: inst = 32'd136314880;
      4628: inst = 32'd268468224;
      4629: inst = 32'd201344101;
      4630: inst = 32'd203482806;
      4631: inst = 32'd136314880;
      4632: inst = 32'd268468224;
      4633: inst = 32'd201344102;
      4634: inst = 32'd203484854;
      4635: inst = 32'd136314880;
      4636: inst = 32'd268468224;
      4637: inst = 32'd201344103;
      4638: inst = 32'd203486869;
      4639: inst = 32'd136314880;
      4640: inst = 32'd268468224;
      4641: inst = 32'd201344104;
      4642: inst = 32'd203488884;
      4643: inst = 32'd136314880;
      4644: inst = 32'd268468224;
      4645: inst = 32'd201344105;
      4646: inst = 32'd203488852;
      4647: inst = 32'd136314880;
      4648: inst = 32'd268468224;
      4649: inst = 32'd201344106;
      4650: inst = 32'd203488722;
      4651: inst = 32'd136314880;
      4652: inst = 32'd268468224;
      4653: inst = 32'd201344107;
      4654: inst = 32'd203488689;
      4655: inst = 32'd136314880;
      4656: inst = 32'd268468224;
      4657: inst = 32'd201344108;
      4658: inst = 32'd203488722;
      4659: inst = 32'd136314880;
      4660: inst = 32'd268468224;
      4661: inst = 32'd201344109;
      4662: inst = 32'd203488754;
      4663: inst = 32'd136314880;
      4664: inst = 32'd268468224;
      4665: inst = 32'd201344110;
      4666: inst = 32'd203488884;
      4667: inst = 32'd136314880;
      4668: inst = 32'd268468224;
      4669: inst = 32'd201344111;
      4670: inst = 32'd203488884;
      4671: inst = 32'd136314880;
      4672: inst = 32'd268468224;
      4673: inst = 32'd201344112;
      4674: inst = 32'd203484822;
      4675: inst = 32'd136314880;
      4676: inst = 32'd268468224;
      4677: inst = 32'd201344113;
      4678: inst = 32'd203484822;
      4679: inst = 32'd136314880;
      4680: inst = 32'd268468224;
      4681: inst = 32'd201344114;
      4682: inst = 32'd203484822;
      4683: inst = 32'd136314880;
      4684: inst = 32'd268468224;
      4685: inst = 32'd201344115;
      4686: inst = 32'd203484822;
      4687: inst = 32'd136314880;
      4688: inst = 32'd268468224;
      4689: inst = 32'd201344116;
      4690: inst = 32'd203484854;
      4691: inst = 32'd136314880;
      4692: inst = 32'd268468224;
      4693: inst = 32'd201344117;
      4694: inst = 32'd203486934;
      4695: inst = 32'd136314880;
      4696: inst = 32'd268468224;
      4697: inst = 32'd201344118;
      4698: inst = 32'd203484886;
      4699: inst = 32'd136314880;
      4700: inst = 32'd268468224;
      4701: inst = 32'd201344119;
      4702: inst = 32'd203484821;
      4703: inst = 32'd136314880;
      4704: inst = 32'd268468224;
      4705: inst = 32'd201344120;
      4706: inst = 32'd203484854;
      4707: inst = 32'd136314880;
      4708: inst = 32'd268468224;
      4709: inst = 32'd201344121;
      4710: inst = 32'd203484854;
      4711: inst = 32'd136314880;
      4712: inst = 32'd268468224;
      4713: inst = 32'd201344122;
      4714: inst = 32'd203484887;
      4715: inst = 32'd136314880;
      4716: inst = 32'd268468224;
      4717: inst = 32'd201344123;
      4718: inst = 32'd203482808;
      4719: inst = 32'd136314880;
      4720: inst = 32'd268468224;
      4721: inst = 32'd201344124;
      4722: inst = 32'd203489278;
      4723: inst = 32'd136314880;
      4724: inst = 32'd268468224;
      4725: inst = 32'd201344125;
      4726: inst = 32'd203489279;
      4727: inst = 32'd136314880;
      4728: inst = 32'd268468224;
      4729: inst = 32'd201344126;
      4730: inst = 32'd203489279;
      4731: inst = 32'd136314880;
      4732: inst = 32'd268468224;
      4733: inst = 32'd201344127;
      4734: inst = 32'd203489279;
      4735: inst = 32'd136314880;
      4736: inst = 32'd268468224;
      4737: inst = 32'd201344128;
      4738: inst = 32'd203489279;
      4739: inst = 32'd136314880;
      4740: inst = 32'd268468224;
      4741: inst = 32'd201344129;
      4742: inst = 32'd203489279;
      4743: inst = 32'd136314880;
      4744: inst = 32'd268468224;
      4745: inst = 32'd201344130;
      4746: inst = 32'd203489279;
      4747: inst = 32'd136314880;
      4748: inst = 32'd268468224;
      4749: inst = 32'd201344131;
      4750: inst = 32'd203489279;
      4751: inst = 32'd136314880;
      4752: inst = 32'd268468224;
      4753: inst = 32'd201344132;
      4754: inst = 32'd203489279;
      4755: inst = 32'd136314880;
      4756: inst = 32'd268468224;
      4757: inst = 32'd201344133;
      4758: inst = 32'd203489279;
      4759: inst = 32'd136314880;
      4760: inst = 32'd268468224;
      4761: inst = 32'd201344134;
      4762: inst = 32'd203489279;
      4763: inst = 32'd136314880;
      4764: inst = 32'd268468224;
      4765: inst = 32'd201344135;
      4766: inst = 32'd203489279;
      4767: inst = 32'd136314880;
      4768: inst = 32'd268468224;
      4769: inst = 32'd201344136;
      4770: inst = 32'd203489279;
      4771: inst = 32'd136314880;
      4772: inst = 32'd268468224;
      4773: inst = 32'd201344137;
      4774: inst = 32'd203489279;
      4775: inst = 32'd136314880;
      4776: inst = 32'd268468224;
      4777: inst = 32'd201344138;
      4778: inst = 32'd203489279;
      4779: inst = 32'd136314880;
      4780: inst = 32'd268468224;
      4781: inst = 32'd201344139;
      4782: inst = 32'd203489279;
      4783: inst = 32'd136314880;
      4784: inst = 32'd268468224;
      4785: inst = 32'd201344140;
      4786: inst = 32'd203489279;
      4787: inst = 32'd136314880;
      4788: inst = 32'd268468224;
      4789: inst = 32'd201344141;
      4790: inst = 32'd203489279;
      4791: inst = 32'd136314880;
      4792: inst = 32'd268468224;
      4793: inst = 32'd201344142;
      4794: inst = 32'd203489279;
      4795: inst = 32'd136314880;
      4796: inst = 32'd268468224;
      4797: inst = 32'd201344143;
      4798: inst = 32'd203489279;
      4799: inst = 32'd136314880;
      4800: inst = 32'd268468224;
      4801: inst = 32'd201344144;
      4802: inst = 32'd203489279;
      4803: inst = 32'd136314880;
      4804: inst = 32'd268468224;
      4805: inst = 32'd201344145;
      4806: inst = 32'd203489279;
      4807: inst = 32'd136314880;
      4808: inst = 32'd268468224;
      4809: inst = 32'd201344146;
      4810: inst = 32'd203489279;
      4811: inst = 32'd136314880;
      4812: inst = 32'd268468224;
      4813: inst = 32'd201344147;
      4814: inst = 32'd203489279;
      4815: inst = 32'd136314880;
      4816: inst = 32'd268468224;
      4817: inst = 32'd201344148;
      4818: inst = 32'd203489279;
      4819: inst = 32'd136314880;
      4820: inst = 32'd268468224;
      4821: inst = 32'd201344149;
      4822: inst = 32'd203489279;
      4823: inst = 32'd136314880;
      4824: inst = 32'd268468224;
      4825: inst = 32'd201344150;
      4826: inst = 32'd203489279;
      4827: inst = 32'd136314880;
      4828: inst = 32'd268468224;
      4829: inst = 32'd201344151;
      4830: inst = 32'd203489279;
      4831: inst = 32'd136314880;
      4832: inst = 32'd268468224;
      4833: inst = 32'd201344152;
      4834: inst = 32'd203489279;
      4835: inst = 32'd136314880;
      4836: inst = 32'd268468224;
      4837: inst = 32'd201344153;
      4838: inst = 32'd203489279;
      4839: inst = 32'd136314880;
      4840: inst = 32'd268468224;
      4841: inst = 32'd201344154;
      4842: inst = 32'd203489279;
      4843: inst = 32'd136314880;
      4844: inst = 32'd268468224;
      4845: inst = 32'd201344155;
      4846: inst = 32'd203489279;
      4847: inst = 32'd136314880;
      4848: inst = 32'd268468224;
      4849: inst = 32'd201344156;
      4850: inst = 32'd203489279;
      4851: inst = 32'd136314880;
      4852: inst = 32'd268468224;
      4853: inst = 32'd201344157;
      4854: inst = 32'd203489279;
      4855: inst = 32'd136314880;
      4856: inst = 32'd268468224;
      4857: inst = 32'd201344158;
      4858: inst = 32'd203489279;
      4859: inst = 32'd136314880;
      4860: inst = 32'd268468224;
      4861: inst = 32'd201344159;
      4862: inst = 32'd203489279;
      4863: inst = 32'd136314880;
      4864: inst = 32'd268468224;
      4865: inst = 32'd201344160;
      4866: inst = 32'd203489279;
      4867: inst = 32'd136314880;
      4868: inst = 32'd268468224;
      4869: inst = 32'd201344161;
      4870: inst = 32'd203489279;
      4871: inst = 32'd136314880;
      4872: inst = 32'd268468224;
      4873: inst = 32'd201344162;
      4874: inst = 32'd203489279;
      4875: inst = 32'd136314880;
      4876: inst = 32'd268468224;
      4877: inst = 32'd201344163;
      4878: inst = 32'd203489278;
      4879: inst = 32'd136314880;
      4880: inst = 32'd268468224;
      4881: inst = 32'd201344164;
      4882: inst = 32'd203482808;
      4883: inst = 32'd136314880;
      4884: inst = 32'd268468224;
      4885: inst = 32'd201344165;
      4886: inst = 32'd203484855;
      4887: inst = 32'd136314880;
      4888: inst = 32'd268468224;
      4889: inst = 32'd201344166;
      4890: inst = 32'd203484854;
      4891: inst = 32'd136314880;
      4892: inst = 32'd268468224;
      4893: inst = 32'd201344167;
      4894: inst = 32'd203484854;
      4895: inst = 32'd136314880;
      4896: inst = 32'd268468224;
      4897: inst = 32'd201344168;
      4898: inst = 32'd203484854;
      4899: inst = 32'd136314880;
      4900: inst = 32'd268468224;
      4901: inst = 32'd201344169;
      4902: inst = 32'd203484854;
      4903: inst = 32'd136314880;
      4904: inst = 32'd268468224;
      4905: inst = 32'd201344170;
      4906: inst = 32'd203484854;
      4907: inst = 32'd136314880;
      4908: inst = 32'd268468224;
      4909: inst = 32'd201344171;
      4910: inst = 32'd203484854;
      4911: inst = 32'd136314880;
      4912: inst = 32'd268468224;
      4913: inst = 32'd201344172;
      4914: inst = 32'd203484854;
      4915: inst = 32'd136314880;
      4916: inst = 32'd268468224;
      4917: inst = 32'd201344173;
      4918: inst = 32'd203484854;
      4919: inst = 32'd136314880;
      4920: inst = 32'd268468224;
      4921: inst = 32'd201344174;
      4922: inst = 32'd203484854;
      4923: inst = 32'd136314880;
      4924: inst = 32'd268468224;
      4925: inst = 32'd201344175;
      4926: inst = 32'd203484854;
      4927: inst = 32'd136314880;
      4928: inst = 32'd268468224;
      4929: inst = 32'd201344176;
      4930: inst = 32'd203484886;
      4931: inst = 32'd136314880;
      4932: inst = 32'd268468224;
      4933: inst = 32'd201344177;
      4934: inst = 32'd203484821;
      4935: inst = 32'd136314880;
      4936: inst = 32'd268468224;
      4937: inst = 32'd201344178;
      4938: inst = 32'd203482708;
      4939: inst = 32'd136314880;
      4940: inst = 32'd268468224;
      4941: inst = 32'd201344179;
      4942: inst = 32'd203480627;
      4943: inst = 32'd136314880;
      4944: inst = 32'd268468224;
      4945: inst = 32'd201344180;
      4946: inst = 32'd203480628;
      4947: inst = 32'd136314880;
      4948: inst = 32'd268468224;
      4949: inst = 32'd201344181;
      4950: inst = 32'd203482708;
      4951: inst = 32'd136314880;
      4952: inst = 32'd268468224;
      4953: inst = 32'd201344182;
      4954: inst = 32'd203484821;
      4955: inst = 32'd136314880;
      4956: inst = 32'd268468224;
      4957: inst = 32'd201344183;
      4958: inst = 32'd203484854;
      4959: inst = 32'd136314880;
      4960: inst = 32'd268468224;
      4961: inst = 32'd201344184;
      4962: inst = 32'd203484854;
      4963: inst = 32'd136314880;
      4964: inst = 32'd268468224;
      4965: inst = 32'd201344185;
      4966: inst = 32'd203484854;
      4967: inst = 32'd136314880;
      4968: inst = 32'd268468224;
      4969: inst = 32'd201344186;
      4970: inst = 32'd203484854;
      4971: inst = 32'd136314880;
      4972: inst = 32'd268468224;
      4973: inst = 32'd201344187;
      4974: inst = 32'd203484854;
      4975: inst = 32'd136314880;
      4976: inst = 32'd268468224;
      4977: inst = 32'd201344188;
      4978: inst = 32'd203484854;
      4979: inst = 32'd136314880;
      4980: inst = 32'd268468224;
      4981: inst = 32'd201344189;
      4982: inst = 32'd203484854;
      4983: inst = 32'd136314880;
      4984: inst = 32'd268468224;
      4985: inst = 32'd201344190;
      4986: inst = 32'd203484854;
      4987: inst = 32'd136314880;
      4988: inst = 32'd268468224;
      4989: inst = 32'd201344191;
      4990: inst = 32'd203484854;
      4991: inst = 32'd136314880;
      4992: inst = 32'd268468224;
      4993: inst = 32'd201344192;
      4994: inst = 32'd203486901;
      4995: inst = 32'd136314880;
      4996: inst = 32'd268468224;
      4997: inst = 32'd201344193;
      4998: inst = 32'd203484821;
      4999: inst = 32'd136314880;
      5000: inst = 32'd268468224;
      5001: inst = 32'd201344194;
      5002: inst = 32'd203484854;
      5003: inst = 32'd136314880;
      5004: inst = 32'd268468224;
      5005: inst = 32'd201344195;
      5006: inst = 32'd203484887;
      5007: inst = 32'd136314880;
      5008: inst = 32'd268468224;
      5009: inst = 32'd201344196;
      5010: inst = 32'd203484920;
      5011: inst = 32'd136314880;
      5012: inst = 32'd268468224;
      5013: inst = 32'd201344197;
      5014: inst = 32'd203484919;
      5015: inst = 32'd136314880;
      5016: inst = 32'd268468224;
      5017: inst = 32'd201344198;
      5018: inst = 32'd203484886;
      5019: inst = 32'd136314880;
      5020: inst = 32'd268468224;
      5021: inst = 32'd201344199;
      5022: inst = 32'd203484854;
      5023: inst = 32'd136314880;
      5024: inst = 32'd268468224;
      5025: inst = 32'd201344200;
      5026: inst = 32'd203486934;
      5027: inst = 32'd136314880;
      5028: inst = 32'd268468224;
      5029: inst = 32'd201344201;
      5030: inst = 32'd203484787;
      5031: inst = 32'd136314880;
      5032: inst = 32'd268468224;
      5033: inst = 32'd201344202;
      5034: inst = 32'd203488981;
      5035: inst = 32'd136314880;
      5036: inst = 32'd268468224;
      5037: inst = 32'd201344203;
      5038: inst = 32'd203486868;
      5039: inst = 32'd136314880;
      5040: inst = 32'd268468224;
      5041: inst = 32'd201344204;
      5042: inst = 32'd203486868;
      5043: inst = 32'd136314880;
      5044: inst = 32'd268468224;
      5045: inst = 32'd201344205;
      5046: inst = 32'd203486933;
      5047: inst = 32'd136314880;
      5048: inst = 32'd268468224;
      5049: inst = 32'd201344206;
      5050: inst = 32'd203482772;
      5051: inst = 32'd136314880;
      5052: inst = 32'd268468224;
      5053: inst = 32'd201344207;
      5054: inst = 32'd203486966;
      5055: inst = 32'd136314880;
      5056: inst = 32'd268468224;
      5057: inst = 32'd201344208;
      5058: inst = 32'd203486870;
      5059: inst = 32'd136314880;
      5060: inst = 32'd268468224;
      5061: inst = 32'd201344209;
      5062: inst = 32'd203486903;
      5063: inst = 32'd136314880;
      5064: inst = 32'd268468224;
      5065: inst = 32'd201344210;
      5066: inst = 32'd203486935;
      5067: inst = 32'd136314880;
      5068: inst = 32'd268468224;
      5069: inst = 32'd201344211;
      5070: inst = 32'd203486967;
      5071: inst = 32'd136314880;
      5072: inst = 32'd268468224;
      5073: inst = 32'd201344212;
      5074: inst = 32'd203486935;
      5075: inst = 32'd136314880;
      5076: inst = 32'd268468224;
      5077: inst = 32'd201344213;
      5078: inst = 32'd203484854;
      5079: inst = 32'd136314880;
      5080: inst = 32'd268468224;
      5081: inst = 32'd201344214;
      5082: inst = 32'd203484853;
      5083: inst = 32'd136314880;
      5084: inst = 32'd268468224;
      5085: inst = 32'd201344215;
      5086: inst = 32'd203484854;
      5087: inst = 32'd136314880;
      5088: inst = 32'd268468224;
      5089: inst = 32'd201344216;
      5090: inst = 32'd203484854;
      5091: inst = 32'd136314880;
      5092: inst = 32'd268468224;
      5093: inst = 32'd201344217;
      5094: inst = 32'd203484854;
      5095: inst = 32'd136314880;
      5096: inst = 32'd268468224;
      5097: inst = 32'd201344218;
      5098: inst = 32'd203484887;
      5099: inst = 32'd136314880;
      5100: inst = 32'd268468224;
      5101: inst = 32'd201344219;
      5102: inst = 32'd203482840;
      5103: inst = 32'd136314880;
      5104: inst = 32'd268468224;
      5105: inst = 32'd201344220;
      5106: inst = 32'd203489278;
      5107: inst = 32'd136314880;
      5108: inst = 32'd268468224;
      5109: inst = 32'd201344221;
      5110: inst = 32'd203489279;
      5111: inst = 32'd136314880;
      5112: inst = 32'd268468224;
      5113: inst = 32'd201344222;
      5114: inst = 32'd203489279;
      5115: inst = 32'd136314880;
      5116: inst = 32'd268468224;
      5117: inst = 32'd201344223;
      5118: inst = 32'd203489279;
      5119: inst = 32'd136314880;
      5120: inst = 32'd268468224;
      5121: inst = 32'd201344224;
      5122: inst = 32'd203489279;
      5123: inst = 32'd136314880;
      5124: inst = 32'd268468224;
      5125: inst = 32'd201344225;
      5126: inst = 32'd203489279;
      5127: inst = 32'd136314880;
      5128: inst = 32'd268468224;
      5129: inst = 32'd201344226;
      5130: inst = 32'd203489279;
      5131: inst = 32'd136314880;
      5132: inst = 32'd268468224;
      5133: inst = 32'd201344227;
      5134: inst = 32'd203489279;
      5135: inst = 32'd136314880;
      5136: inst = 32'd268468224;
      5137: inst = 32'd201344228;
      5138: inst = 32'd203489279;
      5139: inst = 32'd136314880;
      5140: inst = 32'd268468224;
      5141: inst = 32'd201344229;
      5142: inst = 32'd203489279;
      5143: inst = 32'd136314880;
      5144: inst = 32'd268468224;
      5145: inst = 32'd201344230;
      5146: inst = 32'd203489279;
      5147: inst = 32'd136314880;
      5148: inst = 32'd268468224;
      5149: inst = 32'd201344231;
      5150: inst = 32'd203489279;
      5151: inst = 32'd136314880;
      5152: inst = 32'd268468224;
      5153: inst = 32'd201344232;
      5154: inst = 32'd203489279;
      5155: inst = 32'd136314880;
      5156: inst = 32'd268468224;
      5157: inst = 32'd201344233;
      5158: inst = 32'd203489279;
      5159: inst = 32'd136314880;
      5160: inst = 32'd268468224;
      5161: inst = 32'd201344234;
      5162: inst = 32'd203489279;
      5163: inst = 32'd136314880;
      5164: inst = 32'd268468224;
      5165: inst = 32'd201344235;
      5166: inst = 32'd203489279;
      5167: inst = 32'd136314880;
      5168: inst = 32'd268468224;
      5169: inst = 32'd201344236;
      5170: inst = 32'd203489279;
      5171: inst = 32'd136314880;
      5172: inst = 32'd268468224;
      5173: inst = 32'd201344237;
      5174: inst = 32'd203489279;
      5175: inst = 32'd136314880;
      5176: inst = 32'd268468224;
      5177: inst = 32'd201344238;
      5178: inst = 32'd203489279;
      5179: inst = 32'd136314880;
      5180: inst = 32'd268468224;
      5181: inst = 32'd201344239;
      5182: inst = 32'd203489279;
      5183: inst = 32'd136314880;
      5184: inst = 32'd268468224;
      5185: inst = 32'd201344240;
      5186: inst = 32'd203489279;
      5187: inst = 32'd136314880;
      5188: inst = 32'd268468224;
      5189: inst = 32'd201344241;
      5190: inst = 32'd203489279;
      5191: inst = 32'd136314880;
      5192: inst = 32'd268468224;
      5193: inst = 32'd201344242;
      5194: inst = 32'd203489279;
      5195: inst = 32'd136314880;
      5196: inst = 32'd268468224;
      5197: inst = 32'd201344243;
      5198: inst = 32'd203489279;
      5199: inst = 32'd136314880;
      5200: inst = 32'd268468224;
      5201: inst = 32'd201344244;
      5202: inst = 32'd203489279;
      5203: inst = 32'd136314880;
      5204: inst = 32'd268468224;
      5205: inst = 32'd201344245;
      5206: inst = 32'd203489279;
      5207: inst = 32'd136314880;
      5208: inst = 32'd268468224;
      5209: inst = 32'd201344246;
      5210: inst = 32'd203489279;
      5211: inst = 32'd136314880;
      5212: inst = 32'd268468224;
      5213: inst = 32'd201344247;
      5214: inst = 32'd203489279;
      5215: inst = 32'd136314880;
      5216: inst = 32'd268468224;
      5217: inst = 32'd201344248;
      5218: inst = 32'd203489279;
      5219: inst = 32'd136314880;
      5220: inst = 32'd268468224;
      5221: inst = 32'd201344249;
      5222: inst = 32'd203489279;
      5223: inst = 32'd136314880;
      5224: inst = 32'd268468224;
      5225: inst = 32'd201344250;
      5226: inst = 32'd203489279;
      5227: inst = 32'd136314880;
      5228: inst = 32'd268468224;
      5229: inst = 32'd201344251;
      5230: inst = 32'd203489279;
      5231: inst = 32'd136314880;
      5232: inst = 32'd268468224;
      5233: inst = 32'd201344252;
      5234: inst = 32'd203489279;
      5235: inst = 32'd136314880;
      5236: inst = 32'd268468224;
      5237: inst = 32'd201344253;
      5238: inst = 32'd203489279;
      5239: inst = 32'd136314880;
      5240: inst = 32'd268468224;
      5241: inst = 32'd201344254;
      5242: inst = 32'd203489279;
      5243: inst = 32'd136314880;
      5244: inst = 32'd268468224;
      5245: inst = 32'd201344255;
      5246: inst = 32'd203489279;
      5247: inst = 32'd136314880;
      5248: inst = 32'd268468224;
      5249: inst = 32'd201344256;
      5250: inst = 32'd203489279;
      5251: inst = 32'd136314880;
      5252: inst = 32'd268468224;
      5253: inst = 32'd201344257;
      5254: inst = 32'd203489279;
      5255: inst = 32'd136314880;
      5256: inst = 32'd268468224;
      5257: inst = 32'd201344258;
      5258: inst = 32'd203489279;
      5259: inst = 32'd136314880;
      5260: inst = 32'd268468224;
      5261: inst = 32'd201344259;
      5262: inst = 32'd203489278;
      5263: inst = 32'd136314880;
      5264: inst = 32'd268468224;
      5265: inst = 32'd201344260;
      5266: inst = 32'd203482808;
      5267: inst = 32'd136314880;
      5268: inst = 32'd268468224;
      5269: inst = 32'd201344261;
      5270: inst = 32'd203484855;
      5271: inst = 32'd136314880;
      5272: inst = 32'd268468224;
      5273: inst = 32'd201344262;
      5274: inst = 32'd203484854;
      5275: inst = 32'd136314880;
      5276: inst = 32'd268468224;
      5277: inst = 32'd201344263;
      5278: inst = 32'd203484854;
      5279: inst = 32'd136314880;
      5280: inst = 32'd268468224;
      5281: inst = 32'd201344264;
      5282: inst = 32'd203484854;
      5283: inst = 32'd136314880;
      5284: inst = 32'd268468224;
      5285: inst = 32'd201344265;
      5286: inst = 32'd203484854;
      5287: inst = 32'd136314880;
      5288: inst = 32'd268468224;
      5289: inst = 32'd201344266;
      5290: inst = 32'd203484854;
      5291: inst = 32'd136314880;
      5292: inst = 32'd268468224;
      5293: inst = 32'd201344267;
      5294: inst = 32'd203484854;
      5295: inst = 32'd136314880;
      5296: inst = 32'd268468224;
      5297: inst = 32'd201344268;
      5298: inst = 32'd203484854;
      5299: inst = 32'd136314880;
      5300: inst = 32'd268468224;
      5301: inst = 32'd201344269;
      5302: inst = 32'd203484854;
      5303: inst = 32'd136314880;
      5304: inst = 32'd268468224;
      5305: inst = 32'd201344270;
      5306: inst = 32'd203484854;
      5307: inst = 32'd136314880;
      5308: inst = 32'd268468224;
      5309: inst = 32'd201344271;
      5310: inst = 32'd203484854;
      5311: inst = 32'd136314880;
      5312: inst = 32'd268468224;
      5313: inst = 32'd201344272;
      5314: inst = 32'd203486934;
      5315: inst = 32'd136314880;
      5316: inst = 32'd268468224;
      5317: inst = 32'd201344273;
      5318: inst = 32'd203484886;
      5319: inst = 32'd136314880;
      5320: inst = 32'd268468224;
      5321: inst = 32'd201344274;
      5322: inst = 32'd203484853;
      5323: inst = 32'd136314880;
      5324: inst = 32'd268468224;
      5325: inst = 32'd201344275;
      5326: inst = 32'd203484853;
      5327: inst = 32'd136314880;
      5328: inst = 32'd268468224;
      5329: inst = 32'd201344276;
      5330: inst = 32'd203484853;
      5331: inst = 32'd136314880;
      5332: inst = 32'd268468224;
      5333: inst = 32'd201344277;
      5334: inst = 32'd203484854;
      5335: inst = 32'd136314880;
      5336: inst = 32'd268468224;
      5337: inst = 32'd201344278;
      5338: inst = 32'd203484886;
      5339: inst = 32'd136314880;
      5340: inst = 32'd268468224;
      5341: inst = 32'd201344279;
      5342: inst = 32'd203486934;
      5343: inst = 32'd136314880;
      5344: inst = 32'd268468224;
      5345: inst = 32'd201344280;
      5346: inst = 32'd203484854;
      5347: inst = 32'd136314880;
      5348: inst = 32'd268468224;
      5349: inst = 32'd201344281;
      5350: inst = 32'd203484854;
      5351: inst = 32'd136314880;
      5352: inst = 32'd268468224;
      5353: inst = 32'd201344282;
      5354: inst = 32'd203484854;
      5355: inst = 32'd136314880;
      5356: inst = 32'd268468224;
      5357: inst = 32'd201344283;
      5358: inst = 32'd203484854;
      5359: inst = 32'd136314880;
      5360: inst = 32'd268468224;
      5361: inst = 32'd201344284;
      5362: inst = 32'd203484854;
      5363: inst = 32'd136314880;
      5364: inst = 32'd268468224;
      5365: inst = 32'd201344285;
      5366: inst = 32'd203484854;
      5367: inst = 32'd136314880;
      5368: inst = 32'd268468224;
      5369: inst = 32'd201344286;
      5370: inst = 32'd203484854;
      5371: inst = 32'd136314880;
      5372: inst = 32'd268468224;
      5373: inst = 32'd201344287;
      5374: inst = 32'd203484854;
      5375: inst = 32'd136314880;
      5376: inst = 32'd268468224;
      5377: inst = 32'd201344288;
      5378: inst = 32'd203486934;
      5379: inst = 32'd136314880;
      5380: inst = 32'd268468224;
      5381: inst = 32'd201344289;
      5382: inst = 32'd203486934;
      5383: inst = 32'd136314880;
      5384: inst = 32'd268468224;
      5385: inst = 32'd201344290;
      5386: inst = 32'd203486902;
      5387: inst = 32'd136314880;
      5388: inst = 32'd268468224;
      5389: inst = 32'd201344291;
      5390: inst = 32'd203484822;
      5391: inst = 32'd136314880;
      5392: inst = 32'd268468224;
      5393: inst = 32'd201344292;
      5394: inst = 32'd203482742;
      5395: inst = 32'd136314880;
      5396: inst = 32'd268468224;
      5397: inst = 32'd201344293;
      5398: inst = 32'd203482774;
      5399: inst = 32'd136314880;
      5400: inst = 32'd268468224;
      5401: inst = 32'd201344294;
      5402: inst = 32'd203482806;
      5403: inst = 32'd136314880;
      5404: inst = 32'd268468224;
      5405: inst = 32'd201344295;
      5406: inst = 32'd203484887;
      5407: inst = 32'd136314880;
      5408: inst = 32'd268468224;
      5409: inst = 32'd201344296;
      5410: inst = 32'd203482773;
      5411: inst = 32'd136314880;
      5412: inst = 32'd268468224;
      5413: inst = 32'd201344297;
      5414: inst = 32'd203486998;
      5415: inst = 32'd136314880;
      5416: inst = 32'd268468224;
      5417: inst = 32'd201344298;
      5418: inst = 32'd203482804;
      5419: inst = 32'd136314880;
      5420: inst = 32'd268468224;
      5421: inst = 32'd201344299;
      5422: inst = 32'd203484917;
      5423: inst = 32'd136314880;
      5424: inst = 32'd268468224;
      5425: inst = 32'd201344300;
      5426: inst = 32'd203484918;
      5427: inst = 32'd136314880;
      5428: inst = 32'd268468224;
      5429: inst = 32'd201344301;
      5430: inst = 32'd203480757;
      5431: inst = 32'd136314880;
      5432: inst = 32'd268468224;
      5433: inst = 32'd201344302;
      5434: inst = 32'd203484951;
      5435: inst = 32'd136314880;
      5436: inst = 32'd268468224;
      5437: inst = 32'd201344303;
      5438: inst = 32'd203480758;
      5439: inst = 32'd136314880;
      5440: inst = 32'd268468224;
      5441: inst = 32'd201344304;
      5442: inst = 32'd203486903;
      5443: inst = 32'd136314880;
      5444: inst = 32'd268468224;
      5445: inst = 32'd201344305;
      5446: inst = 32'd203484822;
      5447: inst = 32'd136314880;
      5448: inst = 32'd268468224;
      5449: inst = 32'd201344306;
      5450: inst = 32'd203482742;
      5451: inst = 32'd136314880;
      5452: inst = 32'd268468224;
      5453: inst = 32'd201344307;
      5454: inst = 32'd203482742;
      5455: inst = 32'd136314880;
      5456: inst = 32'd268468224;
      5457: inst = 32'd201344308;
      5458: inst = 32'd203484854;
      5459: inst = 32'd136314880;
      5460: inst = 32'd268468224;
      5461: inst = 32'd201344309;
      5462: inst = 32'd203484886;
      5463: inst = 32'd136314880;
      5464: inst = 32'd268468224;
      5465: inst = 32'd201344310;
      5466: inst = 32'd203486934;
      5467: inst = 32'd136314880;
      5468: inst = 32'd268468224;
      5469: inst = 32'd201344311;
      5470: inst = 32'd203486934;
      5471: inst = 32'd136314880;
      5472: inst = 32'd268468224;
      5473: inst = 32'd201344312;
      5474: inst = 32'd203484854;
      5475: inst = 32'd136314880;
      5476: inst = 32'd268468224;
      5477: inst = 32'd201344313;
      5478: inst = 32'd203484854;
      5479: inst = 32'd136314880;
      5480: inst = 32'd268468224;
      5481: inst = 32'd201344314;
      5482: inst = 32'd203484887;
      5483: inst = 32'd136314880;
      5484: inst = 32'd268468224;
      5485: inst = 32'd201344315;
      5486: inst = 32'd203482808;
      5487: inst = 32'd136314880;
      5488: inst = 32'd268468224;
      5489: inst = 32'd201344316;
      5490: inst = 32'd203489277;
      5491: inst = 32'd136314880;
      5492: inst = 32'd268468224;
      5493: inst = 32'd201344317;
      5494: inst = 32'd203489278;
      5495: inst = 32'd136314880;
      5496: inst = 32'd268468224;
      5497: inst = 32'd201344318;
      5498: inst = 32'd203489279;
      5499: inst = 32'd136314880;
      5500: inst = 32'd268468224;
      5501: inst = 32'd201344319;
      5502: inst = 32'd203489279;
      5503: inst = 32'd136314880;
      5504: inst = 32'd268468224;
      5505: inst = 32'd201344320;
      5506: inst = 32'd203489279;
      5507: inst = 32'd136314880;
      5508: inst = 32'd268468224;
      5509: inst = 32'd201344321;
      5510: inst = 32'd203489279;
      5511: inst = 32'd136314880;
      5512: inst = 32'd268468224;
      5513: inst = 32'd201344322;
      5514: inst = 32'd203489279;
      5515: inst = 32'd136314880;
      5516: inst = 32'd268468224;
      5517: inst = 32'd201344323;
      5518: inst = 32'd203489279;
      5519: inst = 32'd136314880;
      5520: inst = 32'd268468224;
      5521: inst = 32'd201344324;
      5522: inst = 32'd203489279;
      5523: inst = 32'd136314880;
      5524: inst = 32'd268468224;
      5525: inst = 32'd201344325;
      5526: inst = 32'd203489279;
      5527: inst = 32'd136314880;
      5528: inst = 32'd268468224;
      5529: inst = 32'd201344326;
      5530: inst = 32'd203489279;
      5531: inst = 32'd136314880;
      5532: inst = 32'd268468224;
      5533: inst = 32'd201344327;
      5534: inst = 32'd203489279;
      5535: inst = 32'd136314880;
      5536: inst = 32'd268468224;
      5537: inst = 32'd201344328;
      5538: inst = 32'd203489279;
      5539: inst = 32'd136314880;
      5540: inst = 32'd268468224;
      5541: inst = 32'd201344329;
      5542: inst = 32'd203489279;
      5543: inst = 32'd136314880;
      5544: inst = 32'd268468224;
      5545: inst = 32'd201344330;
      5546: inst = 32'd203489279;
      5547: inst = 32'd136314880;
      5548: inst = 32'd268468224;
      5549: inst = 32'd201344331;
      5550: inst = 32'd203489279;
      5551: inst = 32'd136314880;
      5552: inst = 32'd268468224;
      5553: inst = 32'd201344332;
      5554: inst = 32'd203489279;
      5555: inst = 32'd136314880;
      5556: inst = 32'd268468224;
      5557: inst = 32'd201344333;
      5558: inst = 32'd203489279;
      5559: inst = 32'd136314880;
      5560: inst = 32'd268468224;
      5561: inst = 32'd201344334;
      5562: inst = 32'd203489279;
      5563: inst = 32'd136314880;
      5564: inst = 32'd268468224;
      5565: inst = 32'd201344335;
      5566: inst = 32'd203489279;
      5567: inst = 32'd136314880;
      5568: inst = 32'd268468224;
      5569: inst = 32'd201344336;
      5570: inst = 32'd203489279;
      5571: inst = 32'd136314880;
      5572: inst = 32'd268468224;
      5573: inst = 32'd201344337;
      5574: inst = 32'd203489279;
      5575: inst = 32'd136314880;
      5576: inst = 32'd268468224;
      5577: inst = 32'd201344338;
      5578: inst = 32'd203489279;
      5579: inst = 32'd136314880;
      5580: inst = 32'd268468224;
      5581: inst = 32'd201344339;
      5582: inst = 32'd203489279;
      5583: inst = 32'd136314880;
      5584: inst = 32'd268468224;
      5585: inst = 32'd201344340;
      5586: inst = 32'd203489279;
      5587: inst = 32'd136314880;
      5588: inst = 32'd268468224;
      5589: inst = 32'd201344341;
      5590: inst = 32'd203489279;
      5591: inst = 32'd136314880;
      5592: inst = 32'd268468224;
      5593: inst = 32'd201344342;
      5594: inst = 32'd203489279;
      5595: inst = 32'd136314880;
      5596: inst = 32'd268468224;
      5597: inst = 32'd201344343;
      5598: inst = 32'd203489279;
      5599: inst = 32'd136314880;
      5600: inst = 32'd268468224;
      5601: inst = 32'd201344344;
      5602: inst = 32'd203489279;
      5603: inst = 32'd136314880;
      5604: inst = 32'd268468224;
      5605: inst = 32'd201344345;
      5606: inst = 32'd203489279;
      5607: inst = 32'd136314880;
      5608: inst = 32'd268468224;
      5609: inst = 32'd201344346;
      5610: inst = 32'd203489279;
      5611: inst = 32'd136314880;
      5612: inst = 32'd268468224;
      5613: inst = 32'd201344347;
      5614: inst = 32'd203489279;
      5615: inst = 32'd136314880;
      5616: inst = 32'd268468224;
      5617: inst = 32'd201344348;
      5618: inst = 32'd203489279;
      5619: inst = 32'd136314880;
      5620: inst = 32'd268468224;
      5621: inst = 32'd201344349;
      5622: inst = 32'd203489279;
      5623: inst = 32'd136314880;
      5624: inst = 32'd268468224;
      5625: inst = 32'd201344350;
      5626: inst = 32'd203489279;
      5627: inst = 32'd136314880;
      5628: inst = 32'd268468224;
      5629: inst = 32'd201344351;
      5630: inst = 32'd203489279;
      5631: inst = 32'd136314880;
      5632: inst = 32'd268468224;
      5633: inst = 32'd201344352;
      5634: inst = 32'd203489279;
      5635: inst = 32'd136314880;
      5636: inst = 32'd268468224;
      5637: inst = 32'd201344353;
      5638: inst = 32'd203489279;
      5639: inst = 32'd136314880;
      5640: inst = 32'd268468224;
      5641: inst = 32'd201344354;
      5642: inst = 32'd203489278;
      5643: inst = 32'd136314880;
      5644: inst = 32'd268468224;
      5645: inst = 32'd201344355;
      5646: inst = 32'd203489277;
      5647: inst = 32'd136314880;
      5648: inst = 32'd268468224;
      5649: inst = 32'd201344356;
      5650: inst = 32'd203482808;
      5651: inst = 32'd136314880;
      5652: inst = 32'd268468224;
      5653: inst = 32'd201344357;
      5654: inst = 32'd203484887;
      5655: inst = 32'd136314880;
      5656: inst = 32'd268468224;
      5657: inst = 32'd201344358;
      5658: inst = 32'd203484854;
      5659: inst = 32'd136314880;
      5660: inst = 32'd268468224;
      5661: inst = 32'd201344359;
      5662: inst = 32'd203484854;
      5663: inst = 32'd136314880;
      5664: inst = 32'd268468224;
      5665: inst = 32'd201344360;
      5666: inst = 32'd203484854;
      5667: inst = 32'd136314880;
      5668: inst = 32'd268468224;
      5669: inst = 32'd201344361;
      5670: inst = 32'd203484854;
      5671: inst = 32'd136314880;
      5672: inst = 32'd268468224;
      5673: inst = 32'd201344362;
      5674: inst = 32'd203484854;
      5675: inst = 32'd136314880;
      5676: inst = 32'd268468224;
      5677: inst = 32'd201344363;
      5678: inst = 32'd203484854;
      5679: inst = 32'd136314880;
      5680: inst = 32'd268468224;
      5681: inst = 32'd201344364;
      5682: inst = 32'd203484854;
      5683: inst = 32'd136314880;
      5684: inst = 32'd268468224;
      5685: inst = 32'd201344365;
      5686: inst = 32'd203484854;
      5687: inst = 32'd136314880;
      5688: inst = 32'd268468224;
      5689: inst = 32'd201344366;
      5690: inst = 32'd203484855;
      5691: inst = 32'd136314880;
      5692: inst = 32'd268468224;
      5693: inst = 32'd201344367;
      5694: inst = 32'd203484855;
      5695: inst = 32'd136314880;
      5696: inst = 32'd268468224;
      5697: inst = 32'd201344368;
      5698: inst = 32'd203484821;
      5699: inst = 32'd136314880;
      5700: inst = 32'd268468224;
      5701: inst = 32'd201344369;
      5702: inst = 32'd203484853;
      5703: inst = 32'd136314880;
      5704: inst = 32'd268468224;
      5705: inst = 32'd201344370;
      5706: inst = 32'd203484854;
      5707: inst = 32'd136314880;
      5708: inst = 32'd268468224;
      5709: inst = 32'd201344371;
      5710: inst = 32'd203484886;
      5711: inst = 32'd136314880;
      5712: inst = 32'd268468224;
      5713: inst = 32'd201344372;
      5714: inst = 32'd203484886;
      5715: inst = 32'd136314880;
      5716: inst = 32'd268468224;
      5717: inst = 32'd201344373;
      5718: inst = 32'd203484854;
      5719: inst = 32'd136314880;
      5720: inst = 32'd268468224;
      5721: inst = 32'd201344374;
      5722: inst = 32'd203484853;
      5723: inst = 32'd136314880;
      5724: inst = 32'd268468224;
      5725: inst = 32'd201344375;
      5726: inst = 32'd203484821;
      5727: inst = 32'd136314880;
      5728: inst = 32'd268468224;
      5729: inst = 32'd201344376;
      5730: inst = 32'd203484854;
      5731: inst = 32'd136314880;
      5732: inst = 32'd268468224;
      5733: inst = 32'd201344377;
      5734: inst = 32'd203484854;
      5735: inst = 32'd136314880;
      5736: inst = 32'd268468224;
      5737: inst = 32'd201344378;
      5738: inst = 32'd203484854;
      5739: inst = 32'd136314880;
      5740: inst = 32'd268468224;
      5741: inst = 32'd201344379;
      5742: inst = 32'd203484854;
      5743: inst = 32'd136314880;
      5744: inst = 32'd268468224;
      5745: inst = 32'd201344380;
      5746: inst = 32'd203484854;
      5747: inst = 32'd136314880;
      5748: inst = 32'd268468224;
      5749: inst = 32'd201344381;
      5750: inst = 32'd203484854;
      5751: inst = 32'd136314880;
      5752: inst = 32'd268468224;
      5753: inst = 32'd201344382;
      5754: inst = 32'd203484854;
      5755: inst = 32'd136314880;
      5756: inst = 32'd268468224;
      5757: inst = 32'd201344383;
      5758: inst = 32'd203484854;
      5759: inst = 32'd136314880;
      5760: inst = 32'd268468224;
      5761: inst = 32'd201344384;
      5762: inst = 32'd203484821;
      5763: inst = 32'd136314880;
      5764: inst = 32'd268468224;
      5765: inst = 32'd201344385;
      5766: inst = 32'd203484854;
      5767: inst = 32'd136314880;
      5768: inst = 32'd268468224;
      5769: inst = 32'd201344386;
      5770: inst = 32'd203486934;
      5771: inst = 32'd136314880;
      5772: inst = 32'd268468224;
      5773: inst = 32'd201344387;
      5774: inst = 32'd203484855;
      5775: inst = 32'd136314880;
      5776: inst = 32'd268468224;
      5777: inst = 32'd201344388;
      5778: inst = 32'd203484855;
      5779: inst = 32'd136314880;
      5780: inst = 32'd268468224;
      5781: inst = 32'd201344389;
      5782: inst = 32'd203484888;
      5783: inst = 32'd136314880;
      5784: inst = 32'd268468224;
      5785: inst = 32'd201344390;
      5786: inst = 32'd203484887;
      5787: inst = 32'd136314880;
      5788: inst = 32'd268468224;
      5789: inst = 32'd201344391;
      5790: inst = 32'd203484854;
      5791: inst = 32'd136314880;
      5792: inst = 32'd268468224;
      5793: inst = 32'd201344392;
      5794: inst = 32'd203484886;
      5795: inst = 32'd136314880;
      5796: inst = 32'd268468224;
      5797: inst = 32'd201344393;
      5798: inst = 32'd203482837;
      5799: inst = 32'd136314880;
      5800: inst = 32'd268468224;
      5801: inst = 32'd201344394;
      5802: inst = 32'd203484918;
      5803: inst = 32'd136314880;
      5804: inst = 32'd268468224;
      5805: inst = 32'd201344395;
      5806: inst = 32'd203482837;
      5807: inst = 32'd136314880;
      5808: inst = 32'd268468224;
      5809: inst = 32'd201344396;
      5810: inst = 32'd203482837;
      5811: inst = 32'd136314880;
      5812: inst = 32'd268468224;
      5813: inst = 32'd201344397;
      5814: inst = 32'd203482871;
      5815: inst = 32'd136314880;
      5816: inst = 32'd268468224;
      5817: inst = 32'd201344398;
      5818: inst = 32'd203482839;
      5819: inst = 32'd136314880;
      5820: inst = 32'd268468224;
      5821: inst = 32'd201344399;
      5822: inst = 32'd203482839;
      5823: inst = 32'd136314880;
      5824: inst = 32'd268468224;
      5825: inst = 32'd201344400;
      5826: inst = 32'd203484855;
      5827: inst = 32'd136314880;
      5828: inst = 32'd268468224;
      5829: inst = 32'd201344401;
      5830: inst = 32'd203486903;
      5831: inst = 32'd136314880;
      5832: inst = 32'd268468224;
      5833: inst = 32'd201344402;
      5834: inst = 32'd203486935;
      5835: inst = 32'd136314880;
      5836: inst = 32'd268468224;
      5837: inst = 32'd201344403;
      5838: inst = 32'd203486903;
      5839: inst = 32'd136314880;
      5840: inst = 32'd268468224;
      5841: inst = 32'd201344404;
      5842: inst = 32'd203484854;
      5843: inst = 32'd136314880;
      5844: inst = 32'd268468224;
      5845: inst = 32'd201344405;
      5846: inst = 32'd203484886;
      5847: inst = 32'd136314880;
      5848: inst = 32'd268468224;
      5849: inst = 32'd201344406;
      5850: inst = 32'd203484854;
      5851: inst = 32'd136314880;
      5852: inst = 32'd268468224;
      5853: inst = 32'd201344407;
      5854: inst = 32'd203484821;
      5855: inst = 32'd136314880;
      5856: inst = 32'd268468224;
      5857: inst = 32'd201344408;
      5858: inst = 32'd203484854;
      5859: inst = 32'd136314880;
      5860: inst = 32'd268468224;
      5861: inst = 32'd201344409;
      5862: inst = 32'd203484854;
      5863: inst = 32'd136314880;
      5864: inst = 32'd268468224;
      5865: inst = 32'd201344410;
      5866: inst = 32'd203484887;
      5867: inst = 32'd136314880;
      5868: inst = 32'd268468224;
      5869: inst = 32'd201344411;
      5870: inst = 32'd203482808;
      5871: inst = 32'd136314880;
      5872: inst = 32'd268468224;
      5873: inst = 32'd201344412;
      5874: inst = 32'd203489277;
      5875: inst = 32'd136314880;
      5876: inst = 32'd268468224;
      5877: inst = 32'd201344413;
      5878: inst = 32'd203489278;
      5879: inst = 32'd136314880;
      5880: inst = 32'd268468224;
      5881: inst = 32'd201344414;
      5882: inst = 32'd203489279;
      5883: inst = 32'd136314880;
      5884: inst = 32'd268468224;
      5885: inst = 32'd201344415;
      5886: inst = 32'd203489279;
      5887: inst = 32'd136314880;
      5888: inst = 32'd268468224;
      5889: inst = 32'd201344416;
      5890: inst = 32'd203489279;
      5891: inst = 32'd136314880;
      5892: inst = 32'd268468224;
      5893: inst = 32'd201344417;
      5894: inst = 32'd203489279;
      5895: inst = 32'd136314880;
      5896: inst = 32'd268468224;
      5897: inst = 32'd201344418;
      5898: inst = 32'd203489279;
      5899: inst = 32'd136314880;
      5900: inst = 32'd268468224;
      5901: inst = 32'd201344419;
      5902: inst = 32'd203489279;
      5903: inst = 32'd136314880;
      5904: inst = 32'd268468224;
      5905: inst = 32'd201344420;
      5906: inst = 32'd203489279;
      5907: inst = 32'd136314880;
      5908: inst = 32'd268468224;
      5909: inst = 32'd201344421;
      5910: inst = 32'd203489279;
      5911: inst = 32'd136314880;
      5912: inst = 32'd268468224;
      5913: inst = 32'd201344422;
      5914: inst = 32'd203489279;
      5915: inst = 32'd136314880;
      5916: inst = 32'd268468224;
      5917: inst = 32'd201344423;
      5918: inst = 32'd203489279;
      5919: inst = 32'd136314880;
      5920: inst = 32'd268468224;
      5921: inst = 32'd201344424;
      5922: inst = 32'd203489279;
      5923: inst = 32'd136314880;
      5924: inst = 32'd268468224;
      5925: inst = 32'd201344425;
      5926: inst = 32'd203489279;
      5927: inst = 32'd136314880;
      5928: inst = 32'd268468224;
      5929: inst = 32'd201344426;
      5930: inst = 32'd203489279;
      5931: inst = 32'd136314880;
      5932: inst = 32'd268468224;
      5933: inst = 32'd201344427;
      5934: inst = 32'd203489279;
      5935: inst = 32'd136314880;
      5936: inst = 32'd268468224;
      5937: inst = 32'd201344428;
      5938: inst = 32'd203489279;
      5939: inst = 32'd136314880;
      5940: inst = 32'd268468224;
      5941: inst = 32'd201344429;
      5942: inst = 32'd203489279;
      5943: inst = 32'd136314880;
      5944: inst = 32'd268468224;
      5945: inst = 32'd201344430;
      5946: inst = 32'd203489279;
      5947: inst = 32'd136314880;
      5948: inst = 32'd268468224;
      5949: inst = 32'd201344431;
      5950: inst = 32'd203489279;
      5951: inst = 32'd136314880;
      5952: inst = 32'd268468224;
      5953: inst = 32'd201344432;
      5954: inst = 32'd203489279;
      5955: inst = 32'd136314880;
      5956: inst = 32'd268468224;
      5957: inst = 32'd201344433;
      5958: inst = 32'd203489279;
      5959: inst = 32'd136314880;
      5960: inst = 32'd268468224;
      5961: inst = 32'd201344434;
      5962: inst = 32'd203489279;
      5963: inst = 32'd136314880;
      5964: inst = 32'd268468224;
      5965: inst = 32'd201344435;
      5966: inst = 32'd203489279;
      5967: inst = 32'd136314880;
      5968: inst = 32'd268468224;
      5969: inst = 32'd201344436;
      5970: inst = 32'd203489279;
      5971: inst = 32'd136314880;
      5972: inst = 32'd268468224;
      5973: inst = 32'd201344437;
      5974: inst = 32'd203489279;
      5975: inst = 32'd136314880;
      5976: inst = 32'd268468224;
      5977: inst = 32'd201344438;
      5978: inst = 32'd203489279;
      5979: inst = 32'd136314880;
      5980: inst = 32'd268468224;
      5981: inst = 32'd201344439;
      5982: inst = 32'd203489279;
      5983: inst = 32'd136314880;
      5984: inst = 32'd268468224;
      5985: inst = 32'd201344440;
      5986: inst = 32'd203489279;
      5987: inst = 32'd136314880;
      5988: inst = 32'd268468224;
      5989: inst = 32'd201344441;
      5990: inst = 32'd203489279;
      5991: inst = 32'd136314880;
      5992: inst = 32'd268468224;
      5993: inst = 32'd201344442;
      5994: inst = 32'd203489279;
      5995: inst = 32'd136314880;
      5996: inst = 32'd268468224;
      5997: inst = 32'd201344443;
      5998: inst = 32'd203489279;
      5999: inst = 32'd136314880;
      6000: inst = 32'd268468224;
      6001: inst = 32'd201344444;
      6002: inst = 32'd203489279;
      6003: inst = 32'd136314880;
      6004: inst = 32'd268468224;
      6005: inst = 32'd201344445;
      6006: inst = 32'd203489279;
      6007: inst = 32'd136314880;
      6008: inst = 32'd268468224;
      6009: inst = 32'd201344446;
      6010: inst = 32'd203489279;
      6011: inst = 32'd136314880;
      6012: inst = 32'd268468224;
      6013: inst = 32'd201344447;
      6014: inst = 32'd203489279;
      6015: inst = 32'd136314880;
      6016: inst = 32'd268468224;
      6017: inst = 32'd201344448;
      6018: inst = 32'd203489279;
      6019: inst = 32'd136314880;
      6020: inst = 32'd268468224;
      6021: inst = 32'd201344449;
      6022: inst = 32'd203489279;
      6023: inst = 32'd136314880;
      6024: inst = 32'd268468224;
      6025: inst = 32'd201344450;
      6026: inst = 32'd203489278;
      6027: inst = 32'd136314880;
      6028: inst = 32'd268468224;
      6029: inst = 32'd201344451;
      6030: inst = 32'd203489277;
      6031: inst = 32'd136314880;
      6032: inst = 32'd268468224;
      6033: inst = 32'd201344452;
      6034: inst = 32'd203482808;
      6035: inst = 32'd136314880;
      6036: inst = 32'd268468224;
      6037: inst = 32'd201344453;
      6038: inst = 32'd203484855;
      6039: inst = 32'd136314880;
      6040: inst = 32'd268468224;
      6041: inst = 32'd201344454;
      6042: inst = 32'd203484854;
      6043: inst = 32'd136314880;
      6044: inst = 32'd268468224;
      6045: inst = 32'd201344455;
      6046: inst = 32'd203484854;
      6047: inst = 32'd136314880;
      6048: inst = 32'd268468224;
      6049: inst = 32'd201344456;
      6050: inst = 32'd203484853;
      6051: inst = 32'd136314880;
      6052: inst = 32'd268468224;
      6053: inst = 32'd201344457;
      6054: inst = 32'd203484854;
      6055: inst = 32'd136314880;
      6056: inst = 32'd268468224;
      6057: inst = 32'd201344458;
      6058: inst = 32'd203484854;
      6059: inst = 32'd136314880;
      6060: inst = 32'd268468224;
      6061: inst = 32'd201344459;
      6062: inst = 32'd203484854;
      6063: inst = 32'd136314880;
      6064: inst = 32'd268468224;
      6065: inst = 32'd201344460;
      6066: inst = 32'd203484854;
      6067: inst = 32'd136314880;
      6068: inst = 32'd268468224;
      6069: inst = 32'd201344461;
      6070: inst = 32'd203484854;
      6071: inst = 32'd136314880;
      6072: inst = 32'd268468224;
      6073: inst = 32'd201344462;
      6074: inst = 32'd203484855;
      6075: inst = 32'd136314880;
      6076: inst = 32'd268468224;
      6077: inst = 32'd201344463;
      6078: inst = 32'd203484855;
      6079: inst = 32'd136314880;
      6080: inst = 32'd268468224;
      6081: inst = 32'd201344464;
      6082: inst = 32'd203484886;
      6083: inst = 32'd136314880;
      6084: inst = 32'd268468224;
      6085: inst = 32'd201344465;
      6086: inst = 32'd203484886;
      6087: inst = 32'd136314880;
      6088: inst = 32'd268468224;
      6089: inst = 32'd201344466;
      6090: inst = 32'd203484854;
      6091: inst = 32'd136314880;
      6092: inst = 32'd268468224;
      6093: inst = 32'd201344467;
      6094: inst = 32'd203484853;
      6095: inst = 32'd136314880;
      6096: inst = 32'd268468224;
      6097: inst = 32'd201344468;
      6098: inst = 32'd203484853;
      6099: inst = 32'd136314880;
      6100: inst = 32'd268468224;
      6101: inst = 32'd201344469;
      6102: inst = 32'd203484854;
      6103: inst = 32'd136314880;
      6104: inst = 32'd268468224;
      6105: inst = 32'd201344470;
      6106: inst = 32'd203484886;
      6107: inst = 32'd136314880;
      6108: inst = 32'd268468224;
      6109: inst = 32'd201344471;
      6110: inst = 32'd203484886;
      6111: inst = 32'd136314880;
      6112: inst = 32'd268468224;
      6113: inst = 32'd201344472;
      6114: inst = 32'd203484854;
      6115: inst = 32'd136314880;
      6116: inst = 32'd268468224;
      6117: inst = 32'd201344473;
      6118: inst = 32'd203484854;
      6119: inst = 32'd136314880;
      6120: inst = 32'd268468224;
      6121: inst = 32'd201344474;
      6122: inst = 32'd203484854;
      6123: inst = 32'd136314880;
      6124: inst = 32'd268468224;
      6125: inst = 32'd201344475;
      6126: inst = 32'd203484854;
      6127: inst = 32'd136314880;
      6128: inst = 32'd268468224;
      6129: inst = 32'd201344476;
      6130: inst = 32'd203484854;
      6131: inst = 32'd136314880;
      6132: inst = 32'd268468224;
      6133: inst = 32'd201344477;
      6134: inst = 32'd203484854;
      6135: inst = 32'd136314880;
      6136: inst = 32'd268468224;
      6137: inst = 32'd201344478;
      6138: inst = 32'd203484854;
      6139: inst = 32'd136314880;
      6140: inst = 32'd268468224;
      6141: inst = 32'd201344479;
      6142: inst = 32'd203484854;
      6143: inst = 32'd136314880;
      6144: inst = 32'd268468224;
      6145: inst = 32'd201344480;
      6146: inst = 32'd203484854;
      6147: inst = 32'd136314880;
      6148: inst = 32'd268468224;
      6149: inst = 32'd201344481;
      6150: inst = 32'd203484854;
      6151: inst = 32'd136314880;
      6152: inst = 32'd268468224;
      6153: inst = 32'd201344482;
      6154: inst = 32'd203484854;
      6155: inst = 32'd136314880;
      6156: inst = 32'd268468224;
      6157: inst = 32'd201344483;
      6158: inst = 32'd203484854;
      6159: inst = 32'd136314880;
      6160: inst = 32'd268468224;
      6161: inst = 32'd201344484;
      6162: inst = 32'd203484854;
      6163: inst = 32'd136314880;
      6164: inst = 32'd268468224;
      6165: inst = 32'd201344485;
      6166: inst = 32'd203484854;
      6167: inst = 32'd136314880;
      6168: inst = 32'd268468224;
      6169: inst = 32'd201344486;
      6170: inst = 32'd203484854;
      6171: inst = 32'd136314880;
      6172: inst = 32'd268468224;
      6173: inst = 32'd201344487;
      6174: inst = 32'd203484854;
      6175: inst = 32'd136314880;
      6176: inst = 32'd268468224;
      6177: inst = 32'd201344488;
      6178: inst = 32'd203484854;
      6179: inst = 32'd136314880;
      6180: inst = 32'd268468224;
      6181: inst = 32'd201344489;
      6182: inst = 32'd203484854;
      6183: inst = 32'd136314880;
      6184: inst = 32'd268468224;
      6185: inst = 32'd201344490;
      6186: inst = 32'd203484886;
      6187: inst = 32'd136314880;
      6188: inst = 32'd268468224;
      6189: inst = 32'd201344491;
      6190: inst = 32'd203484886;
      6191: inst = 32'd136314880;
      6192: inst = 32'd268468224;
      6193: inst = 32'd201344492;
      6194: inst = 32'd203484886;
      6195: inst = 32'd136314880;
      6196: inst = 32'd268468224;
      6197: inst = 32'd201344493;
      6198: inst = 32'd203482838;
      6199: inst = 32'd136314880;
      6200: inst = 32'd268468224;
      6201: inst = 32'd201344494;
      6202: inst = 32'd203482838;
      6203: inst = 32'd136314880;
      6204: inst = 32'd268468224;
      6205: inst = 32'd201344495;
      6206: inst = 32'd203482839;
      6207: inst = 32'd136314880;
      6208: inst = 32'd268468224;
      6209: inst = 32'd201344496;
      6210: inst = 32'd203484854;
      6211: inst = 32'd136314880;
      6212: inst = 32'd268468224;
      6213: inst = 32'd201344497;
      6214: inst = 32'd203484854;
      6215: inst = 32'd136314880;
      6216: inst = 32'd268468224;
      6217: inst = 32'd201344498;
      6218: inst = 32'd203484854;
      6219: inst = 32'd136314880;
      6220: inst = 32'd268468224;
      6221: inst = 32'd201344499;
      6222: inst = 32'd203484854;
      6223: inst = 32'd136314880;
      6224: inst = 32'd268468224;
      6225: inst = 32'd201344500;
      6226: inst = 32'd203484854;
      6227: inst = 32'd136314880;
      6228: inst = 32'd268468224;
      6229: inst = 32'd201344501;
      6230: inst = 32'd203484854;
      6231: inst = 32'd136314880;
      6232: inst = 32'd268468224;
      6233: inst = 32'd201344502;
      6234: inst = 32'd203484854;
      6235: inst = 32'd136314880;
      6236: inst = 32'd268468224;
      6237: inst = 32'd201344503;
      6238: inst = 32'd203484854;
      6239: inst = 32'd136314880;
      6240: inst = 32'd268468224;
      6241: inst = 32'd201344504;
      6242: inst = 32'd203484854;
      6243: inst = 32'd136314880;
      6244: inst = 32'd268468224;
      6245: inst = 32'd201344505;
      6246: inst = 32'd203484854;
      6247: inst = 32'd136314880;
      6248: inst = 32'd268468224;
      6249: inst = 32'd201344506;
      6250: inst = 32'd203484855;
      6251: inst = 32'd136314880;
      6252: inst = 32'd268468224;
      6253: inst = 32'd201344507;
      6254: inst = 32'd203482808;
      6255: inst = 32'd136314880;
      6256: inst = 32'd268468224;
      6257: inst = 32'd201344508;
      6258: inst = 32'd203489278;
      6259: inst = 32'd136314880;
      6260: inst = 32'd268468224;
      6261: inst = 32'd201344509;
      6262: inst = 32'd203489279;
      6263: inst = 32'd136314880;
      6264: inst = 32'd268468224;
      6265: inst = 32'd201344510;
      6266: inst = 32'd203489279;
      6267: inst = 32'd136314880;
      6268: inst = 32'd268468224;
      6269: inst = 32'd201344511;
      6270: inst = 32'd203489279;
      6271: inst = 32'd136314880;
      6272: inst = 32'd268468224;
      6273: inst = 32'd201344512;
      6274: inst = 32'd203489279;
      6275: inst = 32'd136314880;
      6276: inst = 32'd268468224;
      6277: inst = 32'd201344513;
      6278: inst = 32'd203489279;
      6279: inst = 32'd136314880;
      6280: inst = 32'd268468224;
      6281: inst = 32'd201344514;
      6282: inst = 32'd203489279;
      6283: inst = 32'd136314880;
      6284: inst = 32'd268468224;
      6285: inst = 32'd201344515;
      6286: inst = 32'd203489279;
      6287: inst = 32'd136314880;
      6288: inst = 32'd268468224;
      6289: inst = 32'd201344516;
      6290: inst = 32'd203489279;
      6291: inst = 32'd136314880;
      6292: inst = 32'd268468224;
      6293: inst = 32'd201344517;
      6294: inst = 32'd203489279;
      6295: inst = 32'd136314880;
      6296: inst = 32'd268468224;
      6297: inst = 32'd201344518;
      6298: inst = 32'd203489279;
      6299: inst = 32'd136314880;
      6300: inst = 32'd268468224;
      6301: inst = 32'd201344519;
      6302: inst = 32'd203489279;
      6303: inst = 32'd136314880;
      6304: inst = 32'd268468224;
      6305: inst = 32'd201344520;
      6306: inst = 32'd203489279;
      6307: inst = 32'd136314880;
      6308: inst = 32'd268468224;
      6309: inst = 32'd201344521;
      6310: inst = 32'd203489279;
      6311: inst = 32'd136314880;
      6312: inst = 32'd268468224;
      6313: inst = 32'd201344522;
      6314: inst = 32'd203489279;
      6315: inst = 32'd136314880;
      6316: inst = 32'd268468224;
      6317: inst = 32'd201344523;
      6318: inst = 32'd203489279;
      6319: inst = 32'd136314880;
      6320: inst = 32'd268468224;
      6321: inst = 32'd201344524;
      6322: inst = 32'd203489279;
      6323: inst = 32'd136314880;
      6324: inst = 32'd268468224;
      6325: inst = 32'd201344525;
      6326: inst = 32'd203489279;
      6327: inst = 32'd136314880;
      6328: inst = 32'd268468224;
      6329: inst = 32'd201344526;
      6330: inst = 32'd203489279;
      6331: inst = 32'd136314880;
      6332: inst = 32'd268468224;
      6333: inst = 32'd201344527;
      6334: inst = 32'd203489279;
      6335: inst = 32'd136314880;
      6336: inst = 32'd268468224;
      6337: inst = 32'd201344528;
      6338: inst = 32'd203489279;
      6339: inst = 32'd136314880;
      6340: inst = 32'd268468224;
      6341: inst = 32'd201344529;
      6342: inst = 32'd203489279;
      6343: inst = 32'd136314880;
      6344: inst = 32'd268468224;
      6345: inst = 32'd201344530;
      6346: inst = 32'd203489279;
      6347: inst = 32'd136314880;
      6348: inst = 32'd268468224;
      6349: inst = 32'd201344531;
      6350: inst = 32'd203489279;
      6351: inst = 32'd136314880;
      6352: inst = 32'd268468224;
      6353: inst = 32'd201344532;
      6354: inst = 32'd203489279;
      6355: inst = 32'd136314880;
      6356: inst = 32'd268468224;
      6357: inst = 32'd201344533;
      6358: inst = 32'd203489279;
      6359: inst = 32'd136314880;
      6360: inst = 32'd268468224;
      6361: inst = 32'd201344534;
      6362: inst = 32'd203489279;
      6363: inst = 32'd136314880;
      6364: inst = 32'd268468224;
      6365: inst = 32'd201344535;
      6366: inst = 32'd203489279;
      6367: inst = 32'd136314880;
      6368: inst = 32'd268468224;
      6369: inst = 32'd201344536;
      6370: inst = 32'd203489279;
      6371: inst = 32'd136314880;
      6372: inst = 32'd268468224;
      6373: inst = 32'd201344537;
      6374: inst = 32'd203489279;
      6375: inst = 32'd136314880;
      6376: inst = 32'd268468224;
      6377: inst = 32'd201344538;
      6378: inst = 32'd203489279;
      6379: inst = 32'd136314880;
      6380: inst = 32'd268468224;
      6381: inst = 32'd201344539;
      6382: inst = 32'd203489279;
      6383: inst = 32'd136314880;
      6384: inst = 32'd268468224;
      6385: inst = 32'd201344540;
      6386: inst = 32'd203489279;
      6387: inst = 32'd136314880;
      6388: inst = 32'd268468224;
      6389: inst = 32'd201344541;
      6390: inst = 32'd203489279;
      6391: inst = 32'd136314880;
      6392: inst = 32'd268468224;
      6393: inst = 32'd201344542;
      6394: inst = 32'd203489279;
      6395: inst = 32'd136314880;
      6396: inst = 32'd268468224;
      6397: inst = 32'd201344543;
      6398: inst = 32'd203489279;
      6399: inst = 32'd136314880;
      6400: inst = 32'd268468224;
      6401: inst = 32'd201344544;
      6402: inst = 32'd203489279;
      6403: inst = 32'd136314880;
      6404: inst = 32'd268468224;
      6405: inst = 32'd201344545;
      6406: inst = 32'd203489279;
      6407: inst = 32'd136314880;
      6408: inst = 32'd268468224;
      6409: inst = 32'd201344546;
      6410: inst = 32'd203489247;
      6411: inst = 32'd136314880;
      6412: inst = 32'd268468224;
      6413: inst = 32'd201344547;
      6414: inst = 32'd203489279;
      6415: inst = 32'd136314880;
      6416: inst = 32'd268468224;
      6417: inst = 32'd201344548;
      6418: inst = 32'd203482839;
      6419: inst = 32'd136314880;
      6420: inst = 32'd268468224;
      6421: inst = 32'd201344549;
      6422: inst = 32'd203484886;
      6423: inst = 32'd136314880;
      6424: inst = 32'd268468224;
      6425: inst = 32'd201344550;
      6426: inst = 32'd203486901;
      6427: inst = 32'd136314880;
      6428: inst = 32'd268468224;
      6429: inst = 32'd201344551;
      6430: inst = 32'd203484854;
      6431: inst = 32'd136314880;
      6432: inst = 32'd268468224;
      6433: inst = 32'd201344552;
      6434: inst = 32'd203482806;
      6435: inst = 32'd136314880;
      6436: inst = 32'd268468224;
      6437: inst = 32'd201344553;
      6438: inst = 32'd203484854;
      6439: inst = 32'd136314880;
      6440: inst = 32'd268468224;
      6441: inst = 32'd201344554;
      6442: inst = 32'd203486903;
      6443: inst = 32'd136314880;
      6444: inst = 32'd268468224;
      6445: inst = 32'd201344555;
      6446: inst = 32'd203484888;
      6447: inst = 32'd136314880;
      6448: inst = 32'd268468224;
      6449: inst = 32'd201344556;
      6450: inst = 32'd203480824;
      6451: inst = 32'd136314880;
      6452: inst = 32'd268468224;
      6453: inst = 32'd201344557;
      6454: inst = 32'd203480791;
      6455: inst = 32'd136314880;
      6456: inst = 32'd268468224;
      6457: inst = 32'd201344558;
      6458: inst = 32'd203486869;
      6459: inst = 32'd136314880;
      6460: inst = 32'd268468224;
      6461: inst = 32'd201344559;
      6462: inst = 32'd203488883;
      6463: inst = 32'd136314880;
      6464: inst = 32'd268468224;
      6465: inst = 32'd201344560;
      6466: inst = 32'd203486870;
      6467: inst = 32'd136314880;
      6468: inst = 32'd268468224;
      6469: inst = 32'd201344561;
      6470: inst = 32'd203482839;
      6471: inst = 32'd136314880;
      6472: inst = 32'd268468224;
      6473: inst = 32'd201344562;
      6474: inst = 32'd203476759;
      6475: inst = 32'd136314880;
      6476: inst = 32'd268468224;
      6477: inst = 32'd201344563;
      6478: inst = 32'd203474776;
      6479: inst = 32'd136314880;
      6480: inst = 32'd268468224;
      6481: inst = 32'd201344564;
      6482: inst = 32'd203474745;
      6483: inst = 32'd136314880;
      6484: inst = 32'd268468224;
      6485: inst = 32'd201344565;
      6486: inst = 32'd203478777;
      6487: inst = 32'd136314880;
      6488: inst = 32'd268468224;
      6489: inst = 32'd201344566;
      6490: inst = 32'd203484824;
      6491: inst = 32'd136314880;
      6492: inst = 32'd268468224;
      6493: inst = 32'd201344567;
      6494: inst = 32'd203486839;
      6495: inst = 32'd136314880;
      6496: inst = 32'd268468224;
      6497: inst = 32'd201344568;
      6498: inst = 32'd203488886;
      6499: inst = 32'd136314880;
      6500: inst = 32'd268468224;
      6501: inst = 32'd201344569;
      6502: inst = 32'd203486935;
      6503: inst = 32'd136314880;
      6504: inst = 32'd268468224;
      6505: inst = 32'd201344570;
      6506: inst = 32'd203482807;
      6507: inst = 32'd136314880;
      6508: inst = 32'd268468224;
      6509: inst = 32'd201344571;
      6510: inst = 32'd203482840;
      6511: inst = 32'd136314880;
      6512: inst = 32'd268468224;
      6513: inst = 32'd201344572;
      6514: inst = 32'd203484856;
      6515: inst = 32'd136314880;
      6516: inst = 32'd268468224;
      6517: inst = 32'd201344573;
      6518: inst = 32'd203484792;
      6519: inst = 32'd136314880;
      6520: inst = 32'd268468224;
      6521: inst = 32'd201344574;
      6522: inst = 32'd203486839;
      6523: inst = 32'd136314880;
      6524: inst = 32'd268468224;
      6525: inst = 32'd201344575;
      6526: inst = 32'd203488919;
      6527: inst = 32'd136314880;
      6528: inst = 32'd268468224;
      6529: inst = 32'd201344576;
      6530: inst = 32'd203484854;
      6531: inst = 32'd136314880;
      6532: inst = 32'd268468224;
      6533: inst = 32'd201344577;
      6534: inst = 32'd203484854;
      6535: inst = 32'd136314880;
      6536: inst = 32'd268468224;
      6537: inst = 32'd201344578;
      6538: inst = 32'd203484854;
      6539: inst = 32'd136314880;
      6540: inst = 32'd268468224;
      6541: inst = 32'd201344579;
      6542: inst = 32'd203484854;
      6543: inst = 32'd136314880;
      6544: inst = 32'd268468224;
      6545: inst = 32'd201344580;
      6546: inst = 32'd203484854;
      6547: inst = 32'd136314880;
      6548: inst = 32'd268468224;
      6549: inst = 32'd201344581;
      6550: inst = 32'd203484854;
      6551: inst = 32'd136314880;
      6552: inst = 32'd268468224;
      6553: inst = 32'd201344582;
      6554: inst = 32'd203484854;
      6555: inst = 32'd136314880;
      6556: inst = 32'd268468224;
      6557: inst = 32'd201344583;
      6558: inst = 32'd203484854;
      6559: inst = 32'd136314880;
      6560: inst = 32'd268468224;
      6561: inst = 32'd201344584;
      6562: inst = 32'd203484854;
      6563: inst = 32'd136314880;
      6564: inst = 32'd268468224;
      6565: inst = 32'd201344585;
      6566: inst = 32'd203484854;
      6567: inst = 32'd136314880;
      6568: inst = 32'd268468224;
      6569: inst = 32'd201344586;
      6570: inst = 32'd203484854;
      6571: inst = 32'd136314880;
      6572: inst = 32'd268468224;
      6573: inst = 32'd201344587;
      6574: inst = 32'd203484854;
      6575: inst = 32'd136314880;
      6576: inst = 32'd268468224;
      6577: inst = 32'd201344588;
      6578: inst = 32'd203484886;
      6579: inst = 32'd136314880;
      6580: inst = 32'd268468224;
      6581: inst = 32'd201344589;
      6582: inst = 32'd203484886;
      6583: inst = 32'd136314880;
      6584: inst = 32'd268468224;
      6585: inst = 32'd201344590;
      6586: inst = 32'd203482838;
      6587: inst = 32'd136314880;
      6588: inst = 32'd268468224;
      6589: inst = 32'd201344591;
      6590: inst = 32'd203482839;
      6591: inst = 32'd136314880;
      6592: inst = 32'd268468224;
      6593: inst = 32'd201344592;
      6594: inst = 32'd203484854;
      6595: inst = 32'd136314880;
      6596: inst = 32'd268468224;
      6597: inst = 32'd201344593;
      6598: inst = 32'd203484854;
      6599: inst = 32'd136314880;
      6600: inst = 32'd268468224;
      6601: inst = 32'd201344594;
      6602: inst = 32'd203484854;
      6603: inst = 32'd136314880;
      6604: inst = 32'd268468224;
      6605: inst = 32'd201344595;
      6606: inst = 32'd203484854;
      6607: inst = 32'd136314880;
      6608: inst = 32'd268468224;
      6609: inst = 32'd201344596;
      6610: inst = 32'd203484854;
      6611: inst = 32'd136314880;
      6612: inst = 32'd268468224;
      6613: inst = 32'd201344597;
      6614: inst = 32'd203484854;
      6615: inst = 32'd136314880;
      6616: inst = 32'd268468224;
      6617: inst = 32'd201344598;
      6618: inst = 32'd203484854;
      6619: inst = 32'd136314880;
      6620: inst = 32'd268468224;
      6621: inst = 32'd201344599;
      6622: inst = 32'd203484854;
      6623: inst = 32'd136314880;
      6624: inst = 32'd268468224;
      6625: inst = 32'd201344600;
      6626: inst = 32'd203484854;
      6627: inst = 32'd136314880;
      6628: inst = 32'd268468224;
      6629: inst = 32'd201344601;
      6630: inst = 32'd203484854;
      6631: inst = 32'd136314880;
      6632: inst = 32'd268468224;
      6633: inst = 32'd201344602;
      6634: inst = 32'd203484855;
      6635: inst = 32'd136314880;
      6636: inst = 32'd268468224;
      6637: inst = 32'd201344603;
      6638: inst = 32'd203482808;
      6639: inst = 32'd136314880;
      6640: inst = 32'd268468224;
      6641: inst = 32'd201344604;
      6642: inst = 32'd203489278;
      6643: inst = 32'd136314880;
      6644: inst = 32'd268468224;
      6645: inst = 32'd201344605;
      6646: inst = 32'd203489279;
      6647: inst = 32'd136314880;
      6648: inst = 32'd268468224;
      6649: inst = 32'd201344606;
      6650: inst = 32'd203489279;
      6651: inst = 32'd136314880;
      6652: inst = 32'd268468224;
      6653: inst = 32'd201344607;
      6654: inst = 32'd203489279;
      6655: inst = 32'd136314880;
      6656: inst = 32'd268468224;
      6657: inst = 32'd201344608;
      6658: inst = 32'd203489279;
      6659: inst = 32'd136314880;
      6660: inst = 32'd268468224;
      6661: inst = 32'd201344609;
      6662: inst = 32'd203489279;
      6663: inst = 32'd136314880;
      6664: inst = 32'd268468224;
      6665: inst = 32'd201344610;
      6666: inst = 32'd203489279;
      6667: inst = 32'd136314880;
      6668: inst = 32'd268468224;
      6669: inst = 32'd201344611;
      6670: inst = 32'd203489279;
      6671: inst = 32'd136314880;
      6672: inst = 32'd268468224;
      6673: inst = 32'd201344612;
      6674: inst = 32'd203489279;
      6675: inst = 32'd136314880;
      6676: inst = 32'd268468224;
      6677: inst = 32'd201344613;
      6678: inst = 32'd203489279;
      6679: inst = 32'd136314880;
      6680: inst = 32'd268468224;
      6681: inst = 32'd201344614;
      6682: inst = 32'd203489279;
      6683: inst = 32'd136314880;
      6684: inst = 32'd268468224;
      6685: inst = 32'd201344615;
      6686: inst = 32'd203489279;
      6687: inst = 32'd136314880;
      6688: inst = 32'd268468224;
      6689: inst = 32'd201344616;
      6690: inst = 32'd203489279;
      6691: inst = 32'd136314880;
      6692: inst = 32'd268468224;
      6693: inst = 32'd201344617;
      6694: inst = 32'd203489279;
      6695: inst = 32'd136314880;
      6696: inst = 32'd268468224;
      6697: inst = 32'd201344618;
      6698: inst = 32'd203489279;
      6699: inst = 32'd136314880;
      6700: inst = 32'd268468224;
      6701: inst = 32'd201344619;
      6702: inst = 32'd203489279;
      6703: inst = 32'd136314880;
      6704: inst = 32'd268468224;
      6705: inst = 32'd201344620;
      6706: inst = 32'd203489279;
      6707: inst = 32'd136314880;
      6708: inst = 32'd268468224;
      6709: inst = 32'd201344621;
      6710: inst = 32'd203489279;
      6711: inst = 32'd136314880;
      6712: inst = 32'd268468224;
      6713: inst = 32'd201344622;
      6714: inst = 32'd203489279;
      6715: inst = 32'd136314880;
      6716: inst = 32'd268468224;
      6717: inst = 32'd201344623;
      6718: inst = 32'd203489279;
      6719: inst = 32'd136314880;
      6720: inst = 32'd268468224;
      6721: inst = 32'd201344624;
      6722: inst = 32'd203489279;
      6723: inst = 32'd136314880;
      6724: inst = 32'd268468224;
      6725: inst = 32'd201344625;
      6726: inst = 32'd203489279;
      6727: inst = 32'd136314880;
      6728: inst = 32'd268468224;
      6729: inst = 32'd201344626;
      6730: inst = 32'd203489279;
      6731: inst = 32'd136314880;
      6732: inst = 32'd268468224;
      6733: inst = 32'd201344627;
      6734: inst = 32'd203489279;
      6735: inst = 32'd136314880;
      6736: inst = 32'd268468224;
      6737: inst = 32'd201344628;
      6738: inst = 32'd203489279;
      6739: inst = 32'd136314880;
      6740: inst = 32'd268468224;
      6741: inst = 32'd201344629;
      6742: inst = 32'd203489279;
      6743: inst = 32'd136314880;
      6744: inst = 32'd268468224;
      6745: inst = 32'd201344630;
      6746: inst = 32'd203489279;
      6747: inst = 32'd136314880;
      6748: inst = 32'd268468224;
      6749: inst = 32'd201344631;
      6750: inst = 32'd203489279;
      6751: inst = 32'd136314880;
      6752: inst = 32'd268468224;
      6753: inst = 32'd201344632;
      6754: inst = 32'd203489279;
      6755: inst = 32'd136314880;
      6756: inst = 32'd268468224;
      6757: inst = 32'd201344633;
      6758: inst = 32'd203489279;
      6759: inst = 32'd136314880;
      6760: inst = 32'd268468224;
      6761: inst = 32'd201344634;
      6762: inst = 32'd203489279;
      6763: inst = 32'd136314880;
      6764: inst = 32'd268468224;
      6765: inst = 32'd201344635;
      6766: inst = 32'd203489279;
      6767: inst = 32'd136314880;
      6768: inst = 32'd268468224;
      6769: inst = 32'd201344636;
      6770: inst = 32'd203489279;
      6771: inst = 32'd136314880;
      6772: inst = 32'd268468224;
      6773: inst = 32'd201344637;
      6774: inst = 32'd203489279;
      6775: inst = 32'd136314880;
      6776: inst = 32'd268468224;
      6777: inst = 32'd201344638;
      6778: inst = 32'd203489279;
      6779: inst = 32'd136314880;
      6780: inst = 32'd268468224;
      6781: inst = 32'd201344639;
      6782: inst = 32'd203489279;
      6783: inst = 32'd136314880;
      6784: inst = 32'd268468224;
      6785: inst = 32'd201344640;
      6786: inst = 32'd203489279;
      6787: inst = 32'd136314880;
      6788: inst = 32'd268468224;
      6789: inst = 32'd201344641;
      6790: inst = 32'd203489279;
      6791: inst = 32'd136314880;
      6792: inst = 32'd268468224;
      6793: inst = 32'd201344642;
      6794: inst = 32'd203489247;
      6795: inst = 32'd136314880;
      6796: inst = 32'd268468224;
      6797: inst = 32'd201344643;
      6798: inst = 32'd203489279;
      6799: inst = 32'd136314880;
      6800: inst = 32'd268468224;
      6801: inst = 32'd201344644;
      6802: inst = 32'd203482839;
      6803: inst = 32'd136314880;
      6804: inst = 32'd268468224;
      6805: inst = 32'd201344645;
      6806: inst = 32'd203484886;
      6807: inst = 32'd136314880;
      6808: inst = 32'd268468224;
      6809: inst = 32'd201344646;
      6810: inst = 32'd203486901;
      6811: inst = 32'd136314880;
      6812: inst = 32'd268468224;
      6813: inst = 32'd201344647;
      6814: inst = 32'd203484854;
      6815: inst = 32'd136314880;
      6816: inst = 32'd268468224;
      6817: inst = 32'd201344648;
      6818: inst = 32'd203484854;
      6819: inst = 32'd136314880;
      6820: inst = 32'd268468224;
      6821: inst = 32'd201344649;
      6822: inst = 32'd203484887;
      6823: inst = 32'd136314880;
      6824: inst = 32'd268468224;
      6825: inst = 32'd201344650;
      6826: inst = 32'd203486902;
      6827: inst = 32'd136314880;
      6828: inst = 32'd268468224;
      6829: inst = 32'd201344651;
      6830: inst = 32'd203484823;
      6831: inst = 32'd136314880;
      6832: inst = 32'd268468224;
      6833: inst = 32'd201344652;
      6834: inst = 32'd203478711;
      6835: inst = 32'd136314880;
      6836: inst = 32'd268468224;
      6837: inst = 32'd201344653;
      6838: inst = 32'd203482871;
      6839: inst = 32'd136314880;
      6840: inst = 32'd268468224;
      6841: inst = 32'd201344654;
      6842: inst = 32'd203488982;
      6843: inst = 32'd136314880;
      6844: inst = 32'd268468224;
      6845: inst = 32'd201344655;
      6846: inst = 32'd203488786;
      6847: inst = 32'd136314880;
      6848: inst = 32'd268468224;
      6849: inst = 32'd201344656;
      6850: inst = 32'd203488883;
      6851: inst = 32'd136314880;
      6852: inst = 32'd268468224;
      6853: inst = 32'd201344657;
      6854: inst = 32'd203488884;
      6855: inst = 32'd136314880;
      6856: inst = 32'd268468224;
      6857: inst = 32'd201344658;
      6858: inst = 32'd203488948;
      6859: inst = 32'd136314880;
      6860: inst = 32'd268468224;
      6861: inst = 32'd201344659;
      6862: inst = 32'd203486900;
      6863: inst = 32'd136314880;
      6864: inst = 32'd268468224;
      6865: inst = 32'd201344660;
      6866: inst = 32'd203486901;
      6867: inst = 32'd136314880;
      6868: inst = 32'd268468224;
      6869: inst = 32'd201344661;
      6870: inst = 32'd203488917;
      6871: inst = 32'd136314880;
      6872: inst = 32'd268468224;
      6873: inst = 32'd201344662;
      6874: inst = 32'd203488885;
      6875: inst = 32'd136314880;
      6876: inst = 32'd268468224;
      6877: inst = 32'd201344663;
      6878: inst = 32'd203488884;
      6879: inst = 32'd136314880;
      6880: inst = 32'd268468224;
      6881: inst = 32'd201344664;
      6882: inst = 32'd203488883;
      6883: inst = 32'd136314880;
      6884: inst = 32'd268468224;
      6885: inst = 32'd201344665;
      6886: inst = 32'd203488947;
      6887: inst = 32'd136314880;
      6888: inst = 32'd268468224;
      6889: inst = 32'd201344666;
      6890: inst = 32'd203488915;
      6891: inst = 32'd136314880;
      6892: inst = 32'd268468224;
      6893: inst = 32'd201344667;
      6894: inst = 32'd203488916;
      6895: inst = 32'd136314880;
      6896: inst = 32'd268468224;
      6897: inst = 32'd201344668;
      6898: inst = 32'd203488917;
      6899: inst = 32'd136314880;
      6900: inst = 32'd268468224;
      6901: inst = 32'd201344669;
      6902: inst = 32'd203488884;
      6903: inst = 32'd136314880;
      6904: inst = 32'd268468224;
      6905: inst = 32'd201344670;
      6906: inst = 32'd203488916;
      6907: inst = 32'd136314880;
      6908: inst = 32'd268468224;
      6909: inst = 32'd201344671;
      6910: inst = 32'd203488916;
      6911: inst = 32'd136314880;
      6912: inst = 32'd268468224;
      6913: inst = 32'd201344672;
      6914: inst = 32'd203484854;
      6915: inst = 32'd136314880;
      6916: inst = 32'd268468224;
      6917: inst = 32'd201344673;
      6918: inst = 32'd203484854;
      6919: inst = 32'd136314880;
      6920: inst = 32'd268468224;
      6921: inst = 32'd201344674;
      6922: inst = 32'd203484854;
      6923: inst = 32'd136314880;
      6924: inst = 32'd268468224;
      6925: inst = 32'd201344675;
      6926: inst = 32'd203484854;
      6927: inst = 32'd136314880;
      6928: inst = 32'd268468224;
      6929: inst = 32'd201344676;
      6930: inst = 32'd203484854;
      6931: inst = 32'd136314880;
      6932: inst = 32'd268468224;
      6933: inst = 32'd201344677;
      6934: inst = 32'd203484854;
      6935: inst = 32'd136314880;
      6936: inst = 32'd268468224;
      6937: inst = 32'd201344678;
      6938: inst = 32'd203484854;
      6939: inst = 32'd136314880;
      6940: inst = 32'd268468224;
      6941: inst = 32'd201344679;
      6942: inst = 32'd203484854;
      6943: inst = 32'd136314880;
      6944: inst = 32'd268468224;
      6945: inst = 32'd201344680;
      6946: inst = 32'd203484854;
      6947: inst = 32'd136314880;
      6948: inst = 32'd268468224;
      6949: inst = 32'd201344681;
      6950: inst = 32'd203484854;
      6951: inst = 32'd136314880;
      6952: inst = 32'd268468224;
      6953: inst = 32'd201344682;
      6954: inst = 32'd203484854;
      6955: inst = 32'd136314880;
      6956: inst = 32'd268468224;
      6957: inst = 32'd201344683;
      6958: inst = 32'd203484854;
      6959: inst = 32'd136314880;
      6960: inst = 32'd268468224;
      6961: inst = 32'd201344684;
      6962: inst = 32'd203484854;
      6963: inst = 32'd136314880;
      6964: inst = 32'd268468224;
      6965: inst = 32'd201344685;
      6966: inst = 32'd203484854;
      6967: inst = 32'd136314880;
      6968: inst = 32'd268468224;
      6969: inst = 32'd201344686;
      6970: inst = 32'd203484886;
      6971: inst = 32'd136314880;
      6972: inst = 32'd268468224;
      6973: inst = 32'd201344687;
      6974: inst = 32'd203484855;
      6975: inst = 32'd136314880;
      6976: inst = 32'd268468224;
      6977: inst = 32'd201344688;
      6978: inst = 32'd203484854;
      6979: inst = 32'd136314880;
      6980: inst = 32'd268468224;
      6981: inst = 32'd201344689;
      6982: inst = 32'd203484854;
      6983: inst = 32'd136314880;
      6984: inst = 32'd268468224;
      6985: inst = 32'd201344690;
      6986: inst = 32'd203484854;
      6987: inst = 32'd136314880;
      6988: inst = 32'd268468224;
      6989: inst = 32'd201344691;
      6990: inst = 32'd203484854;
      6991: inst = 32'd136314880;
      6992: inst = 32'd268468224;
      6993: inst = 32'd201344692;
      6994: inst = 32'd203484854;
      6995: inst = 32'd136314880;
      6996: inst = 32'd268468224;
      6997: inst = 32'd201344693;
      6998: inst = 32'd203484854;
      6999: inst = 32'd136314880;
      7000: inst = 32'd268468224;
      7001: inst = 32'd201344694;
      7002: inst = 32'd203484854;
      7003: inst = 32'd136314880;
      7004: inst = 32'd268468224;
      7005: inst = 32'd201344695;
      7006: inst = 32'd203484854;
      7007: inst = 32'd136314880;
      7008: inst = 32'd268468224;
      7009: inst = 32'd201344696;
      7010: inst = 32'd203484854;
      7011: inst = 32'd136314880;
      7012: inst = 32'd268468224;
      7013: inst = 32'd201344697;
      7014: inst = 32'd203484854;
      7015: inst = 32'd136314880;
      7016: inst = 32'd268468224;
      7017: inst = 32'd201344698;
      7018: inst = 32'd203484855;
      7019: inst = 32'd136314880;
      7020: inst = 32'd268468224;
      7021: inst = 32'd201344699;
      7022: inst = 32'd203482808;
      7023: inst = 32'd136314880;
      7024: inst = 32'd268468224;
      7025: inst = 32'd201344700;
      7026: inst = 32'd203489278;
      7027: inst = 32'd136314880;
      7028: inst = 32'd268468224;
      7029: inst = 32'd201344701;
      7030: inst = 32'd203489279;
      7031: inst = 32'd136314880;
      7032: inst = 32'd268468224;
      7033: inst = 32'd201344702;
      7034: inst = 32'd203489279;
      7035: inst = 32'd136314880;
      7036: inst = 32'd268468224;
      7037: inst = 32'd201344703;
      7038: inst = 32'd203489279;
      7039: inst = 32'd136314880;
      7040: inst = 32'd268468224;
      7041: inst = 32'd201344704;
      7042: inst = 32'd203489279;
      7043: inst = 32'd136314880;
      7044: inst = 32'd268468224;
      7045: inst = 32'd201344705;
      7046: inst = 32'd203489279;
      7047: inst = 32'd136314880;
      7048: inst = 32'd268468224;
      7049: inst = 32'd201344706;
      7050: inst = 32'd203489279;
      7051: inst = 32'd136314880;
      7052: inst = 32'd268468224;
      7053: inst = 32'd201344707;
      7054: inst = 32'd203489279;
      7055: inst = 32'd136314880;
      7056: inst = 32'd268468224;
      7057: inst = 32'd201344708;
      7058: inst = 32'd203489279;
      7059: inst = 32'd136314880;
      7060: inst = 32'd268468224;
      7061: inst = 32'd201344709;
      7062: inst = 32'd203489279;
      7063: inst = 32'd136314880;
      7064: inst = 32'd268468224;
      7065: inst = 32'd201344710;
      7066: inst = 32'd203489279;
      7067: inst = 32'd136314880;
      7068: inst = 32'd268468224;
      7069: inst = 32'd201344711;
      7070: inst = 32'd203489279;
      7071: inst = 32'd136314880;
      7072: inst = 32'd268468224;
      7073: inst = 32'd201344712;
      7074: inst = 32'd203489279;
      7075: inst = 32'd136314880;
      7076: inst = 32'd268468224;
      7077: inst = 32'd201344713;
      7078: inst = 32'd203489279;
      7079: inst = 32'd136314880;
      7080: inst = 32'd268468224;
      7081: inst = 32'd201344714;
      7082: inst = 32'd203489279;
      7083: inst = 32'd136314880;
      7084: inst = 32'd268468224;
      7085: inst = 32'd201344715;
      7086: inst = 32'd203489279;
      7087: inst = 32'd136314880;
      7088: inst = 32'd268468224;
      7089: inst = 32'd201344716;
      7090: inst = 32'd203489279;
      7091: inst = 32'd136314880;
      7092: inst = 32'd268468224;
      7093: inst = 32'd201344717;
      7094: inst = 32'd203489279;
      7095: inst = 32'd136314880;
      7096: inst = 32'd268468224;
      7097: inst = 32'd201344718;
      7098: inst = 32'd203489279;
      7099: inst = 32'd136314880;
      7100: inst = 32'd268468224;
      7101: inst = 32'd201344719;
      7102: inst = 32'd203489279;
      7103: inst = 32'd136314880;
      7104: inst = 32'd268468224;
      7105: inst = 32'd201344720;
      7106: inst = 32'd203489279;
      7107: inst = 32'd136314880;
      7108: inst = 32'd268468224;
      7109: inst = 32'd201344721;
      7110: inst = 32'd203489279;
      7111: inst = 32'd136314880;
      7112: inst = 32'd268468224;
      7113: inst = 32'd201344722;
      7114: inst = 32'd203489279;
      7115: inst = 32'd136314880;
      7116: inst = 32'd268468224;
      7117: inst = 32'd201344723;
      7118: inst = 32'd203489279;
      7119: inst = 32'd136314880;
      7120: inst = 32'd268468224;
      7121: inst = 32'd201344724;
      7122: inst = 32'd203489279;
      7123: inst = 32'd136314880;
      7124: inst = 32'd268468224;
      7125: inst = 32'd201344725;
      7126: inst = 32'd203489279;
      7127: inst = 32'd136314880;
      7128: inst = 32'd268468224;
      7129: inst = 32'd201344726;
      7130: inst = 32'd203489279;
      7131: inst = 32'd136314880;
      7132: inst = 32'd268468224;
      7133: inst = 32'd201344727;
      7134: inst = 32'd203489279;
      7135: inst = 32'd136314880;
      7136: inst = 32'd268468224;
      7137: inst = 32'd201344728;
      7138: inst = 32'd203489279;
      7139: inst = 32'd136314880;
      7140: inst = 32'd268468224;
      7141: inst = 32'd201344729;
      7142: inst = 32'd203489279;
      7143: inst = 32'd136314880;
      7144: inst = 32'd268468224;
      7145: inst = 32'd201344730;
      7146: inst = 32'd203489279;
      7147: inst = 32'd136314880;
      7148: inst = 32'd268468224;
      7149: inst = 32'd201344731;
      7150: inst = 32'd203489279;
      7151: inst = 32'd136314880;
      7152: inst = 32'd268468224;
      7153: inst = 32'd201344732;
      7154: inst = 32'd203489279;
      7155: inst = 32'd136314880;
      7156: inst = 32'd268468224;
      7157: inst = 32'd201344733;
      7158: inst = 32'd203489279;
      7159: inst = 32'd136314880;
      7160: inst = 32'd268468224;
      7161: inst = 32'd201344734;
      7162: inst = 32'd203489279;
      7163: inst = 32'd136314880;
      7164: inst = 32'd268468224;
      7165: inst = 32'd201344735;
      7166: inst = 32'd203489279;
      7167: inst = 32'd136314880;
      7168: inst = 32'd268468224;
      7169: inst = 32'd201344736;
      7170: inst = 32'd203489279;
      7171: inst = 32'd136314880;
      7172: inst = 32'd268468224;
      7173: inst = 32'd201344737;
      7174: inst = 32'd203489279;
      7175: inst = 32'd136314880;
      7176: inst = 32'd268468224;
      7177: inst = 32'd201344738;
      7178: inst = 32'd203489247;
      7179: inst = 32'd136314880;
      7180: inst = 32'd268468224;
      7181: inst = 32'd201344739;
      7182: inst = 32'd203489279;
      7183: inst = 32'd136314880;
      7184: inst = 32'd268468224;
      7185: inst = 32'd201344740;
      7186: inst = 32'd203482839;
      7187: inst = 32'd136314880;
      7188: inst = 32'd268468224;
      7189: inst = 32'd201344741;
      7190: inst = 32'd203484886;
      7191: inst = 32'd136314880;
      7192: inst = 32'd268468224;
      7193: inst = 32'd201344742;
      7194: inst = 32'd203486901;
      7195: inst = 32'd136314880;
      7196: inst = 32'd268468224;
      7197: inst = 32'd201344743;
      7198: inst = 32'd203484854;
      7199: inst = 32'd136314880;
      7200: inst = 32'd268468224;
      7201: inst = 32'd201344744;
      7202: inst = 32'd203482806;
      7203: inst = 32'd136314880;
      7204: inst = 32'd268468224;
      7205: inst = 32'd201344745;
      7206: inst = 32'd203486934;
      7207: inst = 32'd136314880;
      7208: inst = 32'd268468224;
      7209: inst = 32'd201344746;
      7210: inst = 32'd203486870;
      7211: inst = 32'd136314880;
      7212: inst = 32'd268468224;
      7213: inst = 32'd201344747;
      7214: inst = 32'd203484855;
      7215: inst = 32'd136314880;
      7216: inst = 32'd268468224;
      7217: inst = 32'd201344748;
      7218: inst = 32'd203482872;
      7219: inst = 32'd136314880;
      7220: inst = 32'd268468224;
      7221: inst = 32'd201344749;
      7222: inst = 32'd203482871;
      7223: inst = 32'd136314880;
      7224: inst = 32'd268468224;
      7225: inst = 32'd201344750;
      7226: inst = 32'd203484723;
      7227: inst = 32'd136314880;
      7228: inst = 32'd268468224;
      7229: inst = 32'd201344751;
      7230: inst = 32'd203471752;
      7231: inst = 32'd136314880;
      7232: inst = 32'd268468224;
      7233: inst = 32'd201344752;
      7234: inst = 32'd203471588;
      7235: inst = 32'd136314880;
      7236: inst = 32'd268468224;
      7237: inst = 32'd201344753;
      7238: inst = 32'd203471587;
      7239: inst = 32'd136314880;
      7240: inst = 32'd268468224;
      7241: inst = 32'd201344754;
      7242: inst = 32'd203471587;
      7243: inst = 32'd136314880;
      7244: inst = 32'd268468224;
      7245: inst = 32'd201344755;
      7246: inst = 32'd203471587;
      7247: inst = 32'd136314880;
      7248: inst = 32'd268468224;
      7249: inst = 32'd201344756;
      7250: inst = 32'd203471587;
      7251: inst = 32'd136314880;
      7252: inst = 32'd268468224;
      7253: inst = 32'd201344757;
      7254: inst = 32'd203471587;
      7255: inst = 32'd136314880;
      7256: inst = 32'd268468224;
      7257: inst = 32'd201344758;
      7258: inst = 32'd203469572;
      7259: inst = 32'd136314880;
      7260: inst = 32'd268468224;
      7261: inst = 32'd201344759;
      7262: inst = 32'd203469572;
      7263: inst = 32'd136314880;
      7264: inst = 32'd268468224;
      7265: inst = 32'd201344760;
      7266: inst = 32'd203467523;
      7267: inst = 32'd136314880;
      7268: inst = 32'd268468224;
      7269: inst = 32'd201344761;
      7270: inst = 32'd203469604;
      7271: inst = 32'd136314880;
      7272: inst = 32'd268468224;
      7273: inst = 32'd201344762;
      7274: inst = 32'd203467523;
      7275: inst = 32'd136314880;
      7276: inst = 32'd268468224;
      7277: inst = 32'd201344763;
      7278: inst = 32'd203467523;
      7279: inst = 32'd136314880;
      7280: inst = 32'd268468224;
      7281: inst = 32'd201344764;
      7282: inst = 32'd203469604;
      7283: inst = 32'd136314880;
      7284: inst = 32'd268468224;
      7285: inst = 32'd201344765;
      7286: inst = 32'd203467556;
      7287: inst = 32'd136314880;
      7288: inst = 32'd268468224;
      7289: inst = 32'd201344766;
      7290: inst = 32'd203467588;
      7291: inst = 32'd136314880;
      7292: inst = 32'd268468224;
      7293: inst = 32'd201344767;
      7294: inst = 32'd203465474;
      7295: inst = 32'd136314880;
      7296: inst = 32'd268468224;
      7297: inst = 32'd201344768;
      7298: inst = 32'd203484854;
      7299: inst = 32'd136314880;
      7300: inst = 32'd268468224;
      7301: inst = 32'd201344769;
      7302: inst = 32'd203484854;
      7303: inst = 32'd136314880;
      7304: inst = 32'd268468224;
      7305: inst = 32'd201344770;
      7306: inst = 32'd203484854;
      7307: inst = 32'd136314880;
      7308: inst = 32'd268468224;
      7309: inst = 32'd201344771;
      7310: inst = 32'd203484855;
      7311: inst = 32'd136314880;
      7312: inst = 32'd268468224;
      7313: inst = 32'd201344772;
      7314: inst = 32'd203484855;
      7315: inst = 32'd136314880;
      7316: inst = 32'd268468224;
      7317: inst = 32'd201344773;
      7318: inst = 32'd203484855;
      7319: inst = 32'd136314880;
      7320: inst = 32'd268468224;
      7321: inst = 32'd201344774;
      7322: inst = 32'd203484854;
      7323: inst = 32'd136314880;
      7324: inst = 32'd268468224;
      7325: inst = 32'd201344775;
      7326: inst = 32'd203484854;
      7327: inst = 32'd136314880;
      7328: inst = 32'd268468224;
      7329: inst = 32'd201344776;
      7330: inst = 32'd203484854;
      7331: inst = 32'd136314880;
      7332: inst = 32'd268468224;
      7333: inst = 32'd201344777;
      7334: inst = 32'd203484854;
      7335: inst = 32'd136314880;
      7336: inst = 32'd268468224;
      7337: inst = 32'd201344778;
      7338: inst = 32'd203484854;
      7339: inst = 32'd136314880;
      7340: inst = 32'd268468224;
      7341: inst = 32'd201344779;
      7342: inst = 32'd203484854;
      7343: inst = 32'd136314880;
      7344: inst = 32'd268468224;
      7345: inst = 32'd201344780;
      7346: inst = 32'd203484854;
      7347: inst = 32'd136314880;
      7348: inst = 32'd268468224;
      7349: inst = 32'd201344781;
      7350: inst = 32'd203484854;
      7351: inst = 32'd136314880;
      7352: inst = 32'd268468224;
      7353: inst = 32'd201344782;
      7354: inst = 32'd203484854;
      7355: inst = 32'd136314880;
      7356: inst = 32'd268468224;
      7357: inst = 32'd201344783;
      7358: inst = 32'd203484854;
      7359: inst = 32'd136314880;
      7360: inst = 32'd268468224;
      7361: inst = 32'd201344784;
      7362: inst = 32'd203484854;
      7363: inst = 32'd136314880;
      7364: inst = 32'd268468224;
      7365: inst = 32'd201344785;
      7366: inst = 32'd203484854;
      7367: inst = 32'd136314880;
      7368: inst = 32'd268468224;
      7369: inst = 32'd201344786;
      7370: inst = 32'd203484854;
      7371: inst = 32'd136314880;
      7372: inst = 32'd268468224;
      7373: inst = 32'd201344787;
      7374: inst = 32'd203484854;
      7375: inst = 32'd136314880;
      7376: inst = 32'd268468224;
      7377: inst = 32'd201344788;
      7378: inst = 32'd203484854;
      7379: inst = 32'd136314880;
      7380: inst = 32'd268468224;
      7381: inst = 32'd201344789;
      7382: inst = 32'd203484854;
      7383: inst = 32'd136314880;
      7384: inst = 32'd268468224;
      7385: inst = 32'd201344790;
      7386: inst = 32'd203484854;
      7387: inst = 32'd136314880;
      7388: inst = 32'd268468224;
      7389: inst = 32'd201344791;
      7390: inst = 32'd203484854;
      7391: inst = 32'd136314880;
      7392: inst = 32'd268468224;
      7393: inst = 32'd201344792;
      7394: inst = 32'd203484854;
      7395: inst = 32'd136314880;
      7396: inst = 32'd268468224;
      7397: inst = 32'd201344793;
      7398: inst = 32'd203484854;
      7399: inst = 32'd136314880;
      7400: inst = 32'd268468224;
      7401: inst = 32'd201344794;
      7402: inst = 32'd203484855;
      7403: inst = 32'd136314880;
      7404: inst = 32'd268468224;
      7405: inst = 32'd201344795;
      7406: inst = 32'd203482808;
      7407: inst = 32'd136314880;
      7408: inst = 32'd268468224;
      7409: inst = 32'd201344796;
      7410: inst = 32'd203489278;
      7411: inst = 32'd136314880;
      7412: inst = 32'd268468224;
      7413: inst = 32'd201344797;
      7414: inst = 32'd203489279;
      7415: inst = 32'd136314880;
      7416: inst = 32'd268468224;
      7417: inst = 32'd201344798;
      7418: inst = 32'd203489279;
      7419: inst = 32'd136314880;
      7420: inst = 32'd268468224;
      7421: inst = 32'd201344799;
      7422: inst = 32'd203489279;
      7423: inst = 32'd136314880;
      7424: inst = 32'd268468224;
      7425: inst = 32'd201344800;
      7426: inst = 32'd203489279;
      7427: inst = 32'd136314880;
      7428: inst = 32'd268468224;
      7429: inst = 32'd201344801;
      7430: inst = 32'd203489279;
      7431: inst = 32'd136314880;
      7432: inst = 32'd268468224;
      7433: inst = 32'd201344802;
      7434: inst = 32'd203489279;
      7435: inst = 32'd136314880;
      7436: inst = 32'd268468224;
      7437: inst = 32'd201344803;
      7438: inst = 32'd203489279;
      7439: inst = 32'd136314880;
      7440: inst = 32'd268468224;
      7441: inst = 32'd201344804;
      7442: inst = 32'd203489279;
      7443: inst = 32'd136314880;
      7444: inst = 32'd268468224;
      7445: inst = 32'd201344805;
      7446: inst = 32'd203489279;
      7447: inst = 32'd136314880;
      7448: inst = 32'd268468224;
      7449: inst = 32'd201344806;
      7450: inst = 32'd203489279;
      7451: inst = 32'd136314880;
      7452: inst = 32'd268468224;
      7453: inst = 32'd201344807;
      7454: inst = 32'd203489279;
      7455: inst = 32'd136314880;
      7456: inst = 32'd268468224;
      7457: inst = 32'd201344808;
      7458: inst = 32'd203489279;
      7459: inst = 32'd136314880;
      7460: inst = 32'd268468224;
      7461: inst = 32'd201344809;
      7462: inst = 32'd203489279;
      7463: inst = 32'd136314880;
      7464: inst = 32'd268468224;
      7465: inst = 32'd201344810;
      7466: inst = 32'd203489279;
      7467: inst = 32'd136314880;
      7468: inst = 32'd268468224;
      7469: inst = 32'd201344811;
      7470: inst = 32'd203489279;
      7471: inst = 32'd136314880;
      7472: inst = 32'd268468224;
      7473: inst = 32'd201344812;
      7474: inst = 32'd203489279;
      7475: inst = 32'd136314880;
      7476: inst = 32'd268468224;
      7477: inst = 32'd201344813;
      7478: inst = 32'd203489279;
      7479: inst = 32'd136314880;
      7480: inst = 32'd268468224;
      7481: inst = 32'd201344814;
      7482: inst = 32'd203489279;
      7483: inst = 32'd136314880;
      7484: inst = 32'd268468224;
      7485: inst = 32'd201344815;
      7486: inst = 32'd203489279;
      7487: inst = 32'd136314880;
      7488: inst = 32'd268468224;
      7489: inst = 32'd201344816;
      7490: inst = 32'd203489279;
      7491: inst = 32'd136314880;
      7492: inst = 32'd268468224;
      7493: inst = 32'd201344817;
      7494: inst = 32'd203489279;
      7495: inst = 32'd136314880;
      7496: inst = 32'd268468224;
      7497: inst = 32'd201344818;
      7498: inst = 32'd203489279;
      7499: inst = 32'd136314880;
      7500: inst = 32'd268468224;
      7501: inst = 32'd201344819;
      7502: inst = 32'd203489279;
      7503: inst = 32'd136314880;
      7504: inst = 32'd268468224;
      7505: inst = 32'd201344820;
      7506: inst = 32'd203489279;
      7507: inst = 32'd136314880;
      7508: inst = 32'd268468224;
      7509: inst = 32'd201344821;
      7510: inst = 32'd203489279;
      7511: inst = 32'd136314880;
      7512: inst = 32'd268468224;
      7513: inst = 32'd201344822;
      7514: inst = 32'd203489279;
      7515: inst = 32'd136314880;
      7516: inst = 32'd268468224;
      7517: inst = 32'd201344823;
      7518: inst = 32'd203489279;
      7519: inst = 32'd136314880;
      7520: inst = 32'd268468224;
      7521: inst = 32'd201344824;
      7522: inst = 32'd203489279;
      7523: inst = 32'd136314880;
      7524: inst = 32'd268468224;
      7525: inst = 32'd201344825;
      7526: inst = 32'd203489279;
      7527: inst = 32'd136314880;
      7528: inst = 32'd268468224;
      7529: inst = 32'd201344826;
      7530: inst = 32'd203489279;
      7531: inst = 32'd136314880;
      7532: inst = 32'd268468224;
      7533: inst = 32'd201344827;
      7534: inst = 32'd203489279;
      7535: inst = 32'd136314880;
      7536: inst = 32'd268468224;
      7537: inst = 32'd201344828;
      7538: inst = 32'd203489279;
      7539: inst = 32'd136314880;
      7540: inst = 32'd268468224;
      7541: inst = 32'd201344829;
      7542: inst = 32'd203489279;
      7543: inst = 32'd136314880;
      7544: inst = 32'd268468224;
      7545: inst = 32'd201344830;
      7546: inst = 32'd203489279;
      7547: inst = 32'd136314880;
      7548: inst = 32'd268468224;
      7549: inst = 32'd201344831;
      7550: inst = 32'd203489279;
      7551: inst = 32'd136314880;
      7552: inst = 32'd268468224;
      7553: inst = 32'd201344832;
      7554: inst = 32'd203489279;
      7555: inst = 32'd136314880;
      7556: inst = 32'd268468224;
      7557: inst = 32'd201344833;
      7558: inst = 32'd203489279;
      7559: inst = 32'd136314880;
      7560: inst = 32'd268468224;
      7561: inst = 32'd201344834;
      7562: inst = 32'd203489247;
      7563: inst = 32'd136314880;
      7564: inst = 32'd268468224;
      7565: inst = 32'd201344835;
      7566: inst = 32'd203489279;
      7567: inst = 32'd136314880;
      7568: inst = 32'd268468224;
      7569: inst = 32'd201344836;
      7570: inst = 32'd203482840;
      7571: inst = 32'd136314880;
      7572: inst = 32'd268468224;
      7573: inst = 32'd201344837;
      7574: inst = 32'd203484886;
      7575: inst = 32'd136314880;
      7576: inst = 32'd268468224;
      7577: inst = 32'd201344838;
      7578: inst = 32'd203486869;
      7579: inst = 32'd136314880;
      7580: inst = 32'd268468224;
      7581: inst = 32'd201344839;
      7582: inst = 32'd203484854;
      7583: inst = 32'd136314880;
      7584: inst = 32'd268468224;
      7585: inst = 32'd201344840;
      7586: inst = 32'd203484886;
      7587: inst = 32'd136314880;
      7588: inst = 32'd268468224;
      7589: inst = 32'd201344841;
      7590: inst = 32'd203486934;
      7591: inst = 32'd136314880;
      7592: inst = 32'd268468224;
      7593: inst = 32'd201344842;
      7594: inst = 32'd203484789;
      7595: inst = 32'd136314880;
      7596: inst = 32'd268468224;
      7597: inst = 32'd201344843;
      7598: inst = 32'd203484855;
      7599: inst = 32'd136314880;
      7600: inst = 32'd268468224;
      7601: inst = 32'd201344844;
      7602: inst = 32'd203482872;
      7603: inst = 32'd136314880;
      7604: inst = 32'd268468224;
      7605: inst = 32'd201344845;
      7606: inst = 32'd203484952;
      7607: inst = 32'd136314880;
      7608: inst = 32'd268468224;
      7609: inst = 32'd201344846;
      7610: inst = 32'd203486836;
      7611: inst = 32'd136314880;
      7612: inst = 32'd268468224;
      7613: inst = 32'd201344847;
      7614: inst = 32'd203465413;
      7615: inst = 32'd136314880;
      7616: inst = 32'd268468224;
      7617: inst = 32'd201344848;
      7618: inst = 32'd203480006;
      7619: inst = 32'd136314880;
      7620: inst = 32'd268468224;
      7621: inst = 32'd201344849;
      7622: inst = 32'd203480005;
      7623: inst = 32'd136314880;
      7624: inst = 32'd268468224;
      7625: inst = 32'd201344850;
      7626: inst = 32'd203482053;
      7627: inst = 32'd136314880;
      7628: inst = 32'd268468224;
      7629: inst = 32'd201344851;
      7630: inst = 32'd203482052;
      7631: inst = 32'd136314880;
      7632: inst = 32'd268468224;
      7633: inst = 32'd201344852;
      7634: inst = 32'd203482051;
      7635: inst = 32'd136314880;
      7636: inst = 32'd268468224;
      7637: inst = 32'd201344853;
      7638: inst = 32'd203480004;
      7639: inst = 32'd136314880;
      7640: inst = 32'd268468224;
      7641: inst = 32'd201344854;
      7642: inst = 32'd203480005;
      7643: inst = 32'd136314880;
      7644: inst = 32'd268468224;
      7645: inst = 32'd201344855;
      7646: inst = 32'd203480006;
      7647: inst = 32'd136314880;
      7648: inst = 32'd268468224;
      7649: inst = 32'd201344856;
      7650: inst = 32'd203482054;
      7651: inst = 32'd136314880;
      7652: inst = 32'd268468224;
      7653: inst = 32'd201344857;
      7654: inst = 32'd203482087;
      7655: inst = 32'd136314880;
      7656: inst = 32'd268468224;
      7657: inst = 32'd201344858;
      7658: inst = 32'd203477958;
      7659: inst = 32'd136314880;
      7660: inst = 32'd268468224;
      7661: inst = 32'd201344859;
      7662: inst = 32'd203477989;
      7663: inst = 32'd136314880;
      7664: inst = 32'd268468224;
      7665: inst = 32'd201344860;
      7666: inst = 32'd203478021;
      7667: inst = 32'd136314880;
      7668: inst = 32'd268468224;
      7669: inst = 32'd201344861;
      7670: inst = 32'd203477989;
      7671: inst = 32'd136314880;
      7672: inst = 32'd268468224;
      7673: inst = 32'd201344862;
      7674: inst = 32'd203479973;
      7675: inst = 32'd136314880;
      7676: inst = 32'd268468224;
      7677: inst = 32'd201344863;
      7678: inst = 32'd203477795;
      7679: inst = 32'd136314880;
      7680: inst = 32'd268468224;
      7681: inst = 32'd201344864;
      7682: inst = 32'd203484854;
      7683: inst = 32'd136314880;
      7684: inst = 32'd268468224;
      7685: inst = 32'd201344865;
      7686: inst = 32'd203484855;
      7687: inst = 32'd136314880;
      7688: inst = 32'd268468224;
      7689: inst = 32'd201344866;
      7690: inst = 32'd203484855;
      7691: inst = 32'd136314880;
      7692: inst = 32'd268468224;
      7693: inst = 32'd201344867;
      7694: inst = 32'd203484855;
      7695: inst = 32'd136314880;
      7696: inst = 32'd268468224;
      7697: inst = 32'd201344868;
      7698: inst = 32'd203484855;
      7699: inst = 32'd136314880;
      7700: inst = 32'd268468224;
      7701: inst = 32'd201344869;
      7702: inst = 32'd203484855;
      7703: inst = 32'd136314880;
      7704: inst = 32'd268468224;
      7705: inst = 32'd201344870;
      7706: inst = 32'd203484855;
      7707: inst = 32'd136314880;
      7708: inst = 32'd268468224;
      7709: inst = 32'd201344871;
      7710: inst = 32'd203484854;
      7711: inst = 32'd136314880;
      7712: inst = 32'd268468224;
      7713: inst = 32'd201344872;
      7714: inst = 32'd203484854;
      7715: inst = 32'd136314880;
      7716: inst = 32'd268468224;
      7717: inst = 32'd201344873;
      7718: inst = 32'd203484854;
      7719: inst = 32'd136314880;
      7720: inst = 32'd268468224;
      7721: inst = 32'd201344874;
      7722: inst = 32'd203484854;
      7723: inst = 32'd136314880;
      7724: inst = 32'd268468224;
      7725: inst = 32'd201344875;
      7726: inst = 32'd203484854;
      7727: inst = 32'd136314880;
      7728: inst = 32'd268468224;
      7729: inst = 32'd201344876;
      7730: inst = 32'd203484854;
      7731: inst = 32'd136314880;
      7732: inst = 32'd268468224;
      7733: inst = 32'd201344877;
      7734: inst = 32'd203484854;
      7735: inst = 32'd136314880;
      7736: inst = 32'd268468224;
      7737: inst = 32'd201344878;
      7738: inst = 32'd203484854;
      7739: inst = 32'd136314880;
      7740: inst = 32'd268468224;
      7741: inst = 32'd201344879;
      7742: inst = 32'd203484854;
      7743: inst = 32'd136314880;
      7744: inst = 32'd268468224;
      7745: inst = 32'd201344880;
      7746: inst = 32'd203484854;
      7747: inst = 32'd136314880;
      7748: inst = 32'd268468224;
      7749: inst = 32'd201344881;
      7750: inst = 32'd203484854;
      7751: inst = 32'd136314880;
      7752: inst = 32'd268468224;
      7753: inst = 32'd201344882;
      7754: inst = 32'd203484854;
      7755: inst = 32'd136314880;
      7756: inst = 32'd268468224;
      7757: inst = 32'd201344883;
      7758: inst = 32'd203484854;
      7759: inst = 32'd136314880;
      7760: inst = 32'd268468224;
      7761: inst = 32'd201344884;
      7762: inst = 32'd203484854;
      7763: inst = 32'd136314880;
      7764: inst = 32'd268468224;
      7765: inst = 32'd201344885;
      7766: inst = 32'd203484854;
      7767: inst = 32'd136314880;
      7768: inst = 32'd268468224;
      7769: inst = 32'd201344886;
      7770: inst = 32'd203484854;
      7771: inst = 32'd136314880;
      7772: inst = 32'd268468224;
      7773: inst = 32'd201344887;
      7774: inst = 32'd203484854;
      7775: inst = 32'd136314880;
      7776: inst = 32'd268468224;
      7777: inst = 32'd201344888;
      7778: inst = 32'd203484854;
      7779: inst = 32'd136314880;
      7780: inst = 32'd268468224;
      7781: inst = 32'd201344889;
      7782: inst = 32'd203484854;
      7783: inst = 32'd136314880;
      7784: inst = 32'd268468224;
      7785: inst = 32'd201344890;
      7786: inst = 32'd203484855;
      7787: inst = 32'd136314880;
      7788: inst = 32'd268468224;
      7789: inst = 32'd201344891;
      7790: inst = 32'd203482808;
      7791: inst = 32'd136314880;
      7792: inst = 32'd268468224;
      7793: inst = 32'd201344892;
      7794: inst = 32'd203489278;
      7795: inst = 32'd136314880;
      7796: inst = 32'd268468224;
      7797: inst = 32'd201344893;
      7798: inst = 32'd203489279;
      7799: inst = 32'd136314880;
      7800: inst = 32'd268468224;
      7801: inst = 32'd201344894;
      7802: inst = 32'd203489279;
      7803: inst = 32'd136314880;
      7804: inst = 32'd268468224;
      7805: inst = 32'd201344895;
      7806: inst = 32'd203489279;
      7807: inst = 32'd136314880;
      7808: inst = 32'd268468224;
      7809: inst = 32'd201344896;
      7810: inst = 32'd203489279;
      7811: inst = 32'd136314880;
      7812: inst = 32'd268468224;
      7813: inst = 32'd201344897;
      7814: inst = 32'd203489279;
      7815: inst = 32'd136314880;
      7816: inst = 32'd268468224;
      7817: inst = 32'd201344898;
      7818: inst = 32'd203489279;
      7819: inst = 32'd136314880;
      7820: inst = 32'd268468224;
      7821: inst = 32'd201344899;
      7822: inst = 32'd203489279;
      7823: inst = 32'd136314880;
      7824: inst = 32'd268468224;
      7825: inst = 32'd201344900;
      7826: inst = 32'd203489279;
      7827: inst = 32'd136314880;
      7828: inst = 32'd268468224;
      7829: inst = 32'd201344901;
      7830: inst = 32'd203489279;
      7831: inst = 32'd136314880;
      7832: inst = 32'd268468224;
      7833: inst = 32'd201344902;
      7834: inst = 32'd203489279;
      7835: inst = 32'd136314880;
      7836: inst = 32'd268468224;
      7837: inst = 32'd201344903;
      7838: inst = 32'd203489279;
      7839: inst = 32'd136314880;
      7840: inst = 32'd268468224;
      7841: inst = 32'd201344904;
      7842: inst = 32'd203489279;
      7843: inst = 32'd136314880;
      7844: inst = 32'd268468224;
      7845: inst = 32'd201344905;
      7846: inst = 32'd203489279;
      7847: inst = 32'd136314880;
      7848: inst = 32'd268468224;
      7849: inst = 32'd201344906;
      7850: inst = 32'd203489279;
      7851: inst = 32'd136314880;
      7852: inst = 32'd268468224;
      7853: inst = 32'd201344907;
      7854: inst = 32'd203489279;
      7855: inst = 32'd136314880;
      7856: inst = 32'd268468224;
      7857: inst = 32'd201344908;
      7858: inst = 32'd203489279;
      7859: inst = 32'd136314880;
      7860: inst = 32'd268468224;
      7861: inst = 32'd201344909;
      7862: inst = 32'd203489279;
      7863: inst = 32'd136314880;
      7864: inst = 32'd268468224;
      7865: inst = 32'd201344910;
      7866: inst = 32'd203489279;
      7867: inst = 32'd136314880;
      7868: inst = 32'd268468224;
      7869: inst = 32'd201344911;
      7870: inst = 32'd203489279;
      7871: inst = 32'd136314880;
      7872: inst = 32'd268468224;
      7873: inst = 32'd201344912;
      7874: inst = 32'd203489279;
      7875: inst = 32'd136314880;
      7876: inst = 32'd268468224;
      7877: inst = 32'd201344913;
      7878: inst = 32'd203489279;
      7879: inst = 32'd136314880;
      7880: inst = 32'd268468224;
      7881: inst = 32'd201344914;
      7882: inst = 32'd203489279;
      7883: inst = 32'd136314880;
      7884: inst = 32'd268468224;
      7885: inst = 32'd201344915;
      7886: inst = 32'd203489279;
      7887: inst = 32'd136314880;
      7888: inst = 32'd268468224;
      7889: inst = 32'd201344916;
      7890: inst = 32'd203489279;
      7891: inst = 32'd136314880;
      7892: inst = 32'd268468224;
      7893: inst = 32'd201344917;
      7894: inst = 32'd203489279;
      7895: inst = 32'd136314880;
      7896: inst = 32'd268468224;
      7897: inst = 32'd201344918;
      7898: inst = 32'd203489279;
      7899: inst = 32'd136314880;
      7900: inst = 32'd268468224;
      7901: inst = 32'd201344919;
      7902: inst = 32'd203489279;
      7903: inst = 32'd136314880;
      7904: inst = 32'd268468224;
      7905: inst = 32'd201344920;
      7906: inst = 32'd203489279;
      7907: inst = 32'd136314880;
      7908: inst = 32'd268468224;
      7909: inst = 32'd201344921;
      7910: inst = 32'd203489279;
      7911: inst = 32'd136314880;
      7912: inst = 32'd268468224;
      7913: inst = 32'd201344922;
      7914: inst = 32'd203489279;
      7915: inst = 32'd136314880;
      7916: inst = 32'd268468224;
      7917: inst = 32'd201344923;
      7918: inst = 32'd203489279;
      7919: inst = 32'd136314880;
      7920: inst = 32'd268468224;
      7921: inst = 32'd201344924;
      7922: inst = 32'd203489279;
      7923: inst = 32'd136314880;
      7924: inst = 32'd268468224;
      7925: inst = 32'd201344925;
      7926: inst = 32'd203489279;
      7927: inst = 32'd136314880;
      7928: inst = 32'd268468224;
      7929: inst = 32'd201344926;
      7930: inst = 32'd203489279;
      7931: inst = 32'd136314880;
      7932: inst = 32'd268468224;
      7933: inst = 32'd201344927;
      7934: inst = 32'd203489279;
      7935: inst = 32'd136314880;
      7936: inst = 32'd268468224;
      7937: inst = 32'd201344928;
      7938: inst = 32'd203489279;
      7939: inst = 32'd136314880;
      7940: inst = 32'd268468224;
      7941: inst = 32'd201344929;
      7942: inst = 32'd203489279;
      7943: inst = 32'd136314880;
      7944: inst = 32'd268468224;
      7945: inst = 32'd201344930;
      7946: inst = 32'd203489247;
      7947: inst = 32'd136314880;
      7948: inst = 32'd268468224;
      7949: inst = 32'd201344931;
      7950: inst = 32'd203489279;
      7951: inst = 32'd136314880;
      7952: inst = 32'd268468224;
      7953: inst = 32'd201344932;
      7954: inst = 32'd203482840;
      7955: inst = 32'd136314880;
      7956: inst = 32'd268468224;
      7957: inst = 32'd201344933;
      7958: inst = 32'd203484886;
      7959: inst = 32'd136314880;
      7960: inst = 32'd268468224;
      7961: inst = 32'd201344934;
      7962: inst = 32'd203486869;
      7963: inst = 32'd136314880;
      7964: inst = 32'd268468224;
      7965: inst = 32'd201344935;
      7966: inst = 32'd203484854;
      7967: inst = 32'd136314880;
      7968: inst = 32'd268468224;
      7969: inst = 32'd201344936;
      7970: inst = 32'd203484854;
      7971: inst = 32'd136314880;
      7972: inst = 32'd268468224;
      7973: inst = 32'd201344937;
      7974: inst = 32'd203486934;
      7975: inst = 32'd136314880;
      7976: inst = 32'd268468224;
      7977: inst = 32'd201344938;
      7978: inst = 32'd203486870;
      7979: inst = 32'd136314880;
      7980: inst = 32'd268468224;
      7981: inst = 32'd201344939;
      7982: inst = 32'd203486903;
      7983: inst = 32'd136314880;
      7984: inst = 32'd268468224;
      7985: inst = 32'd201344940;
      7986: inst = 32'd203480759;
      7987: inst = 32'd136314880;
      7988: inst = 32'd268468224;
      7989: inst = 32'd201344941;
      7990: inst = 32'd203482838;
      7991: inst = 32'd136314880;
      7992: inst = 32'd268468224;
      7993: inst = 32'd201344942;
      7994: inst = 32'd203488949;
      7995: inst = 32'd136314880;
      7996: inst = 32'd268468224;
      7997: inst = 32'd201344943;
      7998: inst = 32'd203469638;
      7999: inst = 32'd136314880;
      8000: inst = 32'd268468224;
      8001: inst = 32'd201344944;
      8002: inst = 32'd203477959;
      8003: inst = 32'd136314880;
      8004: inst = 32'd268468224;
      8005: inst = 32'd201344945;
      8006: inst = 32'd203480006;
      8007: inst = 32'd136314880;
      8008: inst = 32'd268468224;
      8009: inst = 32'd201344946;
      8010: inst = 32'd203480004;
      8011: inst = 32'd136314880;
      8012: inst = 32'd268468224;
      8013: inst = 32'd201344947;
      8014: inst = 32'd203480003;
      8015: inst = 32'd136314880;
      8016: inst = 32'd268468224;
      8017: inst = 32'd201344948;
      8018: inst = 32'd203480003;
      8019: inst = 32'd136314880;
      8020: inst = 32'd268468224;
      8021: inst = 32'd201344949;
      8022: inst = 32'd203480003;
      8023: inst = 32'd136314880;
      8024: inst = 32'd268468224;
      8025: inst = 32'd201344950;
      8026: inst = 32'd203480004;
      8027: inst = 32'd136314880;
      8028: inst = 32'd268468224;
      8029: inst = 32'd201344951;
      8030: inst = 32'd203481990;
      8031: inst = 32'd136314880;
      8032: inst = 32'd268468224;
      8033: inst = 32'd201344952;
      8034: inst = 32'd203484039;
      8035: inst = 32'd136314880;
      8036: inst = 32'd268468224;
      8037: inst = 32'd201344953;
      8038: inst = 32'd203482023;
      8039: inst = 32'd136314880;
      8040: inst = 32'd268468224;
      8041: inst = 32'd201344954;
      8042: inst = 32'd203479974;
      8043: inst = 32'd136314880;
      8044: inst = 32'd268468224;
      8045: inst = 32'd201344955;
      8046: inst = 32'd203477989;
      8047: inst = 32'd136314880;
      8048: inst = 32'd268468224;
      8049: inst = 32'd201344956;
      8050: inst = 32'd203475973;
      8051: inst = 32'd136314880;
      8052: inst = 32'd268468224;
      8053: inst = 32'd201344957;
      8054: inst = 32'd203477957;
      8055: inst = 32'd136314880;
      8056: inst = 32'd268468224;
      8057: inst = 32'd201344958;
      8058: inst = 32'd203481957;
      8059: inst = 32'd136314880;
      8060: inst = 32'd268468224;
      8061: inst = 32'd201344959;
      8062: inst = 32'd203479682;
      8063: inst = 32'd136314880;
      8064: inst = 32'd268468224;
      8065: inst = 32'd201344960;
      8066: inst = 32'd203484855;
      8067: inst = 32'd136314880;
      8068: inst = 32'd268468224;
      8069: inst = 32'd201344961;
      8070: inst = 32'd203484855;
      8071: inst = 32'd136314880;
      8072: inst = 32'd268468224;
      8073: inst = 32'd201344962;
      8074: inst = 32'd203484855;
      8075: inst = 32'd136314880;
      8076: inst = 32'd268468224;
      8077: inst = 32'd201344963;
      8078: inst = 32'd203484855;
      8079: inst = 32'd136314880;
      8080: inst = 32'd268468224;
      8081: inst = 32'd201344964;
      8082: inst = 32'd203484855;
      8083: inst = 32'd136314880;
      8084: inst = 32'd268468224;
      8085: inst = 32'd201344965;
      8086: inst = 32'd203484854;
      8087: inst = 32'd136314880;
      8088: inst = 32'd268468224;
      8089: inst = 32'd201344966;
      8090: inst = 32'd203484854;
      8091: inst = 32'd136314880;
      8092: inst = 32'd268468224;
      8093: inst = 32'd201344967;
      8094: inst = 32'd203484854;
      8095: inst = 32'd136314880;
      8096: inst = 32'd268468224;
      8097: inst = 32'd201344968;
      8098: inst = 32'd203484854;
      8099: inst = 32'd136314880;
      8100: inst = 32'd268468224;
      8101: inst = 32'd201344969;
      8102: inst = 32'd203484854;
      8103: inst = 32'd136314880;
      8104: inst = 32'd268468224;
      8105: inst = 32'd201344970;
      8106: inst = 32'd203484854;
      8107: inst = 32'd136314880;
      8108: inst = 32'd268468224;
      8109: inst = 32'd201344971;
      8110: inst = 32'd203484854;
      8111: inst = 32'd136314880;
      8112: inst = 32'd268468224;
      8113: inst = 32'd201344972;
      8114: inst = 32'd203484854;
      8115: inst = 32'd136314880;
      8116: inst = 32'd268468224;
      8117: inst = 32'd201344973;
      8118: inst = 32'd203484854;
      8119: inst = 32'd136314880;
      8120: inst = 32'd268468224;
      8121: inst = 32'd201344974;
      8122: inst = 32'd203484854;
      8123: inst = 32'd136314880;
      8124: inst = 32'd268468224;
      8125: inst = 32'd201344975;
      8126: inst = 32'd203484854;
      8127: inst = 32'd136314880;
      8128: inst = 32'd268468224;
      8129: inst = 32'd201344976;
      8130: inst = 32'd203484854;
      8131: inst = 32'd136314880;
      8132: inst = 32'd268468224;
      8133: inst = 32'd201344977;
      8134: inst = 32'd203484854;
      8135: inst = 32'd136314880;
      8136: inst = 32'd268468224;
      8137: inst = 32'd201344978;
      8138: inst = 32'd203484854;
      8139: inst = 32'd136314880;
      8140: inst = 32'd268468224;
      8141: inst = 32'd201344979;
      8142: inst = 32'd203484854;
      8143: inst = 32'd136314880;
      8144: inst = 32'd268468224;
      8145: inst = 32'd201344980;
      8146: inst = 32'd203484854;
      8147: inst = 32'd136314880;
      8148: inst = 32'd268468224;
      8149: inst = 32'd201344981;
      8150: inst = 32'd203484854;
      8151: inst = 32'd136314880;
      8152: inst = 32'd268468224;
      8153: inst = 32'd201344982;
      8154: inst = 32'd203484854;
      8155: inst = 32'd136314880;
      8156: inst = 32'd268468224;
      8157: inst = 32'd201344983;
      8158: inst = 32'd203484854;
      8159: inst = 32'd136314880;
      8160: inst = 32'd268468224;
      8161: inst = 32'd201344984;
      8162: inst = 32'd203484854;
      8163: inst = 32'd136314880;
      8164: inst = 32'd268468224;
      8165: inst = 32'd201344985;
      8166: inst = 32'd203484854;
      8167: inst = 32'd136314880;
      8168: inst = 32'd268468224;
      8169: inst = 32'd201344986;
      8170: inst = 32'd203484855;
      8171: inst = 32'd136314880;
      8172: inst = 32'd268468224;
      8173: inst = 32'd201344987;
      8174: inst = 32'd203482808;
      8175: inst = 32'd136314880;
      8176: inst = 32'd268468224;
      8177: inst = 32'd201344988;
      8178: inst = 32'd203489278;
      8179: inst = 32'd136314880;
      8180: inst = 32'd268468224;
      8181: inst = 32'd201344989;
      8182: inst = 32'd203489279;
      8183: inst = 32'd136314880;
      8184: inst = 32'd268468224;
      8185: inst = 32'd201344990;
      8186: inst = 32'd203489279;
      8187: inst = 32'd136314880;
      8188: inst = 32'd268468224;
      8189: inst = 32'd201344991;
      8190: inst = 32'd203489279;
      8191: inst = 32'd136314880;
      8192: inst = 32'd268468224;
      8193: inst = 32'd201344992;
      8194: inst = 32'd203489279;
      8195: inst = 32'd136314880;
      8196: inst = 32'd268468224;
      8197: inst = 32'd201344993;
      8198: inst = 32'd203489279;
      8199: inst = 32'd136314880;
      8200: inst = 32'd268468224;
      8201: inst = 32'd201344994;
      8202: inst = 32'd203489279;
      8203: inst = 32'd136314880;
      8204: inst = 32'd268468224;
      8205: inst = 32'd201344995;
      8206: inst = 32'd203489279;
      8207: inst = 32'd136314880;
      8208: inst = 32'd268468224;
      8209: inst = 32'd201344996;
      8210: inst = 32'd203489279;
      8211: inst = 32'd136314880;
      8212: inst = 32'd268468224;
      8213: inst = 32'd201344997;
      8214: inst = 32'd203489279;
      8215: inst = 32'd136314880;
      8216: inst = 32'd268468224;
      8217: inst = 32'd201344998;
      8218: inst = 32'd203489279;
      8219: inst = 32'd136314880;
      8220: inst = 32'd268468224;
      8221: inst = 32'd201344999;
      8222: inst = 32'd203489279;
      8223: inst = 32'd136314880;
      8224: inst = 32'd268468224;
      8225: inst = 32'd201345000;
      8226: inst = 32'd203489279;
      8227: inst = 32'd136314880;
      8228: inst = 32'd268468224;
      8229: inst = 32'd201345001;
      8230: inst = 32'd203489279;
      8231: inst = 32'd136314880;
      8232: inst = 32'd268468224;
      8233: inst = 32'd201345002;
      8234: inst = 32'd203489279;
      8235: inst = 32'd136314880;
      8236: inst = 32'd268468224;
      8237: inst = 32'd201345003;
      8238: inst = 32'd203489279;
      8239: inst = 32'd136314880;
      8240: inst = 32'd268468224;
      8241: inst = 32'd201345004;
      8242: inst = 32'd203489279;
      8243: inst = 32'd136314880;
      8244: inst = 32'd268468224;
      8245: inst = 32'd201345005;
      8246: inst = 32'd203489279;
      8247: inst = 32'd136314880;
      8248: inst = 32'd268468224;
      8249: inst = 32'd201345006;
      8250: inst = 32'd203489279;
      8251: inst = 32'd136314880;
      8252: inst = 32'd268468224;
      8253: inst = 32'd201345007;
      8254: inst = 32'd203489279;
      8255: inst = 32'd136314880;
      8256: inst = 32'd268468224;
      8257: inst = 32'd201345008;
      8258: inst = 32'd203489279;
      8259: inst = 32'd136314880;
      8260: inst = 32'd268468224;
      8261: inst = 32'd201345009;
      8262: inst = 32'd203489279;
      8263: inst = 32'd136314880;
      8264: inst = 32'd268468224;
      8265: inst = 32'd201345010;
      8266: inst = 32'd203489279;
      8267: inst = 32'd136314880;
      8268: inst = 32'd268468224;
      8269: inst = 32'd201345011;
      8270: inst = 32'd203489279;
      8271: inst = 32'd136314880;
      8272: inst = 32'd268468224;
      8273: inst = 32'd201345012;
      8274: inst = 32'd203489279;
      8275: inst = 32'd136314880;
      8276: inst = 32'd268468224;
      8277: inst = 32'd201345013;
      8278: inst = 32'd203489279;
      8279: inst = 32'd136314880;
      8280: inst = 32'd268468224;
      8281: inst = 32'd201345014;
      8282: inst = 32'd203489279;
      8283: inst = 32'd136314880;
      8284: inst = 32'd268468224;
      8285: inst = 32'd201345015;
      8286: inst = 32'd203489279;
      8287: inst = 32'd136314880;
      8288: inst = 32'd268468224;
      8289: inst = 32'd201345016;
      8290: inst = 32'd203489279;
      8291: inst = 32'd136314880;
      8292: inst = 32'd268468224;
      8293: inst = 32'd201345017;
      8294: inst = 32'd203489279;
      8295: inst = 32'd136314880;
      8296: inst = 32'd268468224;
      8297: inst = 32'd201345018;
      8298: inst = 32'd203489279;
      8299: inst = 32'd136314880;
      8300: inst = 32'd268468224;
      8301: inst = 32'd201345019;
      8302: inst = 32'd203489279;
      8303: inst = 32'd136314880;
      8304: inst = 32'd268468224;
      8305: inst = 32'd201345020;
      8306: inst = 32'd203489279;
      8307: inst = 32'd136314880;
      8308: inst = 32'd268468224;
      8309: inst = 32'd201345021;
      8310: inst = 32'd203489279;
      8311: inst = 32'd136314880;
      8312: inst = 32'd268468224;
      8313: inst = 32'd201345022;
      8314: inst = 32'd203489279;
      8315: inst = 32'd136314880;
      8316: inst = 32'd268468224;
      8317: inst = 32'd201345023;
      8318: inst = 32'd203489279;
      8319: inst = 32'd136314880;
      8320: inst = 32'd268468224;
      8321: inst = 32'd201345024;
      8322: inst = 32'd203489279;
      8323: inst = 32'd136314880;
      8324: inst = 32'd268468224;
      8325: inst = 32'd201345025;
      8326: inst = 32'd203489279;
      8327: inst = 32'd136314880;
      8328: inst = 32'd268468224;
      8329: inst = 32'd201345026;
      8330: inst = 32'd203489247;
      8331: inst = 32'd136314880;
      8332: inst = 32'd268468224;
      8333: inst = 32'd201345027;
      8334: inst = 32'd203489279;
      8335: inst = 32'd136314880;
      8336: inst = 32'd268468224;
      8337: inst = 32'd201345028;
      8338: inst = 32'd203482840;
      8339: inst = 32'd136314880;
      8340: inst = 32'd268468224;
      8341: inst = 32'd201345029;
      8342: inst = 32'd203484886;
      8343: inst = 32'd136314880;
      8344: inst = 32'd268468224;
      8345: inst = 32'd201345030;
      8346: inst = 32'd203486869;
      8347: inst = 32'd136314880;
      8348: inst = 32'd268468224;
      8349: inst = 32'd201345031;
      8350: inst = 32'd203484854;
      8351: inst = 32'd136314880;
      8352: inst = 32'd268468224;
      8353: inst = 32'd201345032;
      8354: inst = 32'd203484854;
      8355: inst = 32'd136314880;
      8356: inst = 32'd268468224;
      8357: inst = 32'd201345033;
      8358: inst = 32'd203484854;
      8359: inst = 32'd136314880;
      8360: inst = 32'd268468224;
      8361: inst = 32'd201345034;
      8362: inst = 32'd203486902;
      8363: inst = 32'd136314880;
      8364: inst = 32'd268468224;
      8365: inst = 32'd201345035;
      8366: inst = 32'd203486936;
      8367: inst = 32'd136314880;
      8368: inst = 32'd268468224;
      8369: inst = 32'd201345036;
      8370: inst = 32'd203482839;
      8371: inst = 32'd136314880;
      8372: inst = 32'd268468224;
      8373: inst = 32'd201345037;
      8374: inst = 32'd203482806;
      8375: inst = 32'd136314880;
      8376: inst = 32'd268468224;
      8377: inst = 32'd201345038;
      8378: inst = 32'd203488884;
      8379: inst = 32'd136314880;
      8380: inst = 32'd268468224;
      8381: inst = 32'd201345039;
      8382: inst = 32'd203467460;
      8383: inst = 32'd136314880;
      8384: inst = 32'd268468224;
      8385: inst = 32'd201345040;
      8386: inst = 32'd203480007;
      8387: inst = 32'd136314880;
      8388: inst = 32'd268468224;
      8389: inst = 32'd201345041;
      8390: inst = 32'd203482054;
      8391: inst = 32'd136314880;
      8392: inst = 32'd268468224;
      8393: inst = 32'd201345042;
      8394: inst = 32'd203484069;
      8395: inst = 32'd136314880;
      8396: inst = 32'd268468224;
      8397: inst = 32'd201345043;
      8398: inst = 32'd203484068;
      8399: inst = 32'd136314880;
      8400: inst = 32'd268468224;
      8401: inst = 32'd201345044;
      8402: inst = 32'd203484100;
      8403: inst = 32'd136314880;
      8404: inst = 32'd268468224;
      8405: inst = 32'd201345045;
      8406: inst = 32'd203482052;
      8407: inst = 32'd136314880;
      8408: inst = 32'd268468224;
      8409: inst = 32'd201345046;
      8410: inst = 32'd203482053;
      8411: inst = 32'd136314880;
      8412: inst = 32'd268468224;
      8413: inst = 32'd201345047;
      8414: inst = 32'd203482054;
      8415: inst = 32'd136314880;
      8416: inst = 32'd268468224;
      8417: inst = 32'd201345048;
      8418: inst = 32'd203482023;
      8419: inst = 32'd136314880;
      8420: inst = 32'd268468224;
      8421: inst = 32'd201345049;
      8422: inst = 32'd203482023;
      8423: inst = 32'd136314880;
      8424: inst = 32'd268468224;
      8425: inst = 32'd201345050;
      8426: inst = 32'd203480006;
      8427: inst = 32'd136314880;
      8428: inst = 32'd268468224;
      8429: inst = 32'd201345051;
      8430: inst = 32'd203480037;
      8431: inst = 32'd136314880;
      8432: inst = 32'd268468224;
      8433: inst = 32'd201345052;
      8434: inst = 32'd203477988;
      8435: inst = 32'd136314880;
      8436: inst = 32'd268468224;
      8437: inst = 32'd201345053;
      8438: inst = 32'd203480069;
      8439: inst = 32'd136314880;
      8440: inst = 32'd268468224;
      8441: inst = 32'd201345054;
      8442: inst = 32'd203482021;
      8443: inst = 32'd136314880;
      8444: inst = 32'd268468224;
      8445: inst = 32'd201345055;
      8446: inst = 32'd203477666;
      8447: inst = 32'd136314880;
      8448: inst = 32'd268468224;
      8449: inst = 32'd201345056;
      8450: inst = 32'd203484855;
      8451: inst = 32'd136314880;
      8452: inst = 32'd268468224;
      8453: inst = 32'd201345057;
      8454: inst = 32'd203484855;
      8455: inst = 32'd136314880;
      8456: inst = 32'd268468224;
      8457: inst = 32'd201345058;
      8458: inst = 32'd203484854;
      8459: inst = 32'd136314880;
      8460: inst = 32'd268468224;
      8461: inst = 32'd201345059;
      8462: inst = 32'd203484854;
      8463: inst = 32'd136314880;
      8464: inst = 32'd268468224;
      8465: inst = 32'd201345060;
      8466: inst = 32'd203484854;
      8467: inst = 32'd136314880;
      8468: inst = 32'd268468224;
      8469: inst = 32'd201345061;
      8470: inst = 32'd203484854;
      8471: inst = 32'd136314880;
      8472: inst = 32'd268468224;
      8473: inst = 32'd201345062;
      8474: inst = 32'd203484854;
      8475: inst = 32'd136314880;
      8476: inst = 32'd268468224;
      8477: inst = 32'd201345063;
      8478: inst = 32'd203484854;
      8479: inst = 32'd136314880;
      8480: inst = 32'd268468224;
      8481: inst = 32'd201345064;
      8482: inst = 32'd203484854;
      8483: inst = 32'd136314880;
      8484: inst = 32'd268468224;
      8485: inst = 32'd201345065;
      8486: inst = 32'd203484854;
      8487: inst = 32'd136314880;
      8488: inst = 32'd268468224;
      8489: inst = 32'd201345066;
      8490: inst = 32'd203484854;
      8491: inst = 32'd136314880;
      8492: inst = 32'd268468224;
      8493: inst = 32'd201345067;
      8494: inst = 32'd203484854;
      8495: inst = 32'd136314880;
      8496: inst = 32'd268468224;
      8497: inst = 32'd201345068;
      8498: inst = 32'd203484854;
      8499: inst = 32'd136314880;
      8500: inst = 32'd268468224;
      8501: inst = 32'd201345069;
      8502: inst = 32'd203484854;
      8503: inst = 32'd136314880;
      8504: inst = 32'd268468224;
      8505: inst = 32'd201345070;
      8506: inst = 32'd203484854;
      8507: inst = 32'd136314880;
      8508: inst = 32'd268468224;
      8509: inst = 32'd201345071;
      8510: inst = 32'd203484854;
      8511: inst = 32'd136314880;
      8512: inst = 32'd268468224;
      8513: inst = 32'd201345072;
      8514: inst = 32'd203484854;
      8515: inst = 32'd136314880;
      8516: inst = 32'd268468224;
      8517: inst = 32'd201345073;
      8518: inst = 32'd203484854;
      8519: inst = 32'd136314880;
      8520: inst = 32'd268468224;
      8521: inst = 32'd201345074;
      8522: inst = 32'd203484854;
      8523: inst = 32'd136314880;
      8524: inst = 32'd268468224;
      8525: inst = 32'd201345075;
      8526: inst = 32'd203484854;
      8527: inst = 32'd136314880;
      8528: inst = 32'd268468224;
      8529: inst = 32'd201345076;
      8530: inst = 32'd203484854;
      8531: inst = 32'd136314880;
      8532: inst = 32'd268468224;
      8533: inst = 32'd201345077;
      8534: inst = 32'd203484854;
      8535: inst = 32'd136314880;
      8536: inst = 32'd268468224;
      8537: inst = 32'd201345078;
      8538: inst = 32'd203484854;
      8539: inst = 32'd136314880;
      8540: inst = 32'd268468224;
      8541: inst = 32'd201345079;
      8542: inst = 32'd203484854;
      8543: inst = 32'd136314880;
      8544: inst = 32'd268468224;
      8545: inst = 32'd201345080;
      8546: inst = 32'd203484854;
      8547: inst = 32'd136314880;
      8548: inst = 32'd268468224;
      8549: inst = 32'd201345081;
      8550: inst = 32'd203484854;
      8551: inst = 32'd136314880;
      8552: inst = 32'd268468224;
      8553: inst = 32'd201345082;
      8554: inst = 32'd203484855;
      8555: inst = 32'd136314880;
      8556: inst = 32'd268468224;
      8557: inst = 32'd201345083;
      8558: inst = 32'd203482808;
      8559: inst = 32'd136314880;
      8560: inst = 32'd268468224;
      8561: inst = 32'd201345084;
      8562: inst = 32'd203489278;
      8563: inst = 32'd136314880;
      8564: inst = 32'd268468224;
      8565: inst = 32'd201345085;
      8566: inst = 32'd203489279;
      8567: inst = 32'd136314880;
      8568: inst = 32'd268468224;
      8569: inst = 32'd201345086;
      8570: inst = 32'd203489279;
      8571: inst = 32'd136314880;
      8572: inst = 32'd268468224;
      8573: inst = 32'd201345087;
      8574: inst = 32'd203489279;
      8575: inst = 32'd136314880;
      8576: inst = 32'd268468224;
      8577: inst = 32'd201345088;
      8578: inst = 32'd203489279;
      8579: inst = 32'd136314880;
      8580: inst = 32'd268468224;
      8581: inst = 32'd201345089;
      8582: inst = 32'd203489279;
      8583: inst = 32'd136314880;
      8584: inst = 32'd268468224;
      8585: inst = 32'd201345090;
      8586: inst = 32'd203489279;
      8587: inst = 32'd136314880;
      8588: inst = 32'd268468224;
      8589: inst = 32'd201345091;
      8590: inst = 32'd203489279;
      8591: inst = 32'd136314880;
      8592: inst = 32'd268468224;
      8593: inst = 32'd201345092;
      8594: inst = 32'd203489279;
      8595: inst = 32'd136314880;
      8596: inst = 32'd268468224;
      8597: inst = 32'd201345093;
      8598: inst = 32'd203489279;
      8599: inst = 32'd136314880;
      8600: inst = 32'd268468224;
      8601: inst = 32'd201345094;
      8602: inst = 32'd203489279;
      8603: inst = 32'd136314880;
      8604: inst = 32'd268468224;
      8605: inst = 32'd201345095;
      8606: inst = 32'd203489279;
      8607: inst = 32'd136314880;
      8608: inst = 32'd268468224;
      8609: inst = 32'd201345096;
      8610: inst = 32'd203489279;
      8611: inst = 32'd136314880;
      8612: inst = 32'd268468224;
      8613: inst = 32'd201345097;
      8614: inst = 32'd203489279;
      8615: inst = 32'd136314880;
      8616: inst = 32'd268468224;
      8617: inst = 32'd201345098;
      8618: inst = 32'd203489279;
      8619: inst = 32'd136314880;
      8620: inst = 32'd268468224;
      8621: inst = 32'd201345099;
      8622: inst = 32'd203489279;
      8623: inst = 32'd136314880;
      8624: inst = 32'd268468224;
      8625: inst = 32'd201345100;
      8626: inst = 32'd203489279;
      8627: inst = 32'd136314880;
      8628: inst = 32'd268468224;
      8629: inst = 32'd201345101;
      8630: inst = 32'd203489279;
      8631: inst = 32'd136314880;
      8632: inst = 32'd268468224;
      8633: inst = 32'd201345102;
      8634: inst = 32'd203489279;
      8635: inst = 32'd136314880;
      8636: inst = 32'd268468224;
      8637: inst = 32'd201345103;
      8638: inst = 32'd203489279;
      8639: inst = 32'd136314880;
      8640: inst = 32'd268468224;
      8641: inst = 32'd201345104;
      8642: inst = 32'd203489279;
      8643: inst = 32'd136314880;
      8644: inst = 32'd268468224;
      8645: inst = 32'd201345105;
      8646: inst = 32'd203489279;
      8647: inst = 32'd136314880;
      8648: inst = 32'd268468224;
      8649: inst = 32'd201345106;
      8650: inst = 32'd203489279;
      8651: inst = 32'd136314880;
      8652: inst = 32'd268468224;
      8653: inst = 32'd201345107;
      8654: inst = 32'd203489279;
      8655: inst = 32'd136314880;
      8656: inst = 32'd268468224;
      8657: inst = 32'd201345108;
      8658: inst = 32'd203489279;
      8659: inst = 32'd136314880;
      8660: inst = 32'd268468224;
      8661: inst = 32'd201345109;
      8662: inst = 32'd203489279;
      8663: inst = 32'd136314880;
      8664: inst = 32'd268468224;
      8665: inst = 32'd201345110;
      8666: inst = 32'd203489279;
      8667: inst = 32'd136314880;
      8668: inst = 32'd268468224;
      8669: inst = 32'd201345111;
      8670: inst = 32'd203489279;
      8671: inst = 32'd136314880;
      8672: inst = 32'd268468224;
      8673: inst = 32'd201345112;
      8674: inst = 32'd203489279;
      8675: inst = 32'd136314880;
      8676: inst = 32'd268468224;
      8677: inst = 32'd201345113;
      8678: inst = 32'd203489279;
      8679: inst = 32'd136314880;
      8680: inst = 32'd268468224;
      8681: inst = 32'd201345114;
      8682: inst = 32'd203489279;
      8683: inst = 32'd136314880;
      8684: inst = 32'd268468224;
      8685: inst = 32'd201345115;
      8686: inst = 32'd203489279;
      8687: inst = 32'd136314880;
      8688: inst = 32'd268468224;
      8689: inst = 32'd201345116;
      8690: inst = 32'd203489279;
      8691: inst = 32'd136314880;
      8692: inst = 32'd268468224;
      8693: inst = 32'd201345117;
      8694: inst = 32'd203489279;
      8695: inst = 32'd136314880;
      8696: inst = 32'd268468224;
      8697: inst = 32'd201345118;
      8698: inst = 32'd203489279;
      8699: inst = 32'd136314880;
      8700: inst = 32'd268468224;
      8701: inst = 32'd201345119;
      8702: inst = 32'd203489279;
      8703: inst = 32'd136314880;
      8704: inst = 32'd268468224;
      8705: inst = 32'd201345120;
      8706: inst = 32'd203489279;
      8707: inst = 32'd136314880;
      8708: inst = 32'd268468224;
      8709: inst = 32'd201345121;
      8710: inst = 32'd203489279;
      8711: inst = 32'd136314880;
      8712: inst = 32'd268468224;
      8713: inst = 32'd201345122;
      8714: inst = 32'd203489247;
      8715: inst = 32'd136314880;
      8716: inst = 32'd268468224;
      8717: inst = 32'd201345123;
      8718: inst = 32'd203489279;
      8719: inst = 32'd136314880;
      8720: inst = 32'd268468224;
      8721: inst = 32'd201345124;
      8722: inst = 32'd203482840;
      8723: inst = 32'd136314880;
      8724: inst = 32'd268468224;
      8725: inst = 32'd201345125;
      8726: inst = 32'd203484886;
      8727: inst = 32'd136314880;
      8728: inst = 32'd268468224;
      8729: inst = 32'd201345126;
      8730: inst = 32'd203486869;
      8731: inst = 32'd136314880;
      8732: inst = 32'd268468224;
      8733: inst = 32'd201345127;
      8734: inst = 32'd203484854;
      8735: inst = 32'd136314880;
      8736: inst = 32'd268468224;
      8737: inst = 32'd201345128;
      8738: inst = 32'd203484887;
      8739: inst = 32'd136314880;
      8740: inst = 32'd268468224;
      8741: inst = 32'd201345129;
      8742: inst = 32'd203484822;
      8743: inst = 32'd136314880;
      8744: inst = 32'd268468224;
      8745: inst = 32'd201345130;
      8746: inst = 32'd203486870;
      8747: inst = 32'd136314880;
      8748: inst = 32'd268468224;
      8749: inst = 32'd201345131;
      8750: inst = 32'd203484822;
      8751: inst = 32'd136314880;
      8752: inst = 32'd268468224;
      8753: inst = 32'd201345132;
      8754: inst = 32'd203482839;
      8755: inst = 32'd136314880;
      8756: inst = 32'd268468224;
      8757: inst = 32'd201345133;
      8758: inst = 32'd203484919;
      8759: inst = 32'd136314880;
      8760: inst = 32'd268468224;
      8761: inst = 32'd201345134;
      8762: inst = 32'd203488949;
      8763: inst = 32'd136314880;
      8764: inst = 32'd268468224;
      8765: inst = 32'd201345135;
      8766: inst = 32'd203469573;
      8767: inst = 32'd136314880;
      8768: inst = 32'd268468224;
      8769: inst = 32'd201345136;
      8770: inst = 32'd203482022;
      8771: inst = 32'd136314880;
      8772: inst = 32'd268468224;
      8773: inst = 32'd201345137;
      8774: inst = 32'd203481990;
      8775: inst = 32'd136314880;
      8776: inst = 32'd268468224;
      8777: inst = 32'd201345138;
      8778: inst = 32'd203484006;
      8779: inst = 32'd136314880;
      8780: inst = 32'd268468224;
      8781: inst = 32'd201345139;
      8782: inst = 32'd203484005;
      8783: inst = 32'd136314880;
      8784: inst = 32'd268468224;
      8785: inst = 32'd201345140;
      8786: inst = 32'd203484037;
      8787: inst = 32'd136314880;
      8788: inst = 32'd268468224;
      8789: inst = 32'd201345141;
      8790: inst = 32'd203482020;
      8791: inst = 32'd136314880;
      8792: inst = 32'd268468224;
      8793: inst = 32'd201345142;
      8794: inst = 32'd203479973;
      8795: inst = 32'd136314880;
      8796: inst = 32'd268468224;
      8797: inst = 32'd201345143;
      8798: inst = 32'd203480005;
      8799: inst = 32'd136314880;
      8800: inst = 32'd268468224;
      8801: inst = 32'd201345144;
      8802: inst = 32'd203479974;
      8803: inst = 32'd136314880;
      8804: inst = 32'd268468224;
      8805: inst = 32'd201345145;
      8806: inst = 32'd203479974;
      8807: inst = 32'd136314880;
      8808: inst = 32'd268468224;
      8809: inst = 32'd201345146;
      8810: inst = 32'd203479973;
      8811: inst = 32'd136314880;
      8812: inst = 32'd268468224;
      8813: inst = 32'd201345147;
      8814: inst = 32'd203480004;
      8815: inst = 32'd136314880;
      8816: inst = 32'd268468224;
      8817: inst = 32'd201345148;
      8818: inst = 32'd203480003;
      8819: inst = 32'd136314880;
      8820: inst = 32'd268468224;
      8821: inst = 32'd201345149;
      8822: inst = 32'd203480036;
      8823: inst = 32'd136314880;
      8824: inst = 32'd268468224;
      8825: inst = 32'd201345150;
      8826: inst = 32'd203480037;
      8827: inst = 32'd136314880;
      8828: inst = 32'd268468224;
      8829: inst = 32'd201345151;
      8830: inst = 32'd203471586;
      8831: inst = 32'd136314880;
      8832: inst = 32'd268468224;
      8833: inst = 32'd201345152;
      8834: inst = 32'd203484854;
      8835: inst = 32'd136314880;
      8836: inst = 32'd268468224;
      8837: inst = 32'd201345153;
      8838: inst = 32'd203484854;
      8839: inst = 32'd136314880;
      8840: inst = 32'd268468224;
      8841: inst = 32'd201345154;
      8842: inst = 32'd203484854;
      8843: inst = 32'd136314880;
      8844: inst = 32'd268468224;
      8845: inst = 32'd201345155;
      8846: inst = 32'd203484854;
      8847: inst = 32'd136314880;
      8848: inst = 32'd268468224;
      8849: inst = 32'd201345156;
      8850: inst = 32'd203484854;
      8851: inst = 32'd136314880;
      8852: inst = 32'd268468224;
      8853: inst = 32'd201345157;
      8854: inst = 32'd203484854;
      8855: inst = 32'd136314880;
      8856: inst = 32'd268468224;
      8857: inst = 32'd201345158;
      8858: inst = 32'd203484854;
      8859: inst = 32'd136314880;
      8860: inst = 32'd268468224;
      8861: inst = 32'd201345159;
      8862: inst = 32'd203484854;
      8863: inst = 32'd136314880;
      8864: inst = 32'd268468224;
      8865: inst = 32'd201345160;
      8866: inst = 32'd203484854;
      8867: inst = 32'd136314880;
      8868: inst = 32'd268468224;
      8869: inst = 32'd201345161;
      8870: inst = 32'd203484855;
      8871: inst = 32'd136314880;
      8872: inst = 32'd268468224;
      8873: inst = 32'd201345162;
      8874: inst = 32'd203484855;
      8875: inst = 32'd136314880;
      8876: inst = 32'd268468224;
      8877: inst = 32'd201345163;
      8878: inst = 32'd203484854;
      8879: inst = 32'd136314880;
      8880: inst = 32'd268468224;
      8881: inst = 32'd201345164;
      8882: inst = 32'd203484854;
      8883: inst = 32'd136314880;
      8884: inst = 32'd268468224;
      8885: inst = 32'd201345165;
      8886: inst = 32'd203484854;
      8887: inst = 32'd136314880;
      8888: inst = 32'd268468224;
      8889: inst = 32'd201345166;
      8890: inst = 32'd203484854;
      8891: inst = 32'd136314880;
      8892: inst = 32'd268468224;
      8893: inst = 32'd201345167;
      8894: inst = 32'd203484854;
      8895: inst = 32'd136314880;
      8896: inst = 32'd268468224;
      8897: inst = 32'd201345168;
      8898: inst = 32'd203484854;
      8899: inst = 32'd136314880;
      8900: inst = 32'd268468224;
      8901: inst = 32'd201345169;
      8902: inst = 32'd203484854;
      8903: inst = 32'd136314880;
      8904: inst = 32'd268468224;
      8905: inst = 32'd201345170;
      8906: inst = 32'd203484854;
      8907: inst = 32'd136314880;
      8908: inst = 32'd268468224;
      8909: inst = 32'd201345171;
      8910: inst = 32'd203484854;
      8911: inst = 32'd136314880;
      8912: inst = 32'd268468224;
      8913: inst = 32'd201345172;
      8914: inst = 32'd203484854;
      8915: inst = 32'd136314880;
      8916: inst = 32'd268468224;
      8917: inst = 32'd201345173;
      8918: inst = 32'd203484854;
      8919: inst = 32'd136314880;
      8920: inst = 32'd268468224;
      8921: inst = 32'd201345174;
      8922: inst = 32'd203484854;
      8923: inst = 32'd136314880;
      8924: inst = 32'd268468224;
      8925: inst = 32'd201345175;
      8926: inst = 32'd203484854;
      8927: inst = 32'd136314880;
      8928: inst = 32'd268468224;
      8929: inst = 32'd201345176;
      8930: inst = 32'd203484854;
      8931: inst = 32'd136314880;
      8932: inst = 32'd268468224;
      8933: inst = 32'd201345177;
      8934: inst = 32'd203484854;
      8935: inst = 32'd136314880;
      8936: inst = 32'd268468224;
      8937: inst = 32'd201345178;
      8938: inst = 32'd203484855;
      8939: inst = 32'd136314880;
      8940: inst = 32'd268468224;
      8941: inst = 32'd201345179;
      8942: inst = 32'd203482808;
      8943: inst = 32'd136314880;
      8944: inst = 32'd268468224;
      8945: inst = 32'd201345180;
      8946: inst = 32'd203489278;
      8947: inst = 32'd136314880;
      8948: inst = 32'd268468224;
      8949: inst = 32'd201345181;
      8950: inst = 32'd203489279;
      8951: inst = 32'd136314880;
      8952: inst = 32'd268468224;
      8953: inst = 32'd201345182;
      8954: inst = 32'd203489279;
      8955: inst = 32'd136314880;
      8956: inst = 32'd268468224;
      8957: inst = 32'd201345183;
      8958: inst = 32'd203489279;
      8959: inst = 32'd136314880;
      8960: inst = 32'd268468224;
      8961: inst = 32'd201345184;
      8962: inst = 32'd203489279;
      8963: inst = 32'd136314880;
      8964: inst = 32'd268468224;
      8965: inst = 32'd201345185;
      8966: inst = 32'd203489279;
      8967: inst = 32'd136314880;
      8968: inst = 32'd268468224;
      8969: inst = 32'd201345186;
      8970: inst = 32'd203489279;
      8971: inst = 32'd136314880;
      8972: inst = 32'd268468224;
      8973: inst = 32'd201345187;
      8974: inst = 32'd203489279;
      8975: inst = 32'd136314880;
      8976: inst = 32'd268468224;
      8977: inst = 32'd201345188;
      8978: inst = 32'd203489279;
      8979: inst = 32'd136314880;
      8980: inst = 32'd268468224;
      8981: inst = 32'd201345189;
      8982: inst = 32'd203489279;
      8983: inst = 32'd136314880;
      8984: inst = 32'd268468224;
      8985: inst = 32'd201345190;
      8986: inst = 32'd203489279;
      8987: inst = 32'd136314880;
      8988: inst = 32'd268468224;
      8989: inst = 32'd201345191;
      8990: inst = 32'd203489279;
      8991: inst = 32'd136314880;
      8992: inst = 32'd268468224;
      8993: inst = 32'd201345192;
      8994: inst = 32'd203489279;
      8995: inst = 32'd136314880;
      8996: inst = 32'd268468224;
      8997: inst = 32'd201345193;
      8998: inst = 32'd203489279;
      8999: inst = 32'd136314880;
      9000: inst = 32'd268468224;
      9001: inst = 32'd201345194;
      9002: inst = 32'd203489279;
      9003: inst = 32'd136314880;
      9004: inst = 32'd268468224;
      9005: inst = 32'd201345195;
      9006: inst = 32'd203489279;
      9007: inst = 32'd136314880;
      9008: inst = 32'd268468224;
      9009: inst = 32'd201345196;
      9010: inst = 32'd203489279;
      9011: inst = 32'd136314880;
      9012: inst = 32'd268468224;
      9013: inst = 32'd201345197;
      9014: inst = 32'd203489279;
      9015: inst = 32'd136314880;
      9016: inst = 32'd268468224;
      9017: inst = 32'd201345198;
      9018: inst = 32'd203489279;
      9019: inst = 32'd136314880;
      9020: inst = 32'd268468224;
      9021: inst = 32'd201345199;
      9022: inst = 32'd203489279;
      9023: inst = 32'd136314880;
      9024: inst = 32'd268468224;
      9025: inst = 32'd201345200;
      9026: inst = 32'd203489279;
      9027: inst = 32'd136314880;
      9028: inst = 32'd268468224;
      9029: inst = 32'd201345201;
      9030: inst = 32'd203489279;
      9031: inst = 32'd136314880;
      9032: inst = 32'd268468224;
      9033: inst = 32'd201345202;
      9034: inst = 32'd203489279;
      9035: inst = 32'd136314880;
      9036: inst = 32'd268468224;
      9037: inst = 32'd201345203;
      9038: inst = 32'd203489279;
      9039: inst = 32'd136314880;
      9040: inst = 32'd268468224;
      9041: inst = 32'd201345204;
      9042: inst = 32'd203489279;
      9043: inst = 32'd136314880;
      9044: inst = 32'd268468224;
      9045: inst = 32'd201345205;
      9046: inst = 32'd203489279;
      9047: inst = 32'd136314880;
      9048: inst = 32'd268468224;
      9049: inst = 32'd201345206;
      9050: inst = 32'd203489279;
      9051: inst = 32'd136314880;
      9052: inst = 32'd268468224;
      9053: inst = 32'd201345207;
      9054: inst = 32'd203489279;
      9055: inst = 32'd136314880;
      9056: inst = 32'd268468224;
      9057: inst = 32'd201345208;
      9058: inst = 32'd203489279;
      9059: inst = 32'd136314880;
      9060: inst = 32'd268468224;
      9061: inst = 32'd201345209;
      9062: inst = 32'd203489279;
      9063: inst = 32'd136314880;
      9064: inst = 32'd268468224;
      9065: inst = 32'd201345210;
      9066: inst = 32'd203489279;
      9067: inst = 32'd136314880;
      9068: inst = 32'd268468224;
      9069: inst = 32'd201345211;
      9070: inst = 32'd203489279;
      9071: inst = 32'd136314880;
      9072: inst = 32'd268468224;
      9073: inst = 32'd201345212;
      9074: inst = 32'd203489279;
      9075: inst = 32'd136314880;
      9076: inst = 32'd268468224;
      9077: inst = 32'd201345213;
      9078: inst = 32'd203489279;
      9079: inst = 32'd136314880;
      9080: inst = 32'd268468224;
      9081: inst = 32'd201345214;
      9082: inst = 32'd203489279;
      9083: inst = 32'd136314880;
      9084: inst = 32'd268468224;
      9085: inst = 32'd201345215;
      9086: inst = 32'd203489279;
      9087: inst = 32'd136314880;
      9088: inst = 32'd268468224;
      9089: inst = 32'd201345216;
      9090: inst = 32'd203489279;
      9091: inst = 32'd136314880;
      9092: inst = 32'd268468224;
      9093: inst = 32'd201345217;
      9094: inst = 32'd203489279;
      9095: inst = 32'd136314880;
      9096: inst = 32'd268468224;
      9097: inst = 32'd201345218;
      9098: inst = 32'd203489247;
      9099: inst = 32'd136314880;
      9100: inst = 32'd268468224;
      9101: inst = 32'd201345219;
      9102: inst = 32'd203489279;
      9103: inst = 32'd136314880;
      9104: inst = 32'd268468224;
      9105: inst = 32'd201345220;
      9106: inst = 32'd203482840;
      9107: inst = 32'd136314880;
      9108: inst = 32'd268468224;
      9109: inst = 32'd201345221;
      9110: inst = 32'd203484886;
      9111: inst = 32'd136314880;
      9112: inst = 32'd268468224;
      9113: inst = 32'd201345222;
      9114: inst = 32'd203486869;
      9115: inst = 32'd136314880;
      9116: inst = 32'd268468224;
      9117: inst = 32'd201345223;
      9118: inst = 32'd203484854;
      9119: inst = 32'd136314880;
      9120: inst = 32'd268468224;
      9121: inst = 32'd201345224;
      9122: inst = 32'd203484854;
      9123: inst = 32'd136314880;
      9124: inst = 32'd268468224;
      9125: inst = 32'd201345225;
      9126: inst = 32'd203484822;
      9127: inst = 32'd136314880;
      9128: inst = 32'd268468224;
      9129: inst = 32'd201345226;
      9130: inst = 32'd203488983;
      9131: inst = 32'd136314880;
      9132: inst = 32'd268468224;
      9133: inst = 32'd201345227;
      9134: inst = 32'd203484790;
      9135: inst = 32'd136314880;
      9136: inst = 32'd268468224;
      9137: inst = 32'd201345228;
      9138: inst = 32'd203482806;
      9139: inst = 32'd136314880;
      9140: inst = 32'd268468224;
      9141: inst = 32'd201345229;
      9142: inst = 32'd203484886;
      9143: inst = 32'd136314880;
      9144: inst = 32'd268468224;
      9145: inst = 32'd201345230;
      9146: inst = 32'd203488883;
      9147: inst = 32'd136314880;
      9148: inst = 32'd268468224;
      9149: inst = 32'd201345231;
      9150: inst = 32'd203469541;
      9151: inst = 32'd136314880;
      9152: inst = 32'd268468224;
      9153: inst = 32'd201345232;
      9154: inst = 32'd203482022;
      9155: inst = 32'd136314880;
      9156: inst = 32'd268468224;
      9157: inst = 32'd201345233;
      9158: inst = 32'd203479975;
      9159: inst = 32'd136314880;
      9160: inst = 32'd268468224;
      9161: inst = 32'd201345234;
      9162: inst = 32'd203477960;
      9163: inst = 32'd136314880;
      9164: inst = 32'd268468224;
      9165: inst = 32'd201345235;
      9166: inst = 32'd203475913;
      9167: inst = 32'd136314880;
      9168: inst = 32'd268468224;
      9169: inst = 32'd201345236;
      9170: inst = 32'd203475912;
      9171: inst = 32'd136314880;
      9172: inst = 32'd268468224;
      9173: inst = 32'd201345237;
      9174: inst = 32'd203477959;
      9175: inst = 32'd136314880;
      9176: inst = 32'd268468224;
      9177: inst = 32'd201345238;
      9178: inst = 32'd203480006;
      9179: inst = 32'd136314880;
      9180: inst = 32'd268468224;
      9181: inst = 32'd201345239;
      9182: inst = 32'd203480006;
      9183: inst = 32'd136314880;
      9184: inst = 32'd268468224;
      9185: inst = 32'd201345240;
      9186: inst = 32'd203480006;
      9187: inst = 32'd136314880;
      9188: inst = 32'd268468224;
      9189: inst = 32'd201345241;
      9190: inst = 32'd203480006;
      9191: inst = 32'd136314880;
      9192: inst = 32'd268468224;
      9193: inst = 32'd201345242;
      9194: inst = 32'd203480005;
      9195: inst = 32'd136314880;
      9196: inst = 32'd268468224;
      9197: inst = 32'd201345243;
      9198: inst = 32'd203480037;
      9199: inst = 32'd136314880;
      9200: inst = 32'd268468224;
      9201: inst = 32'd201345244;
      9202: inst = 32'd203479972;
      9203: inst = 32'd136314880;
      9204: inst = 32'd268468224;
      9205: inst = 32'd201345245;
      9206: inst = 32'd203482085;
      9207: inst = 32'd136314880;
      9208: inst = 32'd268468224;
      9209: inst = 32'd201345246;
      9210: inst = 32'd203480037;
      9211: inst = 32'd136314880;
      9212: inst = 32'd268468224;
      9213: inst = 32'd201345247;
      9214: inst = 32'd203471586;
      9215: inst = 32'd136314880;
      9216: inst = 32'd268468224;
      9217: inst = 32'd201345248;
      9218: inst = 32'd203484854;
      9219: inst = 32'd136314880;
      9220: inst = 32'd268468224;
      9221: inst = 32'd201345249;
      9222: inst = 32'd203484854;
      9223: inst = 32'd136314880;
      9224: inst = 32'd268468224;
      9225: inst = 32'd201345250;
      9226: inst = 32'd203484854;
      9227: inst = 32'd136314880;
      9228: inst = 32'd268468224;
      9229: inst = 32'd201345251;
      9230: inst = 32'd203484854;
      9231: inst = 32'd136314880;
      9232: inst = 32'd268468224;
      9233: inst = 32'd201345252;
      9234: inst = 32'd203484886;
      9235: inst = 32'd136314880;
      9236: inst = 32'd268468224;
      9237: inst = 32'd201345253;
      9238: inst = 32'd203484886;
      9239: inst = 32'd136314880;
      9240: inst = 32'd268468224;
      9241: inst = 32'd201345254;
      9242: inst = 32'd203484854;
      9243: inst = 32'd136314880;
      9244: inst = 32'd268468224;
      9245: inst = 32'd201345255;
      9246: inst = 32'd203484854;
      9247: inst = 32'd136314880;
      9248: inst = 32'd268468224;
      9249: inst = 32'd201345256;
      9250: inst = 32'd203484855;
      9251: inst = 32'd136314880;
      9252: inst = 32'd268468224;
      9253: inst = 32'd201345257;
      9254: inst = 32'd203486935;
      9255: inst = 32'd136314880;
      9256: inst = 32'd268468224;
      9257: inst = 32'd201345258;
      9258: inst = 32'd203484855;
      9259: inst = 32'd136314880;
      9260: inst = 32'd268468224;
      9261: inst = 32'd201345259;
      9262: inst = 32'd203484855;
      9263: inst = 32'd136314880;
      9264: inst = 32'd268468224;
      9265: inst = 32'd201345260;
      9266: inst = 32'd203482742;
      9267: inst = 32'd136314880;
      9268: inst = 32'd268468224;
      9269: inst = 32'd201345261;
      9270: inst = 32'd203486967;
      9271: inst = 32'd136314880;
      9272: inst = 32'd268468224;
      9273: inst = 32'd201345262;
      9274: inst = 32'd203484854;
      9275: inst = 32'd136314880;
      9276: inst = 32'd268468224;
      9277: inst = 32'd201345263;
      9278: inst = 32'd203484886;
      9279: inst = 32'd136314880;
      9280: inst = 32'd268468224;
      9281: inst = 32'd201345264;
      9282: inst = 32'd203484854;
      9283: inst = 32'd136314880;
      9284: inst = 32'd268468224;
      9285: inst = 32'd201345265;
      9286: inst = 32'd203484854;
      9287: inst = 32'd136314880;
      9288: inst = 32'd268468224;
      9289: inst = 32'd201345266;
      9290: inst = 32'd203484854;
      9291: inst = 32'd136314880;
      9292: inst = 32'd268468224;
      9293: inst = 32'd201345267;
      9294: inst = 32'd203484854;
      9295: inst = 32'd136314880;
      9296: inst = 32'd268468224;
      9297: inst = 32'd201345268;
      9298: inst = 32'd203484854;
      9299: inst = 32'd136314880;
      9300: inst = 32'd268468224;
      9301: inst = 32'd201345269;
      9302: inst = 32'd203484854;
      9303: inst = 32'd136314880;
      9304: inst = 32'd268468224;
      9305: inst = 32'd201345270;
      9306: inst = 32'd203484854;
      9307: inst = 32'd136314880;
      9308: inst = 32'd268468224;
      9309: inst = 32'd201345271;
      9310: inst = 32'd203484854;
      9311: inst = 32'd136314880;
      9312: inst = 32'd268468224;
      9313: inst = 32'd201345272;
      9314: inst = 32'd203484854;
      9315: inst = 32'd136314880;
      9316: inst = 32'd268468224;
      9317: inst = 32'd201345273;
      9318: inst = 32'd203484854;
      9319: inst = 32'd136314880;
      9320: inst = 32'd268468224;
      9321: inst = 32'd201345274;
      9322: inst = 32'd203484855;
      9323: inst = 32'd136314880;
      9324: inst = 32'd268468224;
      9325: inst = 32'd201345275;
      9326: inst = 32'd203482808;
      9327: inst = 32'd136314880;
      9328: inst = 32'd268468224;
      9329: inst = 32'd201345276;
      9330: inst = 32'd203489278;
      9331: inst = 32'd136314880;
      9332: inst = 32'd268468224;
      9333: inst = 32'd201345277;
      9334: inst = 32'd203489279;
      9335: inst = 32'd136314880;
      9336: inst = 32'd268468224;
      9337: inst = 32'd201345278;
      9338: inst = 32'd203489279;
      9339: inst = 32'd136314880;
      9340: inst = 32'd268468224;
      9341: inst = 32'd201345279;
      9342: inst = 32'd203489279;
      9343: inst = 32'd136314880;
      9344: inst = 32'd268468224;
      9345: inst = 32'd201345280;
      9346: inst = 32'd203489279;
      9347: inst = 32'd136314880;
      9348: inst = 32'd268468224;
      9349: inst = 32'd201345281;
      9350: inst = 32'd203489279;
      9351: inst = 32'd136314880;
      9352: inst = 32'd268468224;
      9353: inst = 32'd201345282;
      9354: inst = 32'd203489279;
      9355: inst = 32'd136314880;
      9356: inst = 32'd268468224;
      9357: inst = 32'd201345283;
      9358: inst = 32'd203489279;
      9359: inst = 32'd136314880;
      9360: inst = 32'd268468224;
      9361: inst = 32'd201345284;
      9362: inst = 32'd203489279;
      9363: inst = 32'd136314880;
      9364: inst = 32'd268468224;
      9365: inst = 32'd201345285;
      9366: inst = 32'd203489279;
      9367: inst = 32'd136314880;
      9368: inst = 32'd268468224;
      9369: inst = 32'd201345286;
      9370: inst = 32'd203489279;
      9371: inst = 32'd136314880;
      9372: inst = 32'd268468224;
      9373: inst = 32'd201345287;
      9374: inst = 32'd203489279;
      9375: inst = 32'd136314880;
      9376: inst = 32'd268468224;
      9377: inst = 32'd201345288;
      9378: inst = 32'd203489279;
      9379: inst = 32'd136314880;
      9380: inst = 32'd268468224;
      9381: inst = 32'd201345289;
      9382: inst = 32'd203489279;
      9383: inst = 32'd136314880;
      9384: inst = 32'd268468224;
      9385: inst = 32'd201345290;
      9386: inst = 32'd203489279;
      9387: inst = 32'd136314880;
      9388: inst = 32'd268468224;
      9389: inst = 32'd201345291;
      9390: inst = 32'd203489279;
      9391: inst = 32'd136314880;
      9392: inst = 32'd268468224;
      9393: inst = 32'd201345292;
      9394: inst = 32'd203489279;
      9395: inst = 32'd136314880;
      9396: inst = 32'd268468224;
      9397: inst = 32'd201345293;
      9398: inst = 32'd203489279;
      9399: inst = 32'd136314880;
      9400: inst = 32'd268468224;
      9401: inst = 32'd201345294;
      9402: inst = 32'd203489279;
      9403: inst = 32'd136314880;
      9404: inst = 32'd268468224;
      9405: inst = 32'd201345295;
      9406: inst = 32'd203489279;
      9407: inst = 32'd136314880;
      9408: inst = 32'd268468224;
      9409: inst = 32'd201345296;
      9410: inst = 32'd203489279;
      9411: inst = 32'd136314880;
      9412: inst = 32'd268468224;
      9413: inst = 32'd201345297;
      9414: inst = 32'd203489279;
      9415: inst = 32'd136314880;
      9416: inst = 32'd268468224;
      9417: inst = 32'd201345298;
      9418: inst = 32'd203489279;
      9419: inst = 32'd136314880;
      9420: inst = 32'd268468224;
      9421: inst = 32'd201345299;
      9422: inst = 32'd203489279;
      9423: inst = 32'd136314880;
      9424: inst = 32'd268468224;
      9425: inst = 32'd201345300;
      9426: inst = 32'd203489279;
      9427: inst = 32'd136314880;
      9428: inst = 32'd268468224;
      9429: inst = 32'd201345301;
      9430: inst = 32'd203489279;
      9431: inst = 32'd136314880;
      9432: inst = 32'd268468224;
      9433: inst = 32'd201345302;
      9434: inst = 32'd203489279;
      9435: inst = 32'd136314880;
      9436: inst = 32'd268468224;
      9437: inst = 32'd201345303;
      9438: inst = 32'd203489279;
      9439: inst = 32'd136314880;
      9440: inst = 32'd268468224;
      9441: inst = 32'd201345304;
      9442: inst = 32'd203489279;
      9443: inst = 32'd136314880;
      9444: inst = 32'd268468224;
      9445: inst = 32'd201345305;
      9446: inst = 32'd203489279;
      9447: inst = 32'd136314880;
      9448: inst = 32'd268468224;
      9449: inst = 32'd201345306;
      9450: inst = 32'd203489279;
      9451: inst = 32'd136314880;
      9452: inst = 32'd268468224;
      9453: inst = 32'd201345307;
      9454: inst = 32'd203489279;
      9455: inst = 32'd136314880;
      9456: inst = 32'd268468224;
      9457: inst = 32'd201345308;
      9458: inst = 32'd203489279;
      9459: inst = 32'd136314880;
      9460: inst = 32'd268468224;
      9461: inst = 32'd201345309;
      9462: inst = 32'd203489279;
      9463: inst = 32'd136314880;
      9464: inst = 32'd268468224;
      9465: inst = 32'd201345310;
      9466: inst = 32'd203489279;
      9467: inst = 32'd136314880;
      9468: inst = 32'd268468224;
      9469: inst = 32'd201345311;
      9470: inst = 32'd203489279;
      9471: inst = 32'd136314880;
      9472: inst = 32'd268468224;
      9473: inst = 32'd201345312;
      9474: inst = 32'd203489279;
      9475: inst = 32'd136314880;
      9476: inst = 32'd268468224;
      9477: inst = 32'd201345313;
      9478: inst = 32'd203489279;
      9479: inst = 32'd136314880;
      9480: inst = 32'd268468224;
      9481: inst = 32'd201345314;
      9482: inst = 32'd203489247;
      9483: inst = 32'd136314880;
      9484: inst = 32'd268468224;
      9485: inst = 32'd201345315;
      9486: inst = 32'd203489279;
      9487: inst = 32'd136314880;
      9488: inst = 32'd268468224;
      9489: inst = 32'd201345316;
      9490: inst = 32'd203482840;
      9491: inst = 32'd136314880;
      9492: inst = 32'd268468224;
      9493: inst = 32'd201345317;
      9494: inst = 32'd203484886;
      9495: inst = 32'd136314880;
      9496: inst = 32'd268468224;
      9497: inst = 32'd201345318;
      9498: inst = 32'd203486901;
      9499: inst = 32'd136314880;
      9500: inst = 32'd268468224;
      9501: inst = 32'd201345319;
      9502: inst = 32'd203484854;
      9503: inst = 32'd136314880;
      9504: inst = 32'd268468224;
      9505: inst = 32'd201345320;
      9506: inst = 32'd203484886;
      9507: inst = 32'd136314880;
      9508: inst = 32'd268468224;
      9509: inst = 32'd201345321;
      9510: inst = 32'd203484854;
      9511: inst = 32'd136314880;
      9512: inst = 32'd268468224;
      9513: inst = 32'd201345322;
      9514: inst = 32'd203486870;
      9515: inst = 32'd136314880;
      9516: inst = 32'd268468224;
      9517: inst = 32'd201345323;
      9518: inst = 32'd203486870;
      9519: inst = 32'd136314880;
      9520: inst = 32'd268468224;
      9521: inst = 32'd201345324;
      9522: inst = 32'd203484887;
      9523: inst = 32'd136314880;
      9524: inst = 32'd268468224;
      9525: inst = 32'd201345325;
      9526: inst = 32'd203484886;
      9527: inst = 32'd136314880;
      9528: inst = 32'd268468224;
      9529: inst = 32'd201345326;
      9530: inst = 32'd203488915;
      9531: inst = 32'd136314880;
      9532: inst = 32'd268468224;
      9533: inst = 32'd201345327;
      9534: inst = 32'd203469573;
      9535: inst = 32'd136314880;
      9536: inst = 32'd268468224;
      9537: inst = 32'd201345328;
      9538: inst = 32'd203482054;
      9539: inst = 32'd136314880;
      9540: inst = 32'd268468224;
      9541: inst = 32'd201345329;
      9542: inst = 32'd203473864;
      9543: inst = 32'd136314880;
      9544: inst = 32'd268468224;
      9545: inst = 32'd201345330;
      9546: inst = 32'd203489144;
      9547: inst = 32'd136314880;
      9548: inst = 32'd268468224;
      9549: inst = 32'd201345331;
      9550: inst = 32'd203487097;
      9551: inst = 32'd136314880;
      9552: inst = 32'd268468224;
      9553: inst = 32'd201345332;
      9554: inst = 32'd203489113;
      9555: inst = 32'd136314880;
      9556: inst = 32'd268468224;
      9557: inst = 32'd201345333;
      9558: inst = 32'd203489079;
      9559: inst = 32'd136314880;
      9560: inst = 32'd268468224;
      9561: inst = 32'd201345334;
      9562: inst = 32'd203475880;
      9563: inst = 32'd136314880;
      9564: inst = 32'd268468224;
      9565: inst = 32'd201345335;
      9566: inst = 32'd203482023;
      9567: inst = 32'd136314880;
      9568: inst = 32'd268468224;
      9569: inst = 32'd201345336;
      9570: inst = 32'd203482022;
      9571: inst = 32'd136314880;
      9572: inst = 32'd268468224;
      9573: inst = 32'd201345337;
      9574: inst = 32'd203480006;
      9575: inst = 32'd136314880;
      9576: inst = 32'd268468224;
      9577: inst = 32'd201345338;
      9578: inst = 32'd203477958;
      9579: inst = 32'd136314880;
      9580: inst = 32'd268468224;
      9581: inst = 32'd201345339;
      9582: inst = 32'd203480038;
      9583: inst = 32'd136314880;
      9584: inst = 32'd268468224;
      9585: inst = 32'd201345340;
      9586: inst = 32'd203480005;
      9587: inst = 32'd136314880;
      9588: inst = 32'd268468224;
      9589: inst = 32'd201345341;
      9590: inst = 32'd203482022;
      9591: inst = 32'd136314880;
      9592: inst = 32'd268468224;
      9593: inst = 32'd201345342;
      9594: inst = 32'd203481990;
      9595: inst = 32'd136314880;
      9596: inst = 32'd268468224;
      9597: inst = 32'd201345343;
      9598: inst = 32'd203475652;
      9599: inst = 32'd136314880;
      9600: inst = 32'd268468224;
      9601: inst = 32'd201345344;
      9602: inst = 32'd203484854;
      9603: inst = 32'd136314880;
      9604: inst = 32'd268468224;
      9605: inst = 32'd201345345;
      9606: inst = 32'd203484854;
      9607: inst = 32'd136314880;
      9608: inst = 32'd268468224;
      9609: inst = 32'd201345346;
      9610: inst = 32'd203484854;
      9611: inst = 32'd136314880;
      9612: inst = 32'd268468224;
      9613: inst = 32'd201345347;
      9614: inst = 32'd203484885;
      9615: inst = 32'd136314880;
      9616: inst = 32'd268468224;
      9617: inst = 32'd201345348;
      9618: inst = 32'd203484885;
      9619: inst = 32'd136314880;
      9620: inst = 32'd268468224;
      9621: inst = 32'd201345349;
      9622: inst = 32'd203484886;
      9623: inst = 32'd136314880;
      9624: inst = 32'd268468224;
      9625: inst = 32'd201345350;
      9626: inst = 32'd203484854;
      9627: inst = 32'd136314880;
      9628: inst = 32'd268468224;
      9629: inst = 32'd201345351;
      9630: inst = 32'd203484854;
      9631: inst = 32'd136314880;
      9632: inst = 32'd268468224;
      9633: inst = 32'd201345352;
      9634: inst = 32'd203482774;
      9635: inst = 32'd136314880;
      9636: inst = 32'd268468224;
      9637: inst = 32'd201345353;
      9638: inst = 32'd203484888;
      9639: inst = 32'd136314880;
      9640: inst = 32'd268468224;
      9641: inst = 32'd201345354;
      9642: inst = 32'd203484855;
      9643: inst = 32'd136314880;
      9644: inst = 32'd268468224;
      9645: inst = 32'd201345355;
      9646: inst = 32'd203486968;
      9647: inst = 32'd136314880;
      9648: inst = 32'd268468224;
      9649: inst = 32'd201345356;
      9650: inst = 32'd203484887;
      9651: inst = 32'd136314880;
      9652: inst = 32'd268468224;
      9653: inst = 32'd201345357;
      9654: inst = 32'd203482774;
      9655: inst = 32'd136314880;
      9656: inst = 32'd268468224;
      9657: inst = 32'd201345358;
      9658: inst = 32'd203482806;
      9659: inst = 32'd136314880;
      9660: inst = 32'd268468224;
      9661: inst = 32'd201345359;
      9662: inst = 32'd203484854;
      9663: inst = 32'd136314880;
      9664: inst = 32'd268468224;
      9665: inst = 32'd201345360;
      9666: inst = 32'd203484854;
      9667: inst = 32'd136314880;
      9668: inst = 32'd268468224;
      9669: inst = 32'd201345361;
      9670: inst = 32'd203484854;
      9671: inst = 32'd136314880;
      9672: inst = 32'd268468224;
      9673: inst = 32'd201345362;
      9674: inst = 32'd203484854;
      9675: inst = 32'd136314880;
      9676: inst = 32'd268468224;
      9677: inst = 32'd201345363;
      9678: inst = 32'd203484854;
      9679: inst = 32'd136314880;
      9680: inst = 32'd268468224;
      9681: inst = 32'd201345364;
      9682: inst = 32'd203484854;
      9683: inst = 32'd136314880;
      9684: inst = 32'd268468224;
      9685: inst = 32'd201345365;
      9686: inst = 32'd203484854;
      9687: inst = 32'd136314880;
      9688: inst = 32'd268468224;
      9689: inst = 32'd201345366;
      9690: inst = 32'd203484854;
      9691: inst = 32'd136314880;
      9692: inst = 32'd268468224;
      9693: inst = 32'd201345367;
      9694: inst = 32'd203484854;
      9695: inst = 32'd136314880;
      9696: inst = 32'd268468224;
      9697: inst = 32'd201345368;
      9698: inst = 32'd203484854;
      9699: inst = 32'd136314880;
      9700: inst = 32'd268468224;
      9701: inst = 32'd201345369;
      9702: inst = 32'd203484854;
      9703: inst = 32'd136314880;
      9704: inst = 32'd268468224;
      9705: inst = 32'd201345370;
      9706: inst = 32'd203484855;
      9707: inst = 32'd136314880;
      9708: inst = 32'd268468224;
      9709: inst = 32'd201345371;
      9710: inst = 32'd203482808;
      9711: inst = 32'd136314880;
      9712: inst = 32'd268468224;
      9713: inst = 32'd201345372;
      9714: inst = 32'd203489278;
      9715: inst = 32'd136314880;
      9716: inst = 32'd268468224;
      9717: inst = 32'd201345373;
      9718: inst = 32'd203489279;
      9719: inst = 32'd136314880;
      9720: inst = 32'd268468224;
      9721: inst = 32'd201345374;
      9722: inst = 32'd203489279;
      9723: inst = 32'd136314880;
      9724: inst = 32'd268468224;
      9725: inst = 32'd201345375;
      9726: inst = 32'd203489279;
      9727: inst = 32'd136314880;
      9728: inst = 32'd268468224;
      9729: inst = 32'd201345376;
      9730: inst = 32'd203489279;
      9731: inst = 32'd136314880;
      9732: inst = 32'd268468224;
      9733: inst = 32'd201345377;
      9734: inst = 32'd203489279;
      9735: inst = 32'd136314880;
      9736: inst = 32'd268468224;
      9737: inst = 32'd201345378;
      9738: inst = 32'd203489279;
      9739: inst = 32'd136314880;
      9740: inst = 32'd268468224;
      9741: inst = 32'd201345379;
      9742: inst = 32'd203489279;
      9743: inst = 32'd136314880;
      9744: inst = 32'd268468224;
      9745: inst = 32'd201345380;
      9746: inst = 32'd203489279;
      9747: inst = 32'd136314880;
      9748: inst = 32'd268468224;
      9749: inst = 32'd201345381;
      9750: inst = 32'd203489279;
      9751: inst = 32'd136314880;
      9752: inst = 32'd268468224;
      9753: inst = 32'd201345382;
      9754: inst = 32'd203489279;
      9755: inst = 32'd136314880;
      9756: inst = 32'd268468224;
      9757: inst = 32'd201345383;
      9758: inst = 32'd203489279;
      9759: inst = 32'd136314880;
      9760: inst = 32'd268468224;
      9761: inst = 32'd201345384;
      9762: inst = 32'd203489279;
      9763: inst = 32'd136314880;
      9764: inst = 32'd268468224;
      9765: inst = 32'd201345385;
      9766: inst = 32'd203489279;
      9767: inst = 32'd136314880;
      9768: inst = 32'd268468224;
      9769: inst = 32'd201345386;
      9770: inst = 32'd203489279;
      9771: inst = 32'd136314880;
      9772: inst = 32'd268468224;
      9773: inst = 32'd201345387;
      9774: inst = 32'd203489279;
      9775: inst = 32'd136314880;
      9776: inst = 32'd268468224;
      9777: inst = 32'd201345388;
      9778: inst = 32'd203489279;
      9779: inst = 32'd136314880;
      9780: inst = 32'd268468224;
      9781: inst = 32'd201345389;
      9782: inst = 32'd203489279;
      9783: inst = 32'd136314880;
      9784: inst = 32'd268468224;
      9785: inst = 32'd201345390;
      9786: inst = 32'd203489279;
      9787: inst = 32'd136314880;
      9788: inst = 32'd268468224;
      9789: inst = 32'd201345391;
      9790: inst = 32'd203489279;
      9791: inst = 32'd136314880;
      9792: inst = 32'd268468224;
      9793: inst = 32'd201345392;
      9794: inst = 32'd203489279;
      9795: inst = 32'd136314880;
      9796: inst = 32'd268468224;
      9797: inst = 32'd201345393;
      9798: inst = 32'd203489279;
      9799: inst = 32'd136314880;
      9800: inst = 32'd268468224;
      9801: inst = 32'd201345394;
      9802: inst = 32'd203489279;
      9803: inst = 32'd136314880;
      9804: inst = 32'd268468224;
      9805: inst = 32'd201345395;
      9806: inst = 32'd203489279;
      9807: inst = 32'd136314880;
      9808: inst = 32'd268468224;
      9809: inst = 32'd201345396;
      9810: inst = 32'd203489279;
      9811: inst = 32'd136314880;
      9812: inst = 32'd268468224;
      9813: inst = 32'd201345397;
      9814: inst = 32'd203489279;
      9815: inst = 32'd136314880;
      9816: inst = 32'd268468224;
      9817: inst = 32'd201345398;
      9818: inst = 32'd203489279;
      9819: inst = 32'd136314880;
      9820: inst = 32'd268468224;
      9821: inst = 32'd201345399;
      9822: inst = 32'd203489279;
      9823: inst = 32'd136314880;
      9824: inst = 32'd268468224;
      9825: inst = 32'd201345400;
      9826: inst = 32'd203489279;
      9827: inst = 32'd136314880;
      9828: inst = 32'd268468224;
      9829: inst = 32'd201345401;
      9830: inst = 32'd203489279;
      9831: inst = 32'd136314880;
      9832: inst = 32'd268468224;
      9833: inst = 32'd201345402;
      9834: inst = 32'd203489279;
      9835: inst = 32'd136314880;
      9836: inst = 32'd268468224;
      9837: inst = 32'd201345403;
      9838: inst = 32'd203489279;
      9839: inst = 32'd136314880;
      9840: inst = 32'd268468224;
      9841: inst = 32'd201345404;
      9842: inst = 32'd203489279;
      9843: inst = 32'd136314880;
      9844: inst = 32'd268468224;
      9845: inst = 32'd201345405;
      9846: inst = 32'd203489279;
      9847: inst = 32'd136314880;
      9848: inst = 32'd268468224;
      9849: inst = 32'd201345406;
      9850: inst = 32'd203489279;
      9851: inst = 32'd136314880;
      9852: inst = 32'd268468224;
      9853: inst = 32'd201345407;
      9854: inst = 32'd203489279;
      9855: inst = 32'd136314880;
      9856: inst = 32'd268468224;
      9857: inst = 32'd201345408;
      9858: inst = 32'd203489279;
      9859: inst = 32'd136314880;
      9860: inst = 32'd268468224;
      9861: inst = 32'd201345409;
      9862: inst = 32'd203489279;
      9863: inst = 32'd136314880;
      9864: inst = 32'd268468224;
      9865: inst = 32'd201345410;
      9866: inst = 32'd203489247;
      9867: inst = 32'd136314880;
      9868: inst = 32'd268468224;
      9869: inst = 32'd201345411;
      9870: inst = 32'd203489279;
      9871: inst = 32'd136314880;
      9872: inst = 32'd268468224;
      9873: inst = 32'd201345412;
      9874: inst = 32'd203482840;
      9875: inst = 32'd136314880;
      9876: inst = 32'd268468224;
      9877: inst = 32'd201345413;
      9878: inst = 32'd203484886;
      9879: inst = 32'd136314880;
      9880: inst = 32'd268468224;
      9881: inst = 32'd201345414;
      9882: inst = 32'd203486901;
      9883: inst = 32'd136314880;
      9884: inst = 32'd268468224;
      9885: inst = 32'd201345415;
      9886: inst = 32'd203484854;
      9887: inst = 32'd136314880;
      9888: inst = 32'd268468224;
      9889: inst = 32'd201345416;
      9890: inst = 32'd203484886;
      9891: inst = 32'd136314880;
      9892: inst = 32'd268468224;
      9893: inst = 32'd201345417;
      9894: inst = 32'd203484854;
      9895: inst = 32'd136314880;
      9896: inst = 32'd268468224;
      9897: inst = 32'd201345418;
      9898: inst = 32'd203486870;
      9899: inst = 32'd136314880;
      9900: inst = 32'd268468224;
      9901: inst = 32'd201345419;
      9902: inst = 32'd203486870;
      9903: inst = 32'd136314880;
      9904: inst = 32'd268468224;
      9905: inst = 32'd201345420;
      9906: inst = 32'd203484887;
      9907: inst = 32'd136314880;
      9908: inst = 32'd268468224;
      9909: inst = 32'd201345421;
      9910: inst = 32'd203484886;
      9911: inst = 32'd136314880;
      9912: inst = 32'd268468224;
      9913: inst = 32'd201345422;
      9914: inst = 32'd203488883;
      9915: inst = 32'd136314880;
      9916: inst = 32'd268468224;
      9917: inst = 32'd201345423;
      9918: inst = 32'd203471621;
      9919: inst = 32'd136314880;
      9920: inst = 32'd268468224;
      9921: inst = 32'd201345424;
      9922: inst = 32'd203481988;
      9923: inst = 32'd136314880;
      9924: inst = 32'd268468224;
      9925: inst = 32'd201345425;
      9926: inst = 32'd203473961;
      9927: inst = 32'd136314880;
      9928: inst = 32'd268468224;
      9929: inst = 32'd201345426;
      9930: inst = 32'd203489242;
      9931: inst = 32'd136314880;
      9932: inst = 32'd268468224;
      9933: inst = 32'd201345427;
      9934: inst = 32'd203481084;
      9935: inst = 32'd136314880;
      9936: inst = 32'd268468224;
      9937: inst = 32'd201345428;
      9938: inst = 32'd203483068;
      9939: inst = 32'd136314880;
      9940: inst = 32'd268468224;
      9941: inst = 32'd201345429;
      9942: inst = 32'd203489080;
      9943: inst = 32'd136314880;
      9944: inst = 32'd268468224;
      9945: inst = 32'd201345430;
      9946: inst = 32'd203475945;
      9947: inst = 32'd136314880;
      9948: inst = 32'd268468224;
      9949: inst = 32'd201345431;
      9950: inst = 32'd203481990;
      9951: inst = 32'd136314880;
      9952: inst = 32'd268468224;
      9953: inst = 32'd201345432;
      9954: inst = 32'd203484069;
      9955: inst = 32'd136314880;
      9956: inst = 32'd268468224;
      9957: inst = 32'd201345433;
      9958: inst = 32'd203480005;
      9959: inst = 32'd136314880;
      9960: inst = 32'd268468224;
      9961: inst = 32'd201345434;
      9962: inst = 32'd203477957;
      9963: inst = 32'd136314880;
      9964: inst = 32'd268468224;
      9965: inst = 32'd201345435;
      9966: inst = 32'd203480006;
      9967: inst = 32'd136314880;
      9968: inst = 32'd268468224;
      9969: inst = 32'd201345436;
      9970: inst = 32'd203482021;
      9971: inst = 32'd136314880;
      9972: inst = 32'd268468224;
      9973: inst = 32'd201345437;
      9974: inst = 32'd203482022;
      9975: inst = 32'd136314880;
      9976: inst = 32'd268468224;
      9977: inst = 32'd201345438;
      9978: inst = 32'd203481990;
      9979: inst = 32'd136314880;
      9980: inst = 32'd268468224;
      9981: inst = 32'd201345439;
      9982: inst = 32'd203475620;
      9983: inst = 32'd136314880;
      9984: inst = 32'd268468224;
      9985: inst = 32'd201345440;
      9986: inst = 32'd203484854;
      9987: inst = 32'd136314880;
      9988: inst = 32'd268468224;
      9989: inst = 32'd201345441;
      9990: inst = 32'd203484854;
      9991: inst = 32'd136314880;
      9992: inst = 32'd268468224;
      9993: inst = 32'd201345442;
      9994: inst = 32'd203484854;
      9995: inst = 32'd136314880;
      9996: inst = 32'd268468224;
      9997: inst = 32'd201345443;
      9998: inst = 32'd203484853;
      9999: inst = 32'd136314880;
      10000: inst = 32'd268468224;
      10001: inst = 32'd201345444;
      10002: inst = 32'd203484885;
      10003: inst = 32'd136314880;
      10004: inst = 32'd268468224;
      10005: inst = 32'd201345445;
      10006: inst = 32'd203484885;
      10007: inst = 32'd136314880;
      10008: inst = 32'd268468224;
      10009: inst = 32'd201345446;
      10010: inst = 32'd203484886;
      10011: inst = 32'd136314880;
      10012: inst = 32'd268468224;
      10013: inst = 32'd201345447;
      10014: inst = 32'd203484855;
      10015: inst = 32'd136314880;
      10016: inst = 32'd268468224;
      10017: inst = 32'd201345448;
      10018: inst = 32'd203484888;
      10019: inst = 32'd136314880;
      10020: inst = 32'd268468224;
      10021: inst = 32'd201345449;
      10022: inst = 32'd203484856;
      10023: inst = 32'd136314880;
      10024: inst = 32'd268468224;
      10025: inst = 32'd201345450;
      10026: inst = 32'd203482808;
      10027: inst = 32'd136314880;
      10028: inst = 32'd268468224;
      10029: inst = 32'd201345451;
      10030: inst = 32'd203482776;
      10031: inst = 32'd136314880;
      10032: inst = 32'd268468224;
      10033: inst = 32'd201345452;
      10034: inst = 32'd203484888;
      10035: inst = 32'd136314880;
      10036: inst = 32'd268468224;
      10037: inst = 32'd201345453;
      10038: inst = 32'd203484887;
      10039: inst = 32'd136314880;
      10040: inst = 32'd268468224;
      10041: inst = 32'd201345454;
      10042: inst = 32'd203482806;
      10043: inst = 32'd136314880;
      10044: inst = 32'd268468224;
      10045: inst = 32'd201345455;
      10046: inst = 32'd203482806;
      10047: inst = 32'd136314880;
      10048: inst = 32'd268468224;
      10049: inst = 32'd201345456;
      10050: inst = 32'd203484854;
      10051: inst = 32'd136314880;
      10052: inst = 32'd268468224;
      10053: inst = 32'd201345457;
      10054: inst = 32'd203484854;
      10055: inst = 32'd136314880;
      10056: inst = 32'd268468224;
      10057: inst = 32'd201345458;
      10058: inst = 32'd203484854;
      10059: inst = 32'd136314880;
      10060: inst = 32'd268468224;
      10061: inst = 32'd201345459;
      10062: inst = 32'd203484854;
      10063: inst = 32'd136314880;
      10064: inst = 32'd268468224;
      10065: inst = 32'd201345460;
      10066: inst = 32'd203484854;
      10067: inst = 32'd136314880;
      10068: inst = 32'd268468224;
      10069: inst = 32'd201345461;
      10070: inst = 32'd203484854;
      10071: inst = 32'd136314880;
      10072: inst = 32'd268468224;
      10073: inst = 32'd201345462;
      10074: inst = 32'd203484854;
      10075: inst = 32'd136314880;
      10076: inst = 32'd268468224;
      10077: inst = 32'd201345463;
      10078: inst = 32'd203484854;
      10079: inst = 32'd136314880;
      10080: inst = 32'd268468224;
      10081: inst = 32'd201345464;
      10082: inst = 32'd203484854;
      10083: inst = 32'd136314880;
      10084: inst = 32'd268468224;
      10085: inst = 32'd201345465;
      10086: inst = 32'd203484854;
      10087: inst = 32'd136314880;
      10088: inst = 32'd268468224;
      10089: inst = 32'd201345466;
      10090: inst = 32'd203484855;
      10091: inst = 32'd136314880;
      10092: inst = 32'd268468224;
      10093: inst = 32'd201345467;
      10094: inst = 32'd203482808;
      10095: inst = 32'd136314880;
      10096: inst = 32'd268468224;
      10097: inst = 32'd201345468;
      10098: inst = 32'd203489278;
      10099: inst = 32'd136314880;
      10100: inst = 32'd268468224;
      10101: inst = 32'd201345469;
      10102: inst = 32'd203489279;
      10103: inst = 32'd136314880;
      10104: inst = 32'd268468224;
      10105: inst = 32'd201345470;
      10106: inst = 32'd203489279;
      10107: inst = 32'd136314880;
      10108: inst = 32'd268468224;
      10109: inst = 32'd201345471;
      10110: inst = 32'd203489279;
      10111: inst = 32'd136314880;
      10112: inst = 32'd268468224;
      10113: inst = 32'd201345472;
      10114: inst = 32'd203489279;
      10115: inst = 32'd136314880;
      10116: inst = 32'd268468224;
      10117: inst = 32'd201345473;
      10118: inst = 32'd203489279;
      10119: inst = 32'd136314880;
      10120: inst = 32'd268468224;
      10121: inst = 32'd201345474;
      10122: inst = 32'd203489279;
      10123: inst = 32'd136314880;
      10124: inst = 32'd268468224;
      10125: inst = 32'd201345475;
      10126: inst = 32'd203489279;
      10127: inst = 32'd136314880;
      10128: inst = 32'd268468224;
      10129: inst = 32'd201345476;
      10130: inst = 32'd203489279;
      10131: inst = 32'd136314880;
      10132: inst = 32'd268468224;
      10133: inst = 32'd201345477;
      10134: inst = 32'd203489279;
      10135: inst = 32'd136314880;
      10136: inst = 32'd268468224;
      10137: inst = 32'd201345478;
      10138: inst = 32'd203489279;
      10139: inst = 32'd136314880;
      10140: inst = 32'd268468224;
      10141: inst = 32'd201345479;
      10142: inst = 32'd203489279;
      10143: inst = 32'd136314880;
      10144: inst = 32'd268468224;
      10145: inst = 32'd201345480;
      10146: inst = 32'd203489279;
      10147: inst = 32'd136314880;
      10148: inst = 32'd268468224;
      10149: inst = 32'd201345481;
      10150: inst = 32'd203489279;
      10151: inst = 32'd136314880;
      10152: inst = 32'd268468224;
      10153: inst = 32'd201345482;
      10154: inst = 32'd203489279;
      10155: inst = 32'd136314880;
      10156: inst = 32'd268468224;
      10157: inst = 32'd201345483;
      10158: inst = 32'd203489279;
      10159: inst = 32'd136314880;
      10160: inst = 32'd268468224;
      10161: inst = 32'd201345484;
      10162: inst = 32'd203489279;
      10163: inst = 32'd136314880;
      10164: inst = 32'd268468224;
      10165: inst = 32'd201345485;
      10166: inst = 32'd203489279;
      10167: inst = 32'd136314880;
      10168: inst = 32'd268468224;
      10169: inst = 32'd201345486;
      10170: inst = 32'd203489279;
      10171: inst = 32'd136314880;
      10172: inst = 32'd268468224;
      10173: inst = 32'd201345487;
      10174: inst = 32'd203489279;
      10175: inst = 32'd136314880;
      10176: inst = 32'd268468224;
      10177: inst = 32'd201345488;
      10178: inst = 32'd203489279;
      10179: inst = 32'd136314880;
      10180: inst = 32'd268468224;
      10181: inst = 32'd201345489;
      10182: inst = 32'd203489279;
      10183: inst = 32'd136314880;
      10184: inst = 32'd268468224;
      10185: inst = 32'd201345490;
      10186: inst = 32'd203489279;
      10187: inst = 32'd136314880;
      10188: inst = 32'd268468224;
      10189: inst = 32'd201345491;
      10190: inst = 32'd203489279;
      10191: inst = 32'd136314880;
      10192: inst = 32'd268468224;
      10193: inst = 32'd201345492;
      10194: inst = 32'd203489279;
      10195: inst = 32'd136314880;
      10196: inst = 32'd268468224;
      10197: inst = 32'd201345493;
      10198: inst = 32'd203489279;
      10199: inst = 32'd136314880;
      10200: inst = 32'd268468224;
      10201: inst = 32'd201345494;
      10202: inst = 32'd203489279;
      10203: inst = 32'd136314880;
      10204: inst = 32'd268468224;
      10205: inst = 32'd201345495;
      10206: inst = 32'd203489279;
      10207: inst = 32'd136314880;
      10208: inst = 32'd268468224;
      10209: inst = 32'd201345496;
      10210: inst = 32'd203489279;
      10211: inst = 32'd136314880;
      10212: inst = 32'd268468224;
      10213: inst = 32'd201345497;
      10214: inst = 32'd203489279;
      10215: inst = 32'd136314880;
      10216: inst = 32'd268468224;
      10217: inst = 32'd201345498;
      10218: inst = 32'd203489279;
      10219: inst = 32'd136314880;
      10220: inst = 32'd268468224;
      10221: inst = 32'd201345499;
      10222: inst = 32'd203489279;
      10223: inst = 32'd136314880;
      10224: inst = 32'd268468224;
      10225: inst = 32'd201345500;
      10226: inst = 32'd203489279;
      10227: inst = 32'd136314880;
      10228: inst = 32'd268468224;
      10229: inst = 32'd201345501;
      10230: inst = 32'd203489279;
      10231: inst = 32'd136314880;
      10232: inst = 32'd268468224;
      10233: inst = 32'd201345502;
      10234: inst = 32'd203489279;
      10235: inst = 32'd136314880;
      10236: inst = 32'd268468224;
      10237: inst = 32'd201345503;
      10238: inst = 32'd203489279;
      10239: inst = 32'd136314880;
      10240: inst = 32'd268468224;
      10241: inst = 32'd201345504;
      10242: inst = 32'd203489279;
      10243: inst = 32'd136314880;
      10244: inst = 32'd268468224;
      10245: inst = 32'd201345505;
      10246: inst = 32'd203489279;
      10247: inst = 32'd136314880;
      10248: inst = 32'd268468224;
      10249: inst = 32'd201345506;
      10250: inst = 32'd203489247;
      10251: inst = 32'd136314880;
      10252: inst = 32'd268468224;
      10253: inst = 32'd201345507;
      10254: inst = 32'd203489279;
      10255: inst = 32'd136314880;
      10256: inst = 32'd268468224;
      10257: inst = 32'd201345508;
      10258: inst = 32'd203482840;
      10259: inst = 32'd136314880;
      10260: inst = 32'd268468224;
      10261: inst = 32'd201345509;
      10262: inst = 32'd203484886;
      10263: inst = 32'd136314880;
      10264: inst = 32'd268468224;
      10265: inst = 32'd201345510;
      10266: inst = 32'd203486901;
      10267: inst = 32'd136314880;
      10268: inst = 32'd268468224;
      10269: inst = 32'd201345511;
      10270: inst = 32'd203484854;
      10271: inst = 32'd136314880;
      10272: inst = 32'd268468224;
      10273: inst = 32'd201345512;
      10274: inst = 32'd203484886;
      10275: inst = 32'd136314880;
      10276: inst = 32'd268468224;
      10277: inst = 32'd201345513;
      10278: inst = 32'd203484854;
      10279: inst = 32'd136314880;
      10280: inst = 32'd268468224;
      10281: inst = 32'd201345514;
      10282: inst = 32'd203486870;
      10283: inst = 32'd136314880;
      10284: inst = 32'd268468224;
      10285: inst = 32'd201345515;
      10286: inst = 32'd203486870;
      10287: inst = 32'd136314880;
      10288: inst = 32'd268468224;
      10289: inst = 32'd201345516;
      10290: inst = 32'd203484887;
      10291: inst = 32'd136314880;
      10292: inst = 32'd268468224;
      10293: inst = 32'd201345517;
      10294: inst = 32'd203484886;
      10295: inst = 32'd136314880;
      10296: inst = 32'd268468224;
      10297: inst = 32'd201345518;
      10298: inst = 32'd203488883;
      10299: inst = 32'd136314880;
      10300: inst = 32'd268468224;
      10301: inst = 32'd201345519;
      10302: inst = 32'd203471621;
      10303: inst = 32'd136314880;
      10304: inst = 32'd268468224;
      10305: inst = 32'd201345520;
      10306: inst = 32'd203486115;
      10307: inst = 32'd136314880;
      10308: inst = 32'd268468224;
      10309: inst = 32'd201345521;
      10310: inst = 32'd203478024;
      10311: inst = 32'd136314880;
      10312: inst = 32'd268468224;
      10313: inst = 32'd201345522;
      10314: inst = 32'd203489275;
      10315: inst = 32'd136314880;
      10316: inst = 32'd268468224;
      10317: inst = 32'd201345523;
      10318: inst = 32'd203483036;
      10319: inst = 32'd136314880;
      10320: inst = 32'd268468224;
      10321: inst = 32'd201345524;
      10322: inst = 32'd203483004;
      10323: inst = 32'd136314880;
      10324: inst = 32'd268468224;
      10325: inst = 32'd201345525;
      10326: inst = 32'd203489049;
      10327: inst = 32'd136314880;
      10328: inst = 32'd268468224;
      10329: inst = 32'd201345526;
      10330: inst = 32'd203477960;
      10331: inst = 32'd136314880;
      10332: inst = 32'd268468224;
      10333: inst = 32'd201345527;
      10334: inst = 32'd203484102;
      10335: inst = 32'd136314880;
      10336: inst = 32'd268468224;
      10337: inst = 32'd201345528;
      10338: inst = 32'd203482052;
      10339: inst = 32'd136314880;
      10340: inst = 32'd268468224;
      10341: inst = 32'd201345529;
      10342: inst = 32'd203480036;
      10343: inst = 32'd136314880;
      10344: inst = 32'd268468224;
      10345: inst = 32'd201345530;
      10346: inst = 32'd203480004;
      10347: inst = 32'd136314880;
      10348: inst = 32'd268468224;
      10349: inst = 32'd201345531;
      10350: inst = 32'd203482052;
      10351: inst = 32'd136314880;
      10352: inst = 32'd268468224;
      10353: inst = 32'd201345532;
      10354: inst = 32'd203484036;
      10355: inst = 32'd136314880;
      10356: inst = 32'd268468224;
      10357: inst = 32'd201345533;
      10358: inst = 32'd203484069;
      10359: inst = 32'd136314880;
      10360: inst = 32'd268468224;
      10361: inst = 32'd201345534;
      10362: inst = 32'd203482021;
      10363: inst = 32'd136314880;
      10364: inst = 32'd268468224;
      10365: inst = 32'd201345535;
      10366: inst = 32'd203471619;
      10367: inst = 32'd136314880;
      10368: inst = 32'd268468224;
      10369: inst = 32'd201345536;
      10370: inst = 32'd203484854;
      10371: inst = 32'd136314880;
      10372: inst = 32'd268468224;
      10373: inst = 32'd201345537;
      10374: inst = 32'd203484854;
      10375: inst = 32'd136314880;
      10376: inst = 32'd268468224;
      10377: inst = 32'd201345538;
      10378: inst = 32'd203484854;
      10379: inst = 32'd136314880;
      10380: inst = 32'd268468224;
      10381: inst = 32'd201345539;
      10382: inst = 32'd203484853;
      10383: inst = 32'd136314880;
      10384: inst = 32'd268468224;
      10385: inst = 32'd201345540;
      10386: inst = 32'd203484885;
      10387: inst = 32'd136314880;
      10388: inst = 32'd268468224;
      10389: inst = 32'd201345541;
      10390: inst = 32'd203484886;
      10391: inst = 32'd136314880;
      10392: inst = 32'd268468224;
      10393: inst = 32'd201345542;
      10394: inst = 32'd203484886;
      10395: inst = 32'd136314880;
      10396: inst = 32'd268468224;
      10397: inst = 32'd201345543;
      10398: inst = 32'd203482839;
      10399: inst = 32'd136314880;
      10400: inst = 32'd268468224;
      10401: inst = 32'd201345544;
      10402: inst = 32'd203484889;
      10403: inst = 32'd136314880;
      10404: inst = 32'd268468224;
      10405: inst = 32'd201345545;
      10406: inst = 32'd203484889;
      10407: inst = 32'd136314880;
      10408: inst = 32'd268468224;
      10409: inst = 32'd201345546;
      10410: inst = 32'd203484922;
      10411: inst = 32'd136314880;
      10412: inst = 32'd268468224;
      10413: inst = 32'd201345547;
      10414: inst = 32'd203484922;
      10415: inst = 32'd136314880;
      10416: inst = 32'd268468224;
      10417: inst = 32'd201345548;
      10418: inst = 32'd203484921;
      10419: inst = 32'd136314880;
      10420: inst = 32'd268468224;
      10421: inst = 32'd201345549;
      10422: inst = 32'd203480727;
      10423: inst = 32'd136314880;
      10424: inst = 32'd268468224;
      10425: inst = 32'd201345550;
      10426: inst = 32'd203482807;
      10427: inst = 32'd136314880;
      10428: inst = 32'd268468224;
      10429: inst = 32'd201345551;
      10430: inst = 32'd203484985;
      10431: inst = 32'd136314880;
      10432: inst = 32'd268468224;
      10433: inst = 32'd201345552;
      10434: inst = 32'd203484854;
      10435: inst = 32'd136314880;
      10436: inst = 32'd268468224;
      10437: inst = 32'd201345553;
      10438: inst = 32'd203484854;
      10439: inst = 32'd136314880;
      10440: inst = 32'd268468224;
      10441: inst = 32'd201345554;
      10442: inst = 32'd203484854;
      10443: inst = 32'd136314880;
      10444: inst = 32'd268468224;
      10445: inst = 32'd201345555;
      10446: inst = 32'd203484854;
      10447: inst = 32'd136314880;
      10448: inst = 32'd268468224;
      10449: inst = 32'd201345556;
      10450: inst = 32'd203484854;
      10451: inst = 32'd136314880;
      10452: inst = 32'd268468224;
      10453: inst = 32'd201345557;
      10454: inst = 32'd203484854;
      10455: inst = 32'd136314880;
      10456: inst = 32'd268468224;
      10457: inst = 32'd201345558;
      10458: inst = 32'd203484854;
      10459: inst = 32'd136314880;
      10460: inst = 32'd268468224;
      10461: inst = 32'd201345559;
      10462: inst = 32'd203484854;
      10463: inst = 32'd136314880;
      10464: inst = 32'd268468224;
      10465: inst = 32'd201345560;
      10466: inst = 32'd203484854;
      10467: inst = 32'd136314880;
      10468: inst = 32'd268468224;
      10469: inst = 32'd201345561;
      10470: inst = 32'd203484854;
      10471: inst = 32'd136314880;
      10472: inst = 32'd268468224;
      10473: inst = 32'd201345562;
      10474: inst = 32'd203484855;
      10475: inst = 32'd136314880;
      10476: inst = 32'd268468224;
      10477: inst = 32'd201345563;
      10478: inst = 32'd203482808;
      10479: inst = 32'd136314880;
      10480: inst = 32'd268468224;
      10481: inst = 32'd201345564;
      10482: inst = 32'd203489278;
      10483: inst = 32'd136314880;
      10484: inst = 32'd268468224;
      10485: inst = 32'd201345565;
      10486: inst = 32'd203489279;
      10487: inst = 32'd136314880;
      10488: inst = 32'd268468224;
      10489: inst = 32'd201345566;
      10490: inst = 32'd203489279;
      10491: inst = 32'd136314880;
      10492: inst = 32'd268468224;
      10493: inst = 32'd201345567;
      10494: inst = 32'd203489279;
      10495: inst = 32'd136314880;
      10496: inst = 32'd268468224;
      10497: inst = 32'd201345568;
      10498: inst = 32'd203489279;
      10499: inst = 32'd136314880;
      10500: inst = 32'd268468224;
      10501: inst = 32'd201345569;
      10502: inst = 32'd203489279;
      10503: inst = 32'd136314880;
      10504: inst = 32'd268468224;
      10505: inst = 32'd201345570;
      10506: inst = 32'd203489279;
      10507: inst = 32'd136314880;
      10508: inst = 32'd268468224;
      10509: inst = 32'd201345571;
      10510: inst = 32'd203489279;
      10511: inst = 32'd136314880;
      10512: inst = 32'd268468224;
      10513: inst = 32'd201345572;
      10514: inst = 32'd203489279;
      10515: inst = 32'd136314880;
      10516: inst = 32'd268468224;
      10517: inst = 32'd201345573;
      10518: inst = 32'd203489279;
      10519: inst = 32'd136314880;
      10520: inst = 32'd268468224;
      10521: inst = 32'd201345574;
      10522: inst = 32'd203489279;
      10523: inst = 32'd136314880;
      10524: inst = 32'd268468224;
      10525: inst = 32'd201345575;
      10526: inst = 32'd203489279;
      10527: inst = 32'd136314880;
      10528: inst = 32'd268468224;
      10529: inst = 32'd201345576;
      10530: inst = 32'd203489279;
      10531: inst = 32'd136314880;
      10532: inst = 32'd268468224;
      10533: inst = 32'd201345577;
      10534: inst = 32'd203489279;
      10535: inst = 32'd136314880;
      10536: inst = 32'd268468224;
      10537: inst = 32'd201345578;
      10538: inst = 32'd203489279;
      10539: inst = 32'd136314880;
      10540: inst = 32'd268468224;
      10541: inst = 32'd201345579;
      10542: inst = 32'd203489279;
      10543: inst = 32'd136314880;
      10544: inst = 32'd268468224;
      10545: inst = 32'd201345580;
      10546: inst = 32'd203489279;
      10547: inst = 32'd136314880;
      10548: inst = 32'd268468224;
      10549: inst = 32'd201345581;
      10550: inst = 32'd203489279;
      10551: inst = 32'd136314880;
      10552: inst = 32'd268468224;
      10553: inst = 32'd201345582;
      10554: inst = 32'd203489279;
      10555: inst = 32'd136314880;
      10556: inst = 32'd268468224;
      10557: inst = 32'd201345583;
      10558: inst = 32'd203489279;
      10559: inst = 32'd136314880;
      10560: inst = 32'd268468224;
      10561: inst = 32'd201345584;
      10562: inst = 32'd203489279;
      10563: inst = 32'd136314880;
      10564: inst = 32'd268468224;
      10565: inst = 32'd201345585;
      10566: inst = 32'd203489279;
      10567: inst = 32'd136314880;
      10568: inst = 32'd268468224;
      10569: inst = 32'd201345586;
      10570: inst = 32'd203489279;
      10571: inst = 32'd136314880;
      10572: inst = 32'd268468224;
      10573: inst = 32'd201345587;
      10574: inst = 32'd203489279;
      10575: inst = 32'd136314880;
      10576: inst = 32'd268468224;
      10577: inst = 32'd201345588;
      10578: inst = 32'd203489279;
      10579: inst = 32'd136314880;
      10580: inst = 32'd268468224;
      10581: inst = 32'd201345589;
      10582: inst = 32'd203489279;
      10583: inst = 32'd136314880;
      10584: inst = 32'd268468224;
      10585: inst = 32'd201345590;
      10586: inst = 32'd203489279;
      10587: inst = 32'd136314880;
      10588: inst = 32'd268468224;
      10589: inst = 32'd201345591;
      10590: inst = 32'd203489279;
      10591: inst = 32'd136314880;
      10592: inst = 32'd268468224;
      10593: inst = 32'd201345592;
      10594: inst = 32'd203489279;
      10595: inst = 32'd136314880;
      10596: inst = 32'd268468224;
      10597: inst = 32'd201345593;
      10598: inst = 32'd203489279;
      10599: inst = 32'd136314880;
      10600: inst = 32'd268468224;
      10601: inst = 32'd201345594;
      10602: inst = 32'd203489279;
      10603: inst = 32'd136314880;
      10604: inst = 32'd268468224;
      10605: inst = 32'd201345595;
      10606: inst = 32'd203489279;
      10607: inst = 32'd136314880;
      10608: inst = 32'd268468224;
      10609: inst = 32'd201345596;
      10610: inst = 32'd203489279;
      10611: inst = 32'd136314880;
      10612: inst = 32'd268468224;
      10613: inst = 32'd201345597;
      10614: inst = 32'd203489279;
      10615: inst = 32'd136314880;
      10616: inst = 32'd268468224;
      10617: inst = 32'd201345598;
      10618: inst = 32'd203489279;
      10619: inst = 32'd136314880;
      10620: inst = 32'd268468224;
      10621: inst = 32'd201345599;
      10622: inst = 32'd203489279;
      10623: inst = 32'd136314880;
      10624: inst = 32'd268468224;
      10625: inst = 32'd201345600;
      10626: inst = 32'd203489279;
      10627: inst = 32'd136314880;
      10628: inst = 32'd268468224;
      10629: inst = 32'd201345601;
      10630: inst = 32'd203489279;
      10631: inst = 32'd136314880;
      10632: inst = 32'd268468224;
      10633: inst = 32'd201345602;
      10634: inst = 32'd203489247;
      10635: inst = 32'd136314880;
      10636: inst = 32'd268468224;
      10637: inst = 32'd201345603;
      10638: inst = 32'd203489279;
      10639: inst = 32'd136314880;
      10640: inst = 32'd268468224;
      10641: inst = 32'd201345604;
      10642: inst = 32'd203482840;
      10643: inst = 32'd136314880;
      10644: inst = 32'd268468224;
      10645: inst = 32'd201345605;
      10646: inst = 32'd203484886;
      10647: inst = 32'd136314880;
      10648: inst = 32'd268468224;
      10649: inst = 32'd201345606;
      10650: inst = 32'd203486901;
      10651: inst = 32'd136314880;
      10652: inst = 32'd268468224;
      10653: inst = 32'd201345607;
      10654: inst = 32'd203484854;
      10655: inst = 32'd136314880;
      10656: inst = 32'd268468224;
      10657: inst = 32'd201345608;
      10658: inst = 32'd203484886;
      10659: inst = 32'd136314880;
      10660: inst = 32'd268468224;
      10661: inst = 32'd201345609;
      10662: inst = 32'd203484854;
      10663: inst = 32'd136314880;
      10664: inst = 32'd268468224;
      10665: inst = 32'd201345610;
      10666: inst = 32'd203486902;
      10667: inst = 32'd136314880;
      10668: inst = 32'd268468224;
      10669: inst = 32'd201345611;
      10670: inst = 32'd203486870;
      10671: inst = 32'd136314880;
      10672: inst = 32'd268468224;
      10673: inst = 32'd201345612;
      10674: inst = 32'd203482839;
      10675: inst = 32'd136314880;
      10676: inst = 32'd268468224;
      10677: inst = 32'd201345613;
      10678: inst = 32'd203484886;
      10679: inst = 32'd136314880;
      10680: inst = 32'd268468224;
      10681: inst = 32'd201345614;
      10682: inst = 32'd203488915;
      10683: inst = 32'd136314880;
      10684: inst = 32'd268468224;
      10685: inst = 32'd201345615;
      10686: inst = 32'd203469573;
      10687: inst = 32'd136314880;
      10688: inst = 32'd268468224;
      10689: inst = 32'd201345616;
      10690: inst = 32'd203484002;
      10691: inst = 32'd136314880;
      10692: inst = 32'd268468224;
      10693: inst = 32'd201345617;
      10694: inst = 32'd203475911;
      10695: inst = 32'd136314880;
      10696: inst = 32'd268468224;
      10697: inst = 32'd201345618;
      10698: inst = 32'd203489211;
      10699: inst = 32'd136314880;
      10700: inst = 32'd268468224;
      10701: inst = 32'd201345619;
      10702: inst = 32'd203485053;
      10703: inst = 32'd136314880;
      10704: inst = 32'd268468224;
      10705: inst = 32'd201345620;
      10706: inst = 32'd203489181;
      10707: inst = 32'd136314880;
      10708: inst = 32'd268468224;
      10709: inst = 32'd201345621;
      10710: inst = 32'd203489016;
      10711: inst = 32'd136314880;
      10712: inst = 32'd268468224;
      10713: inst = 32'd201345622;
      10714: inst = 32'd203477960;
      10715: inst = 32'd136314880;
      10716: inst = 32'd268468224;
      10717: inst = 32'd201345623;
      10718: inst = 32'd203479972;
      10719: inst = 32'd136314880;
      10720: inst = 32'd268468224;
      10721: inst = 32'd201345624;
      10722: inst = 32'd203480004;
      10723: inst = 32'd136314880;
      10724: inst = 32'd268468224;
      10725: inst = 32'd201345625;
      10726: inst = 32'd203480036;
      10727: inst = 32'd136314880;
      10728: inst = 32'd268468224;
      10729: inst = 32'd201345626;
      10730: inst = 32'd203480004;
      10731: inst = 32'd136314880;
      10732: inst = 32'd268468224;
      10733: inst = 32'd201345627;
      10734: inst = 32'd203484068;
      10735: inst = 32'd136314880;
      10736: inst = 32'd268468224;
      10737: inst = 32'd201345628;
      10738: inst = 32'd203484036;
      10739: inst = 32'd136314880;
      10740: inst = 32'd268468224;
      10741: inst = 32'd201345629;
      10742: inst = 32'd203484068;
      10743: inst = 32'd136314880;
      10744: inst = 32'd268468224;
      10745: inst = 32'd201345630;
      10746: inst = 32'd203477957;
      10747: inst = 32'd136314880;
      10748: inst = 32'd268468224;
      10749: inst = 32'd201345631;
      10750: inst = 32'd203469635;
      10751: inst = 32'd136314880;
      10752: inst = 32'd268468224;
      10753: inst = 32'd201345632;
      10754: inst = 32'd203484854;
      10755: inst = 32'd136314880;
      10756: inst = 32'd268468224;
      10757: inst = 32'd201345633;
      10758: inst = 32'd203486902;
      10759: inst = 32'd136314880;
      10760: inst = 32'd268468224;
      10761: inst = 32'd201345634;
      10762: inst = 32'd203484854;
      10763: inst = 32'd136314880;
      10764: inst = 32'd268468224;
      10765: inst = 32'd201345635;
      10766: inst = 32'd203484854;
      10767: inst = 32'd136314880;
      10768: inst = 32'd268468224;
      10769: inst = 32'd201345636;
      10770: inst = 32'd203484886;
      10771: inst = 32'd136314880;
      10772: inst = 32'd268468224;
      10773: inst = 32'd201345637;
      10774: inst = 32'd203484886;
      10775: inst = 32'd136314880;
      10776: inst = 32'd268468224;
      10777: inst = 32'd201345638;
      10778: inst = 32'd203484887;
      10779: inst = 32'd136314880;
      10780: inst = 32'd268468224;
      10781: inst = 32'd201345639;
      10782: inst = 32'd203482840;
      10783: inst = 32'd136314880;
      10784: inst = 32'd268468224;
      10785: inst = 32'd201345640;
      10786: inst = 32'd203482841;
      10787: inst = 32'd136314880;
      10788: inst = 32'd268468224;
      10789: inst = 32'd201345641;
      10790: inst = 32'd203482810;
      10791: inst = 32'd136314880;
      10792: inst = 32'd268468224;
      10793: inst = 32'd201345642;
      10794: inst = 32'd203484923;
      10795: inst = 32'd136314880;
      10796: inst = 32'd268468224;
      10797: inst = 32'd201345643;
      10798: inst = 32'd203484923;
      10799: inst = 32'd136314880;
      10800: inst = 32'd268468224;
      10801: inst = 32'd201345644;
      10802: inst = 32'd203482874;
      10803: inst = 32'd136314880;
      10804: inst = 32'd268468224;
      10805: inst = 32'd201345645;
      10806: inst = 32'd203485019;
      10807: inst = 32'd136314880;
      10808: inst = 32'd268468224;
      10809: inst = 32'd201345646;
      10810: inst = 32'd203482873;
      10811: inst = 32'd136314880;
      10812: inst = 32'd268468224;
      10813: inst = 32'd201345647;
      10814: inst = 32'd203480760;
      10815: inst = 32'd136314880;
      10816: inst = 32'd268468224;
      10817: inst = 32'd201345648;
      10818: inst = 32'd203484854;
      10819: inst = 32'd136314880;
      10820: inst = 32'd268468224;
      10821: inst = 32'd201345649;
      10822: inst = 32'd203484854;
      10823: inst = 32'd136314880;
      10824: inst = 32'd268468224;
      10825: inst = 32'd201345650;
      10826: inst = 32'd203484854;
      10827: inst = 32'd136314880;
      10828: inst = 32'd268468224;
      10829: inst = 32'd201345651;
      10830: inst = 32'd203484854;
      10831: inst = 32'd136314880;
      10832: inst = 32'd268468224;
      10833: inst = 32'd201345652;
      10834: inst = 32'd203484854;
      10835: inst = 32'd136314880;
      10836: inst = 32'd268468224;
      10837: inst = 32'd201345653;
      10838: inst = 32'd203484854;
      10839: inst = 32'd136314880;
      10840: inst = 32'd268468224;
      10841: inst = 32'd201345654;
      10842: inst = 32'd203484854;
      10843: inst = 32'd136314880;
      10844: inst = 32'd268468224;
      10845: inst = 32'd201345655;
      10846: inst = 32'd203484854;
      10847: inst = 32'd136314880;
      10848: inst = 32'd268468224;
      10849: inst = 32'd201345656;
      10850: inst = 32'd203484854;
      10851: inst = 32'd136314880;
      10852: inst = 32'd268468224;
      10853: inst = 32'd201345657;
      10854: inst = 32'd203484854;
      10855: inst = 32'd136314880;
      10856: inst = 32'd268468224;
      10857: inst = 32'd201345658;
      10858: inst = 32'd203484855;
      10859: inst = 32'd136314880;
      10860: inst = 32'd268468224;
      10861: inst = 32'd201345659;
      10862: inst = 32'd203482808;
      10863: inst = 32'd136314880;
      10864: inst = 32'd268468224;
      10865: inst = 32'd201345660;
      10866: inst = 32'd203489278;
      10867: inst = 32'd136314880;
      10868: inst = 32'd268468224;
      10869: inst = 32'd201345661;
      10870: inst = 32'd203489279;
      10871: inst = 32'd136314880;
      10872: inst = 32'd268468224;
      10873: inst = 32'd201345662;
      10874: inst = 32'd203489279;
      10875: inst = 32'd136314880;
      10876: inst = 32'd268468224;
      10877: inst = 32'd201345663;
      10878: inst = 32'd203489279;
      10879: inst = 32'd136314880;
      10880: inst = 32'd268468224;
      10881: inst = 32'd201345664;
      10882: inst = 32'd203489279;
      10883: inst = 32'd136314880;
      10884: inst = 32'd268468224;
      10885: inst = 32'd201345665;
      10886: inst = 32'd203489279;
      10887: inst = 32'd136314880;
      10888: inst = 32'd268468224;
      10889: inst = 32'd201345666;
      10890: inst = 32'd203489279;
      10891: inst = 32'd136314880;
      10892: inst = 32'd268468224;
      10893: inst = 32'd201345667;
      10894: inst = 32'd203489279;
      10895: inst = 32'd136314880;
      10896: inst = 32'd268468224;
      10897: inst = 32'd201345668;
      10898: inst = 32'd203489279;
      10899: inst = 32'd136314880;
      10900: inst = 32'd268468224;
      10901: inst = 32'd201345669;
      10902: inst = 32'd203489279;
      10903: inst = 32'd136314880;
      10904: inst = 32'd268468224;
      10905: inst = 32'd201345670;
      10906: inst = 32'd203489279;
      10907: inst = 32'd136314880;
      10908: inst = 32'd268468224;
      10909: inst = 32'd201345671;
      10910: inst = 32'd203489279;
      10911: inst = 32'd136314880;
      10912: inst = 32'd268468224;
      10913: inst = 32'd201345672;
      10914: inst = 32'd203489279;
      10915: inst = 32'd136314880;
      10916: inst = 32'd268468224;
      10917: inst = 32'd201345673;
      10918: inst = 32'd203489279;
      10919: inst = 32'd136314880;
      10920: inst = 32'd268468224;
      10921: inst = 32'd201345674;
      10922: inst = 32'd203489279;
      10923: inst = 32'd136314880;
      10924: inst = 32'd268468224;
      10925: inst = 32'd201345675;
      10926: inst = 32'd203489279;
      10927: inst = 32'd136314880;
      10928: inst = 32'd268468224;
      10929: inst = 32'd201345676;
      10930: inst = 32'd203489279;
      10931: inst = 32'd136314880;
      10932: inst = 32'd268468224;
      10933: inst = 32'd201345677;
      10934: inst = 32'd203489279;
      10935: inst = 32'd136314880;
      10936: inst = 32'd268468224;
      10937: inst = 32'd201345678;
      10938: inst = 32'd203489279;
      10939: inst = 32'd136314880;
      10940: inst = 32'd268468224;
      10941: inst = 32'd201345679;
      10942: inst = 32'd203489279;
      10943: inst = 32'd136314880;
      10944: inst = 32'd268468224;
      10945: inst = 32'd201345680;
      10946: inst = 32'd203489279;
      10947: inst = 32'd136314880;
      10948: inst = 32'd268468224;
      10949: inst = 32'd201345681;
      10950: inst = 32'd203489279;
      10951: inst = 32'd136314880;
      10952: inst = 32'd268468224;
      10953: inst = 32'd201345682;
      10954: inst = 32'd203489279;
      10955: inst = 32'd136314880;
      10956: inst = 32'd268468224;
      10957: inst = 32'd201345683;
      10958: inst = 32'd203489279;
      10959: inst = 32'd136314880;
      10960: inst = 32'd268468224;
      10961: inst = 32'd201345684;
      10962: inst = 32'd203489279;
      10963: inst = 32'd136314880;
      10964: inst = 32'd268468224;
      10965: inst = 32'd201345685;
      10966: inst = 32'd203489279;
      10967: inst = 32'd136314880;
      10968: inst = 32'd268468224;
      10969: inst = 32'd201345686;
      10970: inst = 32'd203489279;
      10971: inst = 32'd136314880;
      10972: inst = 32'd268468224;
      10973: inst = 32'd201345687;
      10974: inst = 32'd203489279;
      10975: inst = 32'd136314880;
      10976: inst = 32'd268468224;
      10977: inst = 32'd201345688;
      10978: inst = 32'd203489279;
      10979: inst = 32'd136314880;
      10980: inst = 32'd268468224;
      10981: inst = 32'd201345689;
      10982: inst = 32'd203489279;
      10983: inst = 32'd136314880;
      10984: inst = 32'd268468224;
      10985: inst = 32'd201345690;
      10986: inst = 32'd203489279;
      10987: inst = 32'd136314880;
      10988: inst = 32'd268468224;
      10989: inst = 32'd201345691;
      10990: inst = 32'd203489279;
      10991: inst = 32'd136314880;
      10992: inst = 32'd268468224;
      10993: inst = 32'd201345692;
      10994: inst = 32'd203489279;
      10995: inst = 32'd136314880;
      10996: inst = 32'd268468224;
      10997: inst = 32'd201345693;
      10998: inst = 32'd203489279;
      10999: inst = 32'd136314880;
      11000: inst = 32'd268468224;
      11001: inst = 32'd201345694;
      11002: inst = 32'd203489279;
      11003: inst = 32'd136314880;
      11004: inst = 32'd268468224;
      11005: inst = 32'd201345695;
      11006: inst = 32'd203489279;
      11007: inst = 32'd136314880;
      11008: inst = 32'd268468224;
      11009: inst = 32'd201345696;
      11010: inst = 32'd203489278;
      11011: inst = 32'd136314880;
      11012: inst = 32'd268468224;
      11013: inst = 32'd201345697;
      11014: inst = 32'd203489279;
      11015: inst = 32'd136314880;
      11016: inst = 32'd268468224;
      11017: inst = 32'd201345698;
      11018: inst = 32'd203489247;
      11019: inst = 32'd136314880;
      11020: inst = 32'd268468224;
      11021: inst = 32'd201345699;
      11022: inst = 32'd203489279;
      11023: inst = 32'd136314880;
      11024: inst = 32'd268468224;
      11025: inst = 32'd201345700;
      11026: inst = 32'd203482840;
      11027: inst = 32'd136314880;
      11028: inst = 32'd268468224;
      11029: inst = 32'd201345701;
      11030: inst = 32'd203484886;
      11031: inst = 32'd136314880;
      11032: inst = 32'd268468224;
      11033: inst = 32'd201345702;
      11034: inst = 32'd203484853;
      11035: inst = 32'd136314880;
      11036: inst = 32'd268468224;
      11037: inst = 32'd201345703;
      11038: inst = 32'd203484854;
      11039: inst = 32'd136314880;
      11040: inst = 32'd268468224;
      11041: inst = 32'd201345704;
      11042: inst = 32'd203484887;
      11043: inst = 32'd136314880;
      11044: inst = 32'd268468224;
      11045: inst = 32'd201345705;
      11046: inst = 32'd203484854;
      11047: inst = 32'd136314880;
      11048: inst = 32'd268468224;
      11049: inst = 32'd201345706;
      11050: inst = 32'd203486902;
      11051: inst = 32'd136314880;
      11052: inst = 32'd268468224;
      11053: inst = 32'd201345707;
      11054: inst = 32'd203484822;
      11055: inst = 32'd136314880;
      11056: inst = 32'd268468224;
      11057: inst = 32'd201345708;
      11058: inst = 32'd203482839;
      11059: inst = 32'd136314880;
      11060: inst = 32'd268468224;
      11061: inst = 32'd201345709;
      11062: inst = 32'd203484886;
      11063: inst = 32'd136314880;
      11064: inst = 32'd268468224;
      11065: inst = 32'd201345710;
      11066: inst = 32'd203488915;
      11067: inst = 32'd136314880;
      11068: inst = 32'd268468224;
      11069: inst = 32'd201345711;
      11070: inst = 32'd203469573;
      11071: inst = 32'd136314880;
      11072: inst = 32'd268468224;
      11073: inst = 32'd201345712;
      11074: inst = 32'd203484068;
      11075: inst = 32'd136314880;
      11076: inst = 32'd268468224;
      11077: inst = 32'd201345713;
      11078: inst = 32'd203475977;
      11079: inst = 32'd136314880;
      11080: inst = 32'd268468224;
      11081: inst = 32'd201345714;
      11082: inst = 32'd203489113;
      11083: inst = 32'd136314880;
      11084: inst = 32'd268468224;
      11085: inst = 32'd201345715;
      11086: inst = 32'd203483070;
      11087: inst = 32'd136314880;
      11088: inst = 32'd268468224;
      11089: inst = 32'd201345716;
      11090: inst = 32'd203487231;
      11091: inst = 32'd136314880;
      11092: inst = 32'd268468224;
      11093: inst = 32'd201345717;
      11094: inst = 32'd203489016;
      11095: inst = 32'd136314880;
      11096: inst = 32'd268468224;
      11097: inst = 32'd201345718;
      11098: inst = 32'd203478090;
      11099: inst = 32'd136314880;
      11100: inst = 32'd268468224;
      11101: inst = 32'd201345719;
      11102: inst = 32'd203479974;
      11103: inst = 32'd136314880;
      11104: inst = 32'd268468224;
      11105: inst = 32'd201345720;
      11106: inst = 32'd203480006;
      11107: inst = 32'd136314880;
      11108: inst = 32'd268468224;
      11109: inst = 32'd201345721;
      11110: inst = 32'd203480038;
      11111: inst = 32'd136314880;
      11112: inst = 32'd268468224;
      11113: inst = 32'd201345722;
      11114: inst = 32'd203477958;
      11115: inst = 32'd136314880;
      11116: inst = 32'd268468224;
      11117: inst = 32'd201345723;
      11118: inst = 32'd203480005;
      11119: inst = 32'd136314880;
      11120: inst = 32'd268468224;
      11121: inst = 32'd201345724;
      11122: inst = 32'd203482021;
      11123: inst = 32'd136314880;
      11124: inst = 32'd268468224;
      11125: inst = 32'd201345725;
      11126: inst = 32'd203482053;
      11127: inst = 32'd136314880;
      11128: inst = 32'd268468224;
      11129: inst = 32'd201345726;
      11130: inst = 32'd203479974;
      11131: inst = 32'd136314880;
      11132: inst = 32'd268468224;
      11133: inst = 32'd201345727;
      11134: inst = 32'd203471621;
      11135: inst = 32'd136314880;
      11136: inst = 32'd268468224;
      11137: inst = 32'd201345728;
      11138: inst = 32'd203486871;
      11139: inst = 32'd136314880;
      11140: inst = 32'd268468224;
      11141: inst = 32'd201345729;
      11142: inst = 32'd203486903;
      11143: inst = 32'd136314880;
      11144: inst = 32'd268468224;
      11145: inst = 32'd201345730;
      11146: inst = 32'd203486902;
      11147: inst = 32'd136314880;
      11148: inst = 32'd268468224;
      11149: inst = 32'd201345731;
      11150: inst = 32'd203484854;
      11151: inst = 32'd136314880;
      11152: inst = 32'd268468224;
      11153: inst = 32'd201345732;
      11154: inst = 32'd203484854;
      11155: inst = 32'd136314880;
      11156: inst = 32'd268468224;
      11157: inst = 32'd201345733;
      11158: inst = 32'd203482806;
      11159: inst = 32'd136314880;
      11160: inst = 32'd268468224;
      11161: inst = 32'd201345734;
      11162: inst = 32'd203484887;
      11163: inst = 32'd136314880;
      11164: inst = 32'd268468224;
      11165: inst = 32'd201345735;
      11166: inst = 32'd203482873;
      11167: inst = 32'd136314880;
      11168: inst = 32'd268468224;
      11169: inst = 32'd201345736;
      11170: inst = 32'd203484955;
      11171: inst = 32'd136314880;
      11172: inst = 32'd268468224;
      11173: inst = 32'd201345737;
      11174: inst = 32'd203480763;
      11175: inst = 32'd136314880;
      11176: inst = 32'd268468224;
      11177: inst = 32'd201345738;
      11178: inst = 32'd203480795;
      11179: inst = 32'd136314880;
      11180: inst = 32'd268468224;
      11181: inst = 32'd201345739;
      11182: inst = 32'd203482876;
      11183: inst = 32'd136314880;
      11184: inst = 32'd268468224;
      11185: inst = 32'd201345740;
      11186: inst = 32'd203480795;
      11187: inst = 32'd136314880;
      11188: inst = 32'd268468224;
      11189: inst = 32'd201345741;
      11190: inst = 32'd203480794;
      11191: inst = 32'd136314880;
      11192: inst = 32'd268468224;
      11193: inst = 32'd201345742;
      11194: inst = 32'd203485019;
      11195: inst = 32'd136314880;
      11196: inst = 32'd268468224;
      11197: inst = 32'd201345743;
      11198: inst = 32'd203480825;
      11199: inst = 32'd136314880;
      11200: inst = 32'd268468224;
      11201: inst = 32'd201345744;
      11202: inst = 32'd203484854;
      11203: inst = 32'd136314880;
      11204: inst = 32'd268468224;
      11205: inst = 32'd201345745;
      11206: inst = 32'd203484854;
      11207: inst = 32'd136314880;
      11208: inst = 32'd268468224;
      11209: inst = 32'd201345746;
      11210: inst = 32'd203484854;
      11211: inst = 32'd136314880;
      11212: inst = 32'd268468224;
      11213: inst = 32'd201345747;
      11214: inst = 32'd203484854;
      11215: inst = 32'd136314880;
      11216: inst = 32'd268468224;
      11217: inst = 32'd201345748;
      11218: inst = 32'd203484854;
      11219: inst = 32'd136314880;
      11220: inst = 32'd268468224;
      11221: inst = 32'd201345749;
      11222: inst = 32'd203484854;
      11223: inst = 32'd136314880;
      11224: inst = 32'd268468224;
      11225: inst = 32'd201345750;
      11226: inst = 32'd203484854;
      11227: inst = 32'd136314880;
      11228: inst = 32'd268468224;
      11229: inst = 32'd201345751;
      11230: inst = 32'd203484854;
      11231: inst = 32'd136314880;
      11232: inst = 32'd268468224;
      11233: inst = 32'd201345752;
      11234: inst = 32'd203484854;
      11235: inst = 32'd136314880;
      11236: inst = 32'd268468224;
      11237: inst = 32'd201345753;
      11238: inst = 32'd203484854;
      11239: inst = 32'd136314880;
      11240: inst = 32'd268468224;
      11241: inst = 32'd201345754;
      11242: inst = 32'd203484855;
      11243: inst = 32'd136314880;
      11244: inst = 32'd268468224;
      11245: inst = 32'd201345755;
      11246: inst = 32'd203482808;
      11247: inst = 32'd136314880;
      11248: inst = 32'd268468224;
      11249: inst = 32'd201345756;
      11250: inst = 32'd203489278;
      11251: inst = 32'd136314880;
      11252: inst = 32'd268468224;
      11253: inst = 32'd201345757;
      11254: inst = 32'd203489279;
      11255: inst = 32'd136314880;
      11256: inst = 32'd268468224;
      11257: inst = 32'd201345758;
      11258: inst = 32'd203489279;
      11259: inst = 32'd136314880;
      11260: inst = 32'd268468224;
      11261: inst = 32'd201345759;
      11262: inst = 32'd203489279;
      11263: inst = 32'd136314880;
      11264: inst = 32'd268468224;
      11265: inst = 32'd201345760;
      11266: inst = 32'd203489279;
      11267: inst = 32'd136314880;
      11268: inst = 32'd268468224;
      11269: inst = 32'd201345761;
      11270: inst = 32'd203489279;
      11271: inst = 32'd136314880;
      11272: inst = 32'd268468224;
      11273: inst = 32'd201345762;
      11274: inst = 32'd203489279;
      11275: inst = 32'd136314880;
      11276: inst = 32'd268468224;
      11277: inst = 32'd201345763;
      11278: inst = 32'd203489279;
      11279: inst = 32'd136314880;
      11280: inst = 32'd268468224;
      11281: inst = 32'd201345764;
      11282: inst = 32'd203489279;
      11283: inst = 32'd136314880;
      11284: inst = 32'd268468224;
      11285: inst = 32'd201345765;
      11286: inst = 32'd203489279;
      11287: inst = 32'd136314880;
      11288: inst = 32'd268468224;
      11289: inst = 32'd201345766;
      11290: inst = 32'd203489279;
      11291: inst = 32'd136314880;
      11292: inst = 32'd268468224;
      11293: inst = 32'd201345767;
      11294: inst = 32'd203489279;
      11295: inst = 32'd136314880;
      11296: inst = 32'd268468224;
      11297: inst = 32'd201345768;
      11298: inst = 32'd203489279;
      11299: inst = 32'd136314880;
      11300: inst = 32'd268468224;
      11301: inst = 32'd201345769;
      11302: inst = 32'd203489279;
      11303: inst = 32'd136314880;
      11304: inst = 32'd268468224;
      11305: inst = 32'd201345770;
      11306: inst = 32'd203489279;
      11307: inst = 32'd136314880;
      11308: inst = 32'd268468224;
      11309: inst = 32'd201345771;
      11310: inst = 32'd203489279;
      11311: inst = 32'd136314880;
      11312: inst = 32'd268468224;
      11313: inst = 32'd201345772;
      11314: inst = 32'd203489279;
      11315: inst = 32'd136314880;
      11316: inst = 32'd268468224;
      11317: inst = 32'd201345773;
      11318: inst = 32'd203489279;
      11319: inst = 32'd136314880;
      11320: inst = 32'd268468224;
      11321: inst = 32'd201345774;
      11322: inst = 32'd203489279;
      11323: inst = 32'd136314880;
      11324: inst = 32'd268468224;
      11325: inst = 32'd201345775;
      11326: inst = 32'd203489279;
      11327: inst = 32'd136314880;
      11328: inst = 32'd268468224;
      11329: inst = 32'd201345776;
      11330: inst = 32'd203489279;
      11331: inst = 32'd136314880;
      11332: inst = 32'd268468224;
      11333: inst = 32'd201345777;
      11334: inst = 32'd203489279;
      11335: inst = 32'd136314880;
      11336: inst = 32'd268468224;
      11337: inst = 32'd201345778;
      11338: inst = 32'd203489279;
      11339: inst = 32'd136314880;
      11340: inst = 32'd268468224;
      11341: inst = 32'd201345779;
      11342: inst = 32'd203489279;
      11343: inst = 32'd136314880;
      11344: inst = 32'd268468224;
      11345: inst = 32'd201345780;
      11346: inst = 32'd203489279;
      11347: inst = 32'd136314880;
      11348: inst = 32'd268468224;
      11349: inst = 32'd201345781;
      11350: inst = 32'd203489279;
      11351: inst = 32'd136314880;
      11352: inst = 32'd268468224;
      11353: inst = 32'd201345782;
      11354: inst = 32'd203489279;
      11355: inst = 32'd136314880;
      11356: inst = 32'd268468224;
      11357: inst = 32'd201345783;
      11358: inst = 32'd203489279;
      11359: inst = 32'd136314880;
      11360: inst = 32'd268468224;
      11361: inst = 32'd201345784;
      11362: inst = 32'd203489279;
      11363: inst = 32'd136314880;
      11364: inst = 32'd268468224;
      11365: inst = 32'd201345785;
      11366: inst = 32'd203489279;
      11367: inst = 32'd136314880;
      11368: inst = 32'd268468224;
      11369: inst = 32'd201345786;
      11370: inst = 32'd203489279;
      11371: inst = 32'd136314880;
      11372: inst = 32'd268468224;
      11373: inst = 32'd201345787;
      11374: inst = 32'd203489279;
      11375: inst = 32'd136314880;
      11376: inst = 32'd268468224;
      11377: inst = 32'd201345788;
      11378: inst = 32'd203489279;
      11379: inst = 32'd136314880;
      11380: inst = 32'd268468224;
      11381: inst = 32'd201345789;
      11382: inst = 32'd203489279;
      11383: inst = 32'd136314880;
      11384: inst = 32'd268468224;
      11385: inst = 32'd201345790;
      11386: inst = 32'd203489279;
      11387: inst = 32'd136314880;
      11388: inst = 32'd268468224;
      11389: inst = 32'd201345791;
      11390: inst = 32'd203489279;
      11391: inst = 32'd136314880;
      11392: inst = 32'd268468224;
      11393: inst = 32'd201345792;
      11394: inst = 32'd203489278;
      11395: inst = 32'd136314880;
      11396: inst = 32'd268468224;
      11397: inst = 32'd201345793;
      11398: inst = 32'd203489279;
      11399: inst = 32'd136314880;
      11400: inst = 32'd268468224;
      11401: inst = 32'd201345794;
      11402: inst = 32'd203489247;
      11403: inst = 32'd136314880;
      11404: inst = 32'd268468224;
      11405: inst = 32'd201345795;
      11406: inst = 32'd203489279;
      11407: inst = 32'd136314880;
      11408: inst = 32'd268468224;
      11409: inst = 32'd201345796;
      11410: inst = 32'd203482840;
      11411: inst = 32'd136314880;
      11412: inst = 32'd268468224;
      11413: inst = 32'd201345797;
      11414: inst = 32'd203484886;
      11415: inst = 32'd136314880;
      11416: inst = 32'd268468224;
      11417: inst = 32'd201345798;
      11418: inst = 32'd203484853;
      11419: inst = 32'd136314880;
      11420: inst = 32'd268468224;
      11421: inst = 32'd201345799;
      11422: inst = 32'd203484854;
      11423: inst = 32'd136314880;
      11424: inst = 32'd268468224;
      11425: inst = 32'd201345800;
      11426: inst = 32'd203484887;
      11427: inst = 32'd136314880;
      11428: inst = 32'd268468224;
      11429: inst = 32'd201345801;
      11430: inst = 32'd203484854;
      11431: inst = 32'd136314880;
      11432: inst = 32'd268468224;
      11433: inst = 32'd201345802;
      11434: inst = 32'd203486902;
      11435: inst = 32'd136314880;
      11436: inst = 32'd268468224;
      11437: inst = 32'd201345803;
      11438: inst = 32'd203484822;
      11439: inst = 32'd136314880;
      11440: inst = 32'd268468224;
      11441: inst = 32'd201345804;
      11442: inst = 32'd203482839;
      11443: inst = 32'd136314880;
      11444: inst = 32'd268468224;
      11445: inst = 32'd201345805;
      11446: inst = 32'd203482838;
      11447: inst = 32'd136314880;
      11448: inst = 32'd268468224;
      11449: inst = 32'd201345806;
      11450: inst = 32'd203488915;
      11451: inst = 32'd136314880;
      11452: inst = 32'd268468224;
      11453: inst = 32'd201345807;
      11454: inst = 32'd203469573;
      11455: inst = 32'd136314880;
      11456: inst = 32'd268468224;
      11457: inst = 32'd201345808;
      11458: inst = 32'd203482053;
      11459: inst = 32'd136314880;
      11460: inst = 32'd268468224;
      11461: inst = 32'd201345809;
      11462: inst = 32'd203469735;
      11463: inst = 32'd136314880;
      11464: inst = 32'd268468224;
      11465: inst = 32'd201345810;
      11466: inst = 32'd203487098;
      11467: inst = 32'd136314880;
      11468: inst = 32'd268468224;
      11469: inst = 32'd201345811;
      11470: inst = 32'd203481021;
      11471: inst = 32'd136314880;
      11472: inst = 32'd268468224;
      11473: inst = 32'd201345812;
      11474: inst = 32'd203487230;
      11475: inst = 32'd136314880;
      11476: inst = 32'd268468224;
      11477: inst = 32'd201345813;
      11478: inst = 32'd203489145;
      11479: inst = 32'd136314880;
      11480: inst = 32'd268468224;
      11481: inst = 32'd201345814;
      11482: inst = 32'd203473897;
      11483: inst = 32'd136314880;
      11484: inst = 32'd268468224;
      11485: inst = 32'd201345815;
      11486: inst = 32'd203479943;
      11487: inst = 32'd136314880;
      11488: inst = 32'd268468224;
      11489: inst = 32'd201345816;
      11490: inst = 32'd203482023;
      11491: inst = 32'd136314880;
      11492: inst = 32'd268468224;
      11493: inst = 32'd201345817;
      11494: inst = 32'd203480007;
      11495: inst = 32'd136314880;
      11496: inst = 32'd268468224;
      11497: inst = 32'd201345818;
      11498: inst = 32'd203477959;
      11499: inst = 32'd136314880;
      11500: inst = 32'd268468224;
      11501: inst = 32'd201345819;
      11502: inst = 32'd203477990;
      11503: inst = 32'd136314880;
      11504: inst = 32'd268468224;
      11505: inst = 32'd201345820;
      11506: inst = 32'd203477957;
      11507: inst = 32'd136314880;
      11508: inst = 32'd268468224;
      11509: inst = 32'd201345821;
      11510: inst = 32'd203480006;
      11511: inst = 32'd136314880;
      11512: inst = 32'd268468224;
      11513: inst = 32'd201345822;
      11514: inst = 32'd203479943;
      11515: inst = 32'd136314880;
      11516: inst = 32'd268468224;
      11517: inst = 32'd201345823;
      11518: inst = 32'd203473606;
      11519: inst = 32'd136314880;
      11520: inst = 32'd268468224;
      11521: inst = 32'd201345824;
      11522: inst = 32'd203486871;
      11523: inst = 32'd136314880;
      11524: inst = 32'd268468224;
      11525: inst = 32'd201345825;
      11526: inst = 32'd203486903;
      11527: inst = 32'd136314880;
      11528: inst = 32'd268468224;
      11529: inst = 32'd201345826;
      11530: inst = 32'd203486903;
      11531: inst = 32'd136314880;
      11532: inst = 32'd268468224;
      11533: inst = 32'd201345827;
      11534: inst = 32'd203484854;
      11535: inst = 32'd136314880;
      11536: inst = 32'd268468224;
      11537: inst = 32'd201345828;
      11538: inst = 32'd203484854;
      11539: inst = 32'd136314880;
      11540: inst = 32'd268468224;
      11541: inst = 32'd201345829;
      11542: inst = 32'd203482807;
      11543: inst = 32'd136314880;
      11544: inst = 32'd268468224;
      11545: inst = 32'd201345830;
      11546: inst = 32'd203482840;
      11547: inst = 32'd136314880;
      11548: inst = 32'd268468224;
      11549: inst = 32'd201345831;
      11550: inst = 32'd203482874;
      11551: inst = 32'd136314880;
      11552: inst = 32'd268468224;
      11553: inst = 32'd201345832;
      11554: inst = 32'd203442728;
      11555: inst = 32'd136314880;
      11556: inst = 32'd268468224;
      11557: inst = 32'd201345833;
      11558: inst = 32'd203444875;
      11559: inst = 32'd136314880;
      11560: inst = 32'd268468224;
      11561: inst = 32'd201345834;
      11562: inst = 32'd203482909;
      11563: inst = 32'd136314880;
      11564: inst = 32'd268468224;
      11565: inst = 32'd201345835;
      11566: inst = 32'd203444843;
      11567: inst = 32'd136314880;
      11568: inst = 32'd268468224;
      11569: inst = 32'd201345836;
      11570: inst = 32'd203442794;
      11571: inst = 32'd136314880;
      11572: inst = 32'd268468224;
      11573: inst = 32'd201345837;
      11574: inst = 32'd203482940;
      11575: inst = 32'd136314880;
      11576: inst = 32'd268468224;
      11577: inst = 32'd201345838;
      11578: inst = 32'd203478714;
      11579: inst = 32'd136314880;
      11580: inst = 32'd268468224;
      11581: inst = 32'd201345839;
      11582: inst = 32'd203482939;
      11583: inst = 32'd136314880;
      11584: inst = 32'd268468224;
      11585: inst = 32'd201345840;
      11586: inst = 32'd203484854;
      11587: inst = 32'd136314880;
      11588: inst = 32'd268468224;
      11589: inst = 32'd201345841;
      11590: inst = 32'd203484854;
      11591: inst = 32'd136314880;
      11592: inst = 32'd268468224;
      11593: inst = 32'd201345842;
      11594: inst = 32'd203484854;
      11595: inst = 32'd136314880;
      11596: inst = 32'd268468224;
      11597: inst = 32'd201345843;
      11598: inst = 32'd203484854;
      11599: inst = 32'd136314880;
      11600: inst = 32'd268468224;
      11601: inst = 32'd201345844;
      11602: inst = 32'd203484854;
      11603: inst = 32'd136314880;
      11604: inst = 32'd268468224;
      11605: inst = 32'd201345845;
      11606: inst = 32'd203484854;
      11607: inst = 32'd136314880;
      11608: inst = 32'd268468224;
      11609: inst = 32'd201345846;
      11610: inst = 32'd203484854;
      11611: inst = 32'd136314880;
      11612: inst = 32'd268468224;
      11613: inst = 32'd201345847;
      11614: inst = 32'd203484854;
      11615: inst = 32'd136314880;
      11616: inst = 32'd268468224;
      11617: inst = 32'd201345848;
      11618: inst = 32'd203484854;
      11619: inst = 32'd136314880;
      11620: inst = 32'd268468224;
      11621: inst = 32'd201345849;
      11622: inst = 32'd203484854;
      11623: inst = 32'd136314880;
      11624: inst = 32'd268468224;
      11625: inst = 32'd201345850;
      11626: inst = 32'd203484855;
      11627: inst = 32'd136314880;
      11628: inst = 32'd268468224;
      11629: inst = 32'd201345851;
      11630: inst = 32'd203482808;
      11631: inst = 32'd136314880;
      11632: inst = 32'd268468224;
      11633: inst = 32'd201345852;
      11634: inst = 32'd203489278;
      11635: inst = 32'd136314880;
      11636: inst = 32'd268468224;
      11637: inst = 32'd201345853;
      11638: inst = 32'd203489279;
      11639: inst = 32'd136314880;
      11640: inst = 32'd268468224;
      11641: inst = 32'd201345854;
      11642: inst = 32'd203489279;
      11643: inst = 32'd136314880;
      11644: inst = 32'd268468224;
      11645: inst = 32'd201345855;
      11646: inst = 32'd203489279;
      11647: inst = 32'd136314880;
      11648: inst = 32'd268468224;
      11649: inst = 32'd201345856;
      11650: inst = 32'd203489279;
      11651: inst = 32'd136314880;
      11652: inst = 32'd268468224;
      11653: inst = 32'd201345857;
      11654: inst = 32'd203489279;
      11655: inst = 32'd136314880;
      11656: inst = 32'd268468224;
      11657: inst = 32'd201345858;
      11658: inst = 32'd203489279;
      11659: inst = 32'd136314880;
      11660: inst = 32'd268468224;
      11661: inst = 32'd201345859;
      11662: inst = 32'd203489279;
      11663: inst = 32'd136314880;
      11664: inst = 32'd268468224;
      11665: inst = 32'd201345860;
      11666: inst = 32'd203489279;
      11667: inst = 32'd136314880;
      11668: inst = 32'd268468224;
      11669: inst = 32'd201345861;
      11670: inst = 32'd203489279;
      11671: inst = 32'd136314880;
      11672: inst = 32'd268468224;
      11673: inst = 32'd201345862;
      11674: inst = 32'd203489279;
      11675: inst = 32'd136314880;
      11676: inst = 32'd268468224;
      11677: inst = 32'd201345863;
      11678: inst = 32'd203489279;
      11679: inst = 32'd136314880;
      11680: inst = 32'd268468224;
      11681: inst = 32'd201345864;
      11682: inst = 32'd203489279;
      11683: inst = 32'd136314880;
      11684: inst = 32'd268468224;
      11685: inst = 32'd201345865;
      11686: inst = 32'd203489279;
      11687: inst = 32'd136314880;
      11688: inst = 32'd268468224;
      11689: inst = 32'd201345866;
      11690: inst = 32'd203489279;
      11691: inst = 32'd136314880;
      11692: inst = 32'd268468224;
      11693: inst = 32'd201345867;
      11694: inst = 32'd203489279;
      11695: inst = 32'd136314880;
      11696: inst = 32'd268468224;
      11697: inst = 32'd201345868;
      11698: inst = 32'd203489279;
      11699: inst = 32'd136314880;
      11700: inst = 32'd268468224;
      11701: inst = 32'd201345869;
      11702: inst = 32'd203489279;
      11703: inst = 32'd136314880;
      11704: inst = 32'd268468224;
      11705: inst = 32'd201345870;
      11706: inst = 32'd203489279;
      11707: inst = 32'd136314880;
      11708: inst = 32'd268468224;
      11709: inst = 32'd201345871;
      11710: inst = 32'd203489279;
      11711: inst = 32'd136314880;
      11712: inst = 32'd268468224;
      11713: inst = 32'd201345872;
      11714: inst = 32'd203489279;
      11715: inst = 32'd136314880;
      11716: inst = 32'd268468224;
      11717: inst = 32'd201345873;
      11718: inst = 32'd203489279;
      11719: inst = 32'd136314880;
      11720: inst = 32'd268468224;
      11721: inst = 32'd201345874;
      11722: inst = 32'd203489279;
      11723: inst = 32'd136314880;
      11724: inst = 32'd268468224;
      11725: inst = 32'd201345875;
      11726: inst = 32'd203489279;
      11727: inst = 32'd136314880;
      11728: inst = 32'd268468224;
      11729: inst = 32'd201345876;
      11730: inst = 32'd203489279;
      11731: inst = 32'd136314880;
      11732: inst = 32'd268468224;
      11733: inst = 32'd201345877;
      11734: inst = 32'd203489279;
      11735: inst = 32'd136314880;
      11736: inst = 32'd268468224;
      11737: inst = 32'd201345878;
      11738: inst = 32'd203489279;
      11739: inst = 32'd136314880;
      11740: inst = 32'd268468224;
      11741: inst = 32'd201345879;
      11742: inst = 32'd203489279;
      11743: inst = 32'd136314880;
      11744: inst = 32'd268468224;
      11745: inst = 32'd201345880;
      11746: inst = 32'd203489279;
      11747: inst = 32'd136314880;
      11748: inst = 32'd268468224;
      11749: inst = 32'd201345881;
      11750: inst = 32'd203489279;
      11751: inst = 32'd136314880;
      11752: inst = 32'd268468224;
      11753: inst = 32'd201345882;
      11754: inst = 32'd203489279;
      11755: inst = 32'd136314880;
      11756: inst = 32'd268468224;
      11757: inst = 32'd201345883;
      11758: inst = 32'd203489279;
      11759: inst = 32'd136314880;
      11760: inst = 32'd268468224;
      11761: inst = 32'd201345884;
      11762: inst = 32'd203489279;
      11763: inst = 32'd136314880;
      11764: inst = 32'd268468224;
      11765: inst = 32'd201345885;
      11766: inst = 32'd203489279;
      11767: inst = 32'd136314880;
      11768: inst = 32'd268468224;
      11769: inst = 32'd201345886;
      11770: inst = 32'd203489279;
      11771: inst = 32'd136314880;
      11772: inst = 32'd268468224;
      11773: inst = 32'd201345887;
      11774: inst = 32'd203489279;
      11775: inst = 32'd136314880;
      11776: inst = 32'd268468224;
      11777: inst = 32'd201345888;
      11778: inst = 32'd203489278;
      11779: inst = 32'd136314880;
      11780: inst = 32'd268468224;
      11781: inst = 32'd201345889;
      11782: inst = 32'd203489279;
      11783: inst = 32'd136314880;
      11784: inst = 32'd268468224;
      11785: inst = 32'd201345890;
      11786: inst = 32'd203489247;
      11787: inst = 32'd136314880;
      11788: inst = 32'd268468224;
      11789: inst = 32'd201345891;
      11790: inst = 32'd203489279;
      11791: inst = 32'd136314880;
      11792: inst = 32'd268468224;
      11793: inst = 32'd201345892;
      11794: inst = 32'd203482840;
      11795: inst = 32'd136314880;
      11796: inst = 32'd268468224;
      11797: inst = 32'd201345893;
      11798: inst = 32'd203484886;
      11799: inst = 32'd136314880;
      11800: inst = 32'd268468224;
      11801: inst = 32'd201345894;
      11802: inst = 32'd203484853;
      11803: inst = 32'd136314880;
      11804: inst = 32'd268468224;
      11805: inst = 32'd201345895;
      11806: inst = 32'd203484854;
      11807: inst = 32'd136314880;
      11808: inst = 32'd268468224;
      11809: inst = 32'd201345896;
      11810: inst = 32'd203484887;
      11811: inst = 32'd136314880;
      11812: inst = 32'd268468224;
      11813: inst = 32'd201345897;
      11814: inst = 32'd203484854;
      11815: inst = 32'd136314880;
      11816: inst = 32'd268468224;
      11817: inst = 32'd201345898;
      11818: inst = 32'd203486902;
      11819: inst = 32'd136314880;
      11820: inst = 32'd268468224;
      11821: inst = 32'd201345899;
      11822: inst = 32'd203484854;
      11823: inst = 32'd136314880;
      11824: inst = 32'd268468224;
      11825: inst = 32'd201345900;
      11826: inst = 32'd203482839;
      11827: inst = 32'd136314880;
      11828: inst = 32'd268468224;
      11829: inst = 32'd201345901;
      11830: inst = 32'd203482838;
      11831: inst = 32'd136314880;
      11832: inst = 32'd268468224;
      11833: inst = 32'd201345902;
      11834: inst = 32'd203488915;
      11835: inst = 32'd136314880;
      11836: inst = 32'd268468224;
      11837: inst = 32'd201345903;
      11838: inst = 32'd203469573;
      11839: inst = 32'd136314880;
      11840: inst = 32'd268468224;
      11841: inst = 32'd201345904;
      11842: inst = 32'd203484133;
      11843: inst = 32'd136314880;
      11844: inst = 32'd268468224;
      11845: inst = 32'd201345905;
      11846: inst = 32'd203475911;
      11847: inst = 32'd136314880;
      11848: inst = 32'd268468224;
      11849: inst = 32'd201345906;
      11850: inst = 32'd203489048;
      11851: inst = 32'd136314880;
      11852: inst = 32'd268468224;
      11853: inst = 32'd201345907;
      11854: inst = 32'd203489082;
      11855: inst = 32'd136314880;
      11856: inst = 32'd268468224;
      11857: inst = 32'd201345908;
      11858: inst = 32'd203489113;
      11859: inst = 32'd136314880;
      11860: inst = 32'd268468224;
      11861: inst = 32'd201345909;
      11862: inst = 32'd203489078;
      11863: inst = 32'd136314880;
      11864: inst = 32'd268468224;
      11865: inst = 32'd201345910;
      11866: inst = 32'd203477991;
      11867: inst = 32'd136314880;
      11868: inst = 32'd268468224;
      11869: inst = 32'd201345911;
      11870: inst = 32'd203482087;
      11871: inst = 32'd136314880;
      11872: inst = 32'd268468224;
      11873: inst = 32'd201345912;
      11874: inst = 32'd203482023;
      11875: inst = 32'd136314880;
      11876: inst = 32'd268468224;
      11877: inst = 32'd201345913;
      11878: inst = 32'd203479975;
      11879: inst = 32'd136314880;
      11880: inst = 32'd268468224;
      11881: inst = 32'd201345914;
      11882: inst = 32'd203480006;
      11883: inst = 32'd136314880;
      11884: inst = 32'd268468224;
      11885: inst = 32'd201345915;
      11886: inst = 32'd203480037;
      11887: inst = 32'd136314880;
      11888: inst = 32'd268468224;
      11889: inst = 32'd201345916;
      11890: inst = 32'd203480003;
      11891: inst = 32'd136314880;
      11892: inst = 32'd268468224;
      11893: inst = 32'd201345917;
      11894: inst = 32'd203480004;
      11895: inst = 32'd136314880;
      11896: inst = 32'd268468224;
      11897: inst = 32'd201345918;
      11898: inst = 32'd203479974;
      11899: inst = 32'd136314880;
      11900: inst = 32'd268468224;
      11901: inst = 32'd201345919;
      11902: inst = 32'd203473605;
      11903: inst = 32'd136314880;
      11904: inst = 32'd268468224;
      11905: inst = 32'd201345920;
      11906: inst = 32'd203486871;
      11907: inst = 32'd136314880;
      11908: inst = 32'd268468224;
      11909: inst = 32'd201345921;
      11910: inst = 32'd203486903;
      11911: inst = 32'd136314880;
      11912: inst = 32'd268468224;
      11913: inst = 32'd201345922;
      11914: inst = 32'd203486903;
      11915: inst = 32'd136314880;
      11916: inst = 32'd268468224;
      11917: inst = 32'd201345923;
      11918: inst = 32'd203484854;
      11919: inst = 32'd136314880;
      11920: inst = 32'd268468224;
      11921: inst = 32'd201345924;
      11922: inst = 32'd203484854;
      11923: inst = 32'd136314880;
      11924: inst = 32'd268468224;
      11925: inst = 32'd201345925;
      11926: inst = 32'd203482807;
      11927: inst = 32'd136314880;
      11928: inst = 32'd268468224;
      11929: inst = 32'd201345926;
      11930: inst = 32'd203482840;
      11931: inst = 32'd136314880;
      11932: inst = 32'd268468224;
      11933: inst = 32'd201345927;
      11934: inst = 32'd203482874;
      11935: inst = 32'd136314880;
      11936: inst = 32'd268468224;
      11937: inst = 32'd201345928;
      11938: inst = 32'd203444841;
      11939: inst = 32'd136314880;
      11940: inst = 32'd268468224;
      11941: inst = 32'd201345929;
      11942: inst = 32'd203444875;
      11943: inst = 32'd136314880;
      11944: inst = 32'd268468224;
      11945: inst = 32'd201345930;
      11946: inst = 32'd203480764;
      11947: inst = 32'd136314880;
      11948: inst = 32'd268468224;
      11949: inst = 32'd201345931;
      11950: inst = 32'd203442763;
      11951: inst = 32'd136314880;
      11952: inst = 32'd268468224;
      11953: inst = 32'd201345932;
      11954: inst = 32'd203444908;
      11955: inst = 32'd136314880;
      11956: inst = 32'd268468224;
      11957: inst = 32'd201345933;
      11958: inst = 32'd203478715;
      11959: inst = 32'd136314880;
      11960: inst = 32'd268468224;
      11961: inst = 32'd201345934;
      11962: inst = 32'd203482972;
      11963: inst = 32'd136314880;
      11964: inst = 32'd268468224;
      11965: inst = 32'd201345935;
      11966: inst = 32'd203480827;
      11967: inst = 32'd136314880;
      11968: inst = 32'd268468224;
      11969: inst = 32'd201345936;
      11970: inst = 32'd203484854;
      11971: inst = 32'd136314880;
      11972: inst = 32'd268468224;
      11973: inst = 32'd201345937;
      11974: inst = 32'd203484854;
      11975: inst = 32'd136314880;
      11976: inst = 32'd268468224;
      11977: inst = 32'd201345938;
      11978: inst = 32'd203484854;
      11979: inst = 32'd136314880;
      11980: inst = 32'd268468224;
      11981: inst = 32'd201345939;
      11982: inst = 32'd203484854;
      11983: inst = 32'd136314880;
      11984: inst = 32'd268468224;
      11985: inst = 32'd201345940;
      11986: inst = 32'd203484854;
      11987: inst = 32'd136314880;
      11988: inst = 32'd268468224;
      11989: inst = 32'd201345941;
      11990: inst = 32'd203484854;
      11991: inst = 32'd136314880;
      11992: inst = 32'd268468224;
      11993: inst = 32'd201345942;
      11994: inst = 32'd203484854;
      11995: inst = 32'd136314880;
      11996: inst = 32'd268468224;
      11997: inst = 32'd201345943;
      11998: inst = 32'd203484854;
      11999: inst = 32'd136314880;
      12000: inst = 32'd268468224;
      12001: inst = 32'd201345944;
      12002: inst = 32'd203484854;
      12003: inst = 32'd136314880;
      12004: inst = 32'd268468224;
      12005: inst = 32'd201345945;
      12006: inst = 32'd203484854;
      12007: inst = 32'd136314880;
      12008: inst = 32'd268468224;
      12009: inst = 32'd201345946;
      12010: inst = 32'd203484855;
      12011: inst = 32'd136314880;
      12012: inst = 32'd268468224;
      12013: inst = 32'd201345947;
      12014: inst = 32'd203482808;
      12015: inst = 32'd136314880;
      12016: inst = 32'd268468224;
      12017: inst = 32'd201345948;
      12018: inst = 32'd203489278;
      12019: inst = 32'd136314880;
      12020: inst = 32'd268468224;
      12021: inst = 32'd201345949;
      12022: inst = 32'd203489279;
      12023: inst = 32'd136314880;
      12024: inst = 32'd268468224;
      12025: inst = 32'd201345950;
      12026: inst = 32'd203489279;
      12027: inst = 32'd136314880;
      12028: inst = 32'd268468224;
      12029: inst = 32'd201345951;
      12030: inst = 32'd203489279;
      12031: inst = 32'd136314880;
      12032: inst = 32'd268468224;
      12033: inst = 32'd201345952;
      12034: inst = 32'd203489279;
      12035: inst = 32'd136314880;
      12036: inst = 32'd268468224;
      12037: inst = 32'd201345953;
      12038: inst = 32'd203489279;
      12039: inst = 32'd136314880;
      12040: inst = 32'd268468224;
      12041: inst = 32'd201345954;
      12042: inst = 32'd203489279;
      12043: inst = 32'd136314880;
      12044: inst = 32'd268468224;
      12045: inst = 32'd201345955;
      12046: inst = 32'd203489279;
      12047: inst = 32'd136314880;
      12048: inst = 32'd268468224;
      12049: inst = 32'd201345956;
      12050: inst = 32'd203489279;
      12051: inst = 32'd136314880;
      12052: inst = 32'd268468224;
      12053: inst = 32'd201345957;
      12054: inst = 32'd203489279;
      12055: inst = 32'd136314880;
      12056: inst = 32'd268468224;
      12057: inst = 32'd201345958;
      12058: inst = 32'd203489279;
      12059: inst = 32'd136314880;
      12060: inst = 32'd268468224;
      12061: inst = 32'd201345959;
      12062: inst = 32'd203489279;
      12063: inst = 32'd136314880;
      12064: inst = 32'd268468224;
      12065: inst = 32'd201345960;
      12066: inst = 32'd203489279;
      12067: inst = 32'd136314880;
      12068: inst = 32'd268468224;
      12069: inst = 32'd201345961;
      12070: inst = 32'd203489279;
      12071: inst = 32'd136314880;
      12072: inst = 32'd268468224;
      12073: inst = 32'd201345962;
      12074: inst = 32'd203489279;
      12075: inst = 32'd136314880;
      12076: inst = 32'd268468224;
      12077: inst = 32'd201345963;
      12078: inst = 32'd203489279;
      12079: inst = 32'd136314880;
      12080: inst = 32'd268468224;
      12081: inst = 32'd201345964;
      12082: inst = 32'd203489279;
      12083: inst = 32'd136314880;
      12084: inst = 32'd268468224;
      12085: inst = 32'd201345965;
      12086: inst = 32'd203489279;
      12087: inst = 32'd136314880;
      12088: inst = 32'd268468224;
      12089: inst = 32'd201345966;
      12090: inst = 32'd203489279;
      12091: inst = 32'd136314880;
      12092: inst = 32'd268468224;
      12093: inst = 32'd201345967;
      12094: inst = 32'd203489279;
      12095: inst = 32'd136314880;
      12096: inst = 32'd268468224;
      12097: inst = 32'd201345968;
      12098: inst = 32'd203489279;
      12099: inst = 32'd136314880;
      12100: inst = 32'd268468224;
      12101: inst = 32'd201345969;
      12102: inst = 32'd203489279;
      12103: inst = 32'd136314880;
      12104: inst = 32'd268468224;
      12105: inst = 32'd201345970;
      12106: inst = 32'd203489279;
      12107: inst = 32'd136314880;
      12108: inst = 32'd268468224;
      12109: inst = 32'd201345971;
      12110: inst = 32'd203489279;
      12111: inst = 32'd136314880;
      12112: inst = 32'd268468224;
      12113: inst = 32'd201345972;
      12114: inst = 32'd203489279;
      12115: inst = 32'd136314880;
      12116: inst = 32'd268468224;
      12117: inst = 32'd201345973;
      12118: inst = 32'd203489279;
      12119: inst = 32'd136314880;
      12120: inst = 32'd268468224;
      12121: inst = 32'd201345974;
      12122: inst = 32'd203489279;
      12123: inst = 32'd136314880;
      12124: inst = 32'd268468224;
      12125: inst = 32'd201345975;
      12126: inst = 32'd203489279;
      12127: inst = 32'd136314880;
      12128: inst = 32'd268468224;
      12129: inst = 32'd201345976;
      12130: inst = 32'd203489279;
      12131: inst = 32'd136314880;
      12132: inst = 32'd268468224;
      12133: inst = 32'd201345977;
      12134: inst = 32'd203489279;
      12135: inst = 32'd136314880;
      12136: inst = 32'd268468224;
      12137: inst = 32'd201345978;
      12138: inst = 32'd203489279;
      12139: inst = 32'd136314880;
      12140: inst = 32'd268468224;
      12141: inst = 32'd201345979;
      12142: inst = 32'd203489279;
      12143: inst = 32'd136314880;
      12144: inst = 32'd268468224;
      12145: inst = 32'd201345980;
      12146: inst = 32'd203489279;
      12147: inst = 32'd136314880;
      12148: inst = 32'd268468224;
      12149: inst = 32'd201345981;
      12150: inst = 32'd203489279;
      12151: inst = 32'd136314880;
      12152: inst = 32'd268468224;
      12153: inst = 32'd201345982;
      12154: inst = 32'd203489279;
      12155: inst = 32'd136314880;
      12156: inst = 32'd268468224;
      12157: inst = 32'd201345983;
      12158: inst = 32'd203489279;
      12159: inst = 32'd136314880;
      12160: inst = 32'd268468224;
      12161: inst = 32'd201345984;
      12162: inst = 32'd203489278;
      12163: inst = 32'd136314880;
      12164: inst = 32'd268468224;
      12165: inst = 32'd201345985;
      12166: inst = 32'd203489279;
      12167: inst = 32'd136314880;
      12168: inst = 32'd268468224;
      12169: inst = 32'd201345986;
      12170: inst = 32'd203489247;
      12171: inst = 32'd136314880;
      12172: inst = 32'd268468224;
      12173: inst = 32'd201345987;
      12174: inst = 32'd203489278;
      12175: inst = 32'd136314880;
      12176: inst = 32'd268468224;
      12177: inst = 32'd201345988;
      12178: inst = 32'd203482839;
      12179: inst = 32'd136314880;
      12180: inst = 32'd268468224;
      12181: inst = 32'd201345989;
      12182: inst = 32'd203484886;
      12183: inst = 32'd136314880;
      12184: inst = 32'd268468224;
      12185: inst = 32'd201345990;
      12186: inst = 32'd203484853;
      12187: inst = 32'd136314880;
      12188: inst = 32'd268468224;
      12189: inst = 32'd201345991;
      12190: inst = 32'd203484854;
      12191: inst = 32'd136314880;
      12192: inst = 32'd268468224;
      12193: inst = 32'd201345992;
      12194: inst = 32'd203484887;
      12195: inst = 32'd136314880;
      12196: inst = 32'd268468224;
      12197: inst = 32'd201345993;
      12198: inst = 32'd203484854;
      12199: inst = 32'd136314880;
      12200: inst = 32'd268468224;
      12201: inst = 32'd201345994;
      12202: inst = 32'd203486902;
      12203: inst = 32'd136314880;
      12204: inst = 32'd268468224;
      12205: inst = 32'd201345995;
      12206: inst = 32'd203484823;
      12207: inst = 32'd136314880;
      12208: inst = 32'd268468224;
      12209: inst = 32'd201345996;
      12210: inst = 32'd203482839;
      12211: inst = 32'd136314880;
      12212: inst = 32'd268468224;
      12213: inst = 32'd201345997;
      12214: inst = 32'd203482838;
      12215: inst = 32'd136314880;
      12216: inst = 32'd268468224;
      12217: inst = 32'd201345998;
      12218: inst = 32'd203488915;
      12219: inst = 32'd136314880;
      12220: inst = 32'd268468224;
      12221: inst = 32'd201345999;
      12222: inst = 32'd203469573;
      12223: inst = 32'd136314880;
      12224: inst = 32'd268468224;
      12225: inst = 32'd201346000;
      12226: inst = 32'd203484002;
      12227: inst = 32'd136314880;
      12228: inst = 32'd268468224;
      12229: inst = 32'd201346001;
      12230: inst = 32'd203482022;
      12231: inst = 32'd136314880;
      12232: inst = 32'd268468224;
      12233: inst = 32'd201346002;
      12234: inst = 32'd203477962;
      12235: inst = 32'd136314880;
      12236: inst = 32'd268468224;
      12237: inst = 32'd201346003;
      12238: inst = 32'd203475948;
      12239: inst = 32'd136314880;
      12240: inst = 32'd268468224;
      12241: inst = 32'd201346004;
      12242: inst = 32'd203473866;
      12243: inst = 32'd136314880;
      12244: inst = 32'd268468224;
      12245: inst = 32'd201346005;
      12246: inst = 32'd203475879;
      12247: inst = 32'd136314880;
      12248: inst = 32'd268468224;
      12249: inst = 32'd201346006;
      12250: inst = 32'd203480005;
      12251: inst = 32'd136314880;
      12252: inst = 32'd268468224;
      12253: inst = 32'd201346007;
      12254: inst = 32'd203479972;
      12255: inst = 32'd136314880;
      12256: inst = 32'd268468224;
      12257: inst = 32'd201346008;
      12258: inst = 32'd203482021;
      12259: inst = 32'd136314880;
      12260: inst = 32'd268468224;
      12261: inst = 32'd201346009;
      12262: inst = 32'd203482021;
      12263: inst = 32'd136314880;
      12264: inst = 32'd268468224;
      12265: inst = 32'd201346010;
      12266: inst = 32'd203482020;
      12267: inst = 32'd136314880;
      12268: inst = 32'd268468224;
      12269: inst = 32'd201346011;
      12270: inst = 32'd203482051;
      12271: inst = 32'd136314880;
      12272: inst = 32'd268468224;
      12273: inst = 32'd201346012;
      12274: inst = 32'd203482049;
      12275: inst = 32'd136314880;
      12276: inst = 32'd268468224;
      12277: inst = 32'd201346013;
      12278: inst = 32'd203482082;
      12279: inst = 32'd136314880;
      12280: inst = 32'd268468224;
      12281: inst = 32'd201346014;
      12282: inst = 32'd203480004;
      12283: inst = 32'd136314880;
      12284: inst = 32'd268468224;
      12285: inst = 32'd201346015;
      12286: inst = 32'd203471619;
      12287: inst = 32'd136314880;
      12288: inst = 32'd268468224;
      12289: inst = 32'd201346016;
      12290: inst = 32'd203484822;
      12291: inst = 32'd136314880;
      12292: inst = 32'd268468224;
      12293: inst = 32'd201346017;
      12294: inst = 32'd203486935;
      12295: inst = 32'd136314880;
      12296: inst = 32'd268468224;
      12297: inst = 32'd201346018;
      12298: inst = 32'd203486967;
      12299: inst = 32'd136314880;
      12300: inst = 32'd268468224;
      12301: inst = 32'd201346019;
      12302: inst = 32'd203484855;
      12303: inst = 32'd136314880;
      12304: inst = 32'd268468224;
      12305: inst = 32'd201346020;
      12306: inst = 32'd203482807;
      12307: inst = 32'd136314880;
      12308: inst = 32'd268468224;
      12309: inst = 32'd201346021;
      12310: inst = 32'd203482808;
      12311: inst = 32'd136314880;
      12312: inst = 32'd268468224;
      12313: inst = 32'd201346022;
      12314: inst = 32'd203482808;
      12315: inst = 32'd136314880;
      12316: inst = 32'd268468224;
      12317: inst = 32'd201346023;
      12318: inst = 32'd203482874;
      12319: inst = 32'd136314880;
      12320: inst = 32'd268468224;
      12321: inst = 32'd201346024;
      12322: inst = 32'd203482874;
      12323: inst = 32'd136314880;
      12324: inst = 32'd268468224;
      12325: inst = 32'd201346025;
      12326: inst = 32'd203482907;
      12327: inst = 32'd136314880;
      12328: inst = 32'd268468224;
      12329: inst = 32'd201346026;
      12330: inst = 32'd203482874;
      12331: inst = 32'd136314880;
      12332: inst = 32'd268468224;
      12333: inst = 32'd201346027;
      12334: inst = 32'd203482842;
      12335: inst = 32'd136314880;
      12336: inst = 32'd268468224;
      12337: inst = 32'd201346028;
      12338: inst = 32'd203482842;
      12339: inst = 32'd136314880;
      12340: inst = 32'd268468224;
      12341: inst = 32'd201346029;
      12342: inst = 32'd203484988;
      12343: inst = 32'd136314880;
      12344: inst = 32'd268468224;
      12345: inst = 32'd201346030;
      12346: inst = 32'd203482810;
      12347: inst = 32'd136314880;
      12348: inst = 32'd268468224;
      12349: inst = 32'd201346031;
      12350: inst = 32'd203482843;
      12351: inst = 32'd136314880;
      12352: inst = 32'd268468224;
      12353: inst = 32'd201346032;
      12354: inst = 32'd203486904;
      12355: inst = 32'd136314880;
      12356: inst = 32'd268468224;
      12357: inst = 32'd201346033;
      12358: inst = 32'd203486934;
      12359: inst = 32'd136314880;
      12360: inst = 32'd268468224;
      12361: inst = 32'd201346034;
      12362: inst = 32'd203484853;
      12363: inst = 32'd136314880;
      12364: inst = 32'd268468224;
      12365: inst = 32'd201346035;
      12366: inst = 32'd203484886;
      12367: inst = 32'd136314880;
      12368: inst = 32'd268468224;
      12369: inst = 32'd201346036;
      12370: inst = 32'd203482774;
      12371: inst = 32'd136314880;
      12372: inst = 32'd268468224;
      12373: inst = 32'd201346037;
      12374: inst = 32'd203484855;
      12375: inst = 32'd136314880;
      12376: inst = 32'd268468224;
      12377: inst = 32'd201346038;
      12378: inst = 32'd203484887;
      12379: inst = 32'd136314880;
      12380: inst = 32'd268468224;
      12381: inst = 32'd201346039;
      12382: inst = 32'd203482806;
      12383: inst = 32'd136314880;
      12384: inst = 32'd268468224;
      12385: inst = 32'd201346040;
      12386: inst = 32'd203484887;
      12387: inst = 32'd136314880;
      12388: inst = 32'd268468224;
      12389: inst = 32'd201346041;
      12390: inst = 32'd203482776;
      12391: inst = 32'd136314880;
      12392: inst = 32'd268468224;
      12393: inst = 32'd201346042;
      12394: inst = 32'd203476405;
      12395: inst = 32'd136314880;
      12396: inst = 32'd268468224;
      12397: inst = 32'd201346043;
      12398: inst = 32'd203472212;
      12399: inst = 32'd136314880;
      12400: inst = 32'd268468224;
      12401: inst = 32'd201346044;
      12402: inst = 32'd203474324;
      12403: inst = 32'd136314880;
      12404: inst = 32'd268468224;
      12405: inst = 32'd201346045;
      12406: inst = 32'd203472276;
      12407: inst = 32'd136314880;
      12408: inst = 32'd268468224;
      12409: inst = 32'd201346046;
      12410: inst = 32'd203472277;
      12411: inst = 32'd136314880;
      12412: inst = 32'd268468224;
      12413: inst = 32'd201346047;
      12414: inst = 32'd203472246;
      12415: inst = 32'd136314880;
      12416: inst = 32'd268468224;
      12417: inst = 32'd201346048;
      12418: inst = 32'd203474293;
      12419: inst = 32'd136314880;
      12420: inst = 32'd268468224;
      12421: inst = 32'd201346049;
      12422: inst = 32'd203472245;
      12423: inst = 32'd136314880;
      12424: inst = 32'd268468224;
      12425: inst = 32'd201346050;
      12426: inst = 32'd203472244;
      12427: inst = 32'd136314880;
      12428: inst = 32'd268468224;
      12429: inst = 32'd201346051;
      12430: inst = 32'd203472276;
      12431: inst = 32'd136314880;
      12432: inst = 32'd268468224;
      12433: inst = 32'd201346052;
      12434: inst = 32'd203470228;
      12435: inst = 32'd136314880;
      12436: inst = 32'd268468224;
      12437: inst = 32'd201346053;
      12438: inst = 32'd203470228;
      12439: inst = 32'd136314880;
      12440: inst = 32'd268468224;
      12441: inst = 32'd201346054;
      12442: inst = 32'd203470260;
      12443: inst = 32'd136314880;
      12444: inst = 32'd268468224;
      12445: inst = 32'd201346055;
      12446: inst = 32'd203472308;
      12447: inst = 32'd136314880;
      12448: inst = 32'd268468224;
      12449: inst = 32'd201346056;
      12450: inst = 32'd203472276;
      12451: inst = 32'd136314880;
      12452: inst = 32'd268468224;
      12453: inst = 32'd201346057;
      12454: inst = 32'd203472276;
      12455: inst = 32'd136314880;
      12456: inst = 32'd268468224;
      12457: inst = 32'd201346058;
      12458: inst = 32'd203472276;
      12459: inst = 32'd136314880;
      12460: inst = 32'd268468224;
      12461: inst = 32'd201346059;
      12462: inst = 32'd203472276;
      12463: inst = 32'd136314880;
      12464: inst = 32'd268468224;
      12465: inst = 32'd201346060;
      12466: inst = 32'd203470228;
      12467: inst = 32'd136314880;
      12468: inst = 32'd268468224;
      12469: inst = 32'd201346061;
      12470: inst = 32'd203470260;
      12471: inst = 32'd136314880;
      12472: inst = 32'd268468224;
      12473: inst = 32'd201346062;
      12474: inst = 32'd203470259;
      12475: inst = 32'd136314880;
      12476: inst = 32'd268468224;
      12477: inst = 32'd201346063;
      12478: inst = 32'd203470259;
      12479: inst = 32'd136314880;
      12480: inst = 32'd268468224;
      12481: inst = 32'd201346064;
      12482: inst = 32'd203470259;
      12483: inst = 32'd136314880;
      12484: inst = 32'd268468224;
      12485: inst = 32'd201346065;
      12486: inst = 32'd203470259;
      12487: inst = 32'd136314880;
      12488: inst = 32'd268468224;
      12489: inst = 32'd201346066;
      12490: inst = 32'd203470260;
      12491: inst = 32'd136314880;
      12492: inst = 32'd268468224;
      12493: inst = 32'd201346067;
      12494: inst = 32'd203470228;
      12495: inst = 32'd136314880;
      12496: inst = 32'd268468224;
      12497: inst = 32'd201346068;
      12498: inst = 32'd203472276;
      12499: inst = 32'd136314880;
      12500: inst = 32'd268468224;
      12501: inst = 32'd201346069;
      12502: inst = 32'd203472276;
      12503: inst = 32'd136314880;
      12504: inst = 32'd268468224;
      12505: inst = 32'd201346070;
      12506: inst = 32'd203472276;
      12507: inst = 32'd136314880;
      12508: inst = 32'd268468224;
      12509: inst = 32'd201346071;
      12510: inst = 32'd203472276;
      12511: inst = 32'd136314880;
      12512: inst = 32'd268468224;
      12513: inst = 32'd201346072;
      12514: inst = 32'd203472308;
      12515: inst = 32'd136314880;
      12516: inst = 32'd268468224;
      12517: inst = 32'd201346073;
      12518: inst = 32'd203470260;
      12519: inst = 32'd136314880;
      12520: inst = 32'd268468224;
      12521: inst = 32'd201346074;
      12522: inst = 32'd203470228;
      12523: inst = 32'd136314880;
      12524: inst = 32'd268468224;
      12525: inst = 32'd201346075;
      12526: inst = 32'd203470228;
      12527: inst = 32'd136314880;
      12528: inst = 32'd268468224;
      12529: inst = 32'd201346076;
      12530: inst = 32'd203472276;
      12531: inst = 32'd136314880;
      12532: inst = 32'd268468224;
      12533: inst = 32'd201346077;
      12534: inst = 32'd203472244;
      12535: inst = 32'd136314880;
      12536: inst = 32'd268468224;
      12537: inst = 32'd201346078;
      12538: inst = 32'd203472245;
      12539: inst = 32'd136314880;
      12540: inst = 32'd268468224;
      12541: inst = 32'd201346079;
      12542: inst = 32'd203474293;
      12543: inst = 32'd136314880;
      12544: inst = 32'd268468224;
      12545: inst = 32'd201346080;
      12546: inst = 32'd203472275;
      12547: inst = 32'd136314880;
      12548: inst = 32'd268468224;
      12549: inst = 32'd201346081;
      12550: inst = 32'd203474323;
      12551: inst = 32'd136314880;
      12552: inst = 32'd268468224;
      12553: inst = 32'd201346082;
      12554: inst = 32'd203474323;
      12555: inst = 32'd136314880;
      12556: inst = 32'd268468224;
      12557: inst = 32'd201346083;
      12558: inst = 32'd203474323;
      12559: inst = 32'd136314880;
      12560: inst = 32'd268468224;
      12561: inst = 32'd201346084;
      12562: inst = 32'd203472242;
      12563: inst = 32'd136314880;
      12564: inst = 32'd268468224;
      12565: inst = 32'd201346085;
      12566: inst = 32'd203476403;
      12567: inst = 32'd136314880;
      12568: inst = 32'd268468224;
      12569: inst = 32'd201346086;
      12570: inst = 32'd203484822;
      12571: inst = 32'd136314880;
      12572: inst = 32'd268468224;
      12573: inst = 32'd201346087;
      12574: inst = 32'd203484855;
      12575: inst = 32'd136314880;
      12576: inst = 32'd268468224;
      12577: inst = 32'd201346088;
      12578: inst = 32'd203482839;
      12579: inst = 32'd136314880;
      12580: inst = 32'd268468224;
      12581: inst = 32'd201346089;
      12582: inst = 32'd203484854;
      12583: inst = 32'd136314880;
      12584: inst = 32'd268468224;
      12585: inst = 32'd201346090;
      12586: inst = 32'd203486901;
      12587: inst = 32'd136314880;
      12588: inst = 32'd268468224;
      12589: inst = 32'd201346091;
      12590: inst = 32'd203484854;
      12591: inst = 32'd136314880;
      12592: inst = 32'd268468224;
      12593: inst = 32'd201346092;
      12594: inst = 32'd203482840;
      12595: inst = 32'd136314880;
      12596: inst = 32'd268468224;
      12597: inst = 32'd201346093;
      12598: inst = 32'd203484855;
      12599: inst = 32'd136314880;
      12600: inst = 32'd268468224;
      12601: inst = 32'd201346094;
      12602: inst = 32'd203488883;
      12603: inst = 32'd136314880;
      12604: inst = 32'd268468224;
      12605: inst = 32'd201346095;
      12606: inst = 32'd203471619;
      12607: inst = 32'd136314880;
      12608: inst = 32'd268468224;
      12609: inst = 32'd201346096;
      12610: inst = 32'd203480005;
      12611: inst = 32'd136314880;
      12612: inst = 32'd268468224;
      12613: inst = 32'd201346097;
      12614: inst = 32'd203480005;
      12615: inst = 32'd136314880;
      12616: inst = 32'd268468224;
      12617: inst = 32'd201346098;
      12618: inst = 32'd203480005;
      12619: inst = 32'd136314880;
      12620: inst = 32'd268468224;
      12621: inst = 32'd201346099;
      12622: inst = 32'd203480005;
      12623: inst = 32'd136314880;
      12624: inst = 32'd268468224;
      12625: inst = 32'd201346100;
      12626: inst = 32'd203480006;
      12627: inst = 32'd136314880;
      12628: inst = 32'd268468224;
      12629: inst = 32'd201346101;
      12630: inst = 32'd203480006;
      12631: inst = 32'd136314880;
      12632: inst = 32'd268468224;
      12633: inst = 32'd201346102;
      12634: inst = 32'd203480006;
      12635: inst = 32'd136314880;
      12636: inst = 32'd268468224;
      12637: inst = 32'd201346103;
      12638: inst = 32'd203480006;
      12639: inst = 32'd136314880;
      12640: inst = 32'd268468224;
      12641: inst = 32'd201346104;
      12642: inst = 32'd203477893;
      12643: inst = 32'd136314880;
      12644: inst = 32'd268468224;
      12645: inst = 32'd201346105;
      12646: inst = 32'd203480071;
      12647: inst = 32'd136314880;
      12648: inst = 32'd268468224;
      12649: inst = 32'd201346106;
      12650: inst = 32'd203477959;
      12651: inst = 32'd136314880;
      12652: inst = 32'd268468224;
      12653: inst = 32'd201346107;
      12654: inst = 32'd203475878;
      12655: inst = 32'd136314880;
      12656: inst = 32'd268468224;
      12657: inst = 32'd201346108;
      12658: inst = 32'd203480104;
      12659: inst = 32'd136314880;
      12660: inst = 32'd268468224;
      12661: inst = 32'd201346109;
      12662: inst = 32'd203477959;
      12663: inst = 32'd136314880;
      12664: inst = 32'd268468224;
      12665: inst = 32'd201346110;
      12666: inst = 32'd203475911;
      12667: inst = 32'd136314880;
      12668: inst = 32'd268468224;
      12669: inst = 32'd201346111;
      12670: inst = 32'd203471620;
      12671: inst = 32'd136314880;
      12672: inst = 32'd268468224;
      12673: inst = 32'd201346112;
      12674: inst = 32'd203489048;
      12675: inst = 32'd136314880;
      12676: inst = 32'd268468224;
      12677: inst = 32'd201346113;
      12678: inst = 32'd203484855;
      12679: inst = 32'd136314880;
      12680: inst = 32'd268468224;
      12681: inst = 32'd201346114;
      12682: inst = 32'd203482774;
      12683: inst = 32'd136314880;
      12684: inst = 32'd268468224;
      12685: inst = 32'd201346115;
      12686: inst = 32'd203482807;
      12687: inst = 32'd136314880;
      12688: inst = 32'd268468224;
      12689: inst = 32'd201346116;
      12690: inst = 32'd203484888;
      12691: inst = 32'd136314880;
      12692: inst = 32'd268468224;
      12693: inst = 32'd201346117;
      12694: inst = 32'd203484921;
      12695: inst = 32'd136314880;
      12696: inst = 32'd268468224;
      12697: inst = 32'd201346118;
      12698: inst = 32'd203482841;
      12699: inst = 32'd136314880;
      12700: inst = 32'd268468224;
      12701: inst = 32'd201346119;
      12702: inst = 32'd203480793;
      12703: inst = 32'd136314880;
      12704: inst = 32'd268468224;
      12705: inst = 32'd201346120;
      12706: inst = 32'd203444840;
      12707: inst = 32'd136314880;
      12708: inst = 32'd268468224;
      12709: inst = 32'd201346121;
      12710: inst = 32'd203482907;
      12711: inst = 32'd136314880;
      12712: inst = 32'd268468224;
      12713: inst = 32'd201346122;
      12714: inst = 32'd203444841;
      12715: inst = 32'd136314880;
      12716: inst = 32'd268468224;
      12717: inst = 32'd201346123;
      12718: inst = 32'd203480794;
      12719: inst = 32'd136314880;
      12720: inst = 32'd268468224;
      12721: inst = 32'd201346124;
      12722: inst = 32'd203446954;
      12723: inst = 32'd136314880;
      12724: inst = 32'd268468224;
      12725: inst = 32'd201346125;
      12726: inst = 32'd203480730;
      12727: inst = 32'd136314880;
      12728: inst = 32'd268468224;
      12729: inst = 32'd201346126;
      12730: inst = 32'd203480730;
      12731: inst = 32'd136314880;
      12732: inst = 32'd268468224;
      12733: inst = 32'd201346127;
      12734: inst = 32'd203482842;
      12735: inst = 32'd136314880;
      12736: inst = 32'd268468224;
      12737: inst = 32'd201346128;
      12738: inst = 32'd203484792;
      12739: inst = 32'd136314880;
      12740: inst = 32'd268468224;
      12741: inst = 32'd201346129;
      12742: inst = 32'd203484823;
      12743: inst = 32'd136314880;
      12744: inst = 32'd268468224;
      12745: inst = 32'd201346130;
      12746: inst = 32'd203482774;
      12747: inst = 32'd136314880;
      12748: inst = 32'd268468224;
      12749: inst = 32'd201346131;
      12750: inst = 32'd203484887;
      12751: inst = 32'd136314880;
      12752: inst = 32'd268468224;
      12753: inst = 32'd201346132;
      12754: inst = 32'd203484856;
      12755: inst = 32'd136314880;
      12756: inst = 32'd268468224;
      12757: inst = 32'd201346133;
      12758: inst = 32'd203482808;
      12759: inst = 32'd136314880;
      12760: inst = 32'd268468224;
      12761: inst = 32'd201346134;
      12762: inst = 32'd203480694;
      12763: inst = 32'd136314880;
      12764: inst = 32'd268468224;
      12765: inst = 32'd201346135;
      12766: inst = 32'd203484919;
      12767: inst = 32'd136314880;
      12768: inst = 32'd268468224;
      12769: inst = 32'd201346136;
      12770: inst = 32'd203482806;
      12771: inst = 32'd136314880;
      12772: inst = 32'd268468224;
      12773: inst = 32'd201346137;
      12774: inst = 32'd203484888;
      12775: inst = 32'd136314880;
      12776: inst = 32'd268468224;
      12777: inst = 32'd201346138;
      12778: inst = 32'd203482776;
      12779: inst = 32'd136314880;
      12780: inst = 32'd268468224;
      12781: inst = 32'd201346139;
      12782: inst = 32'd203482776;
      12783: inst = 32'd136314880;
      12784: inst = 32'd268468224;
      12785: inst = 32'd201346140;
      12786: inst = 32'd203484856;
      12787: inst = 32'd136314880;
      12788: inst = 32'd268468224;
      12789: inst = 32'd201346141;
      12790: inst = 32'd203482807;
      12791: inst = 32'd136314880;
      12792: inst = 32'd268468224;
      12793: inst = 32'd201346142;
      12794: inst = 32'd203482808;
      12795: inst = 32'd136314880;
      12796: inst = 32'd268468224;
      12797: inst = 32'd201346143;
      12798: inst = 32'd203482810;
      12799: inst = 32'd136314880;
      12800: inst = 32'd268468224;
      12801: inst = 32'd201346144;
      12802: inst = 32'd203484824;
      12803: inst = 32'd136314880;
      12804: inst = 32'd268468224;
      12805: inst = 32'd201346145;
      12806: inst = 32'd203484857;
      12807: inst = 32'd136314880;
      12808: inst = 32'd268468224;
      12809: inst = 32'd201346146;
      12810: inst = 32'd203484889;
      12811: inst = 32'd136314880;
      12812: inst = 32'd268468224;
      12813: inst = 32'd201346147;
      12814: inst = 32'd203484920;
      12815: inst = 32'd136314880;
      12816: inst = 32'd268468224;
      12817: inst = 32'd201346148;
      12818: inst = 32'd203482872;
      12819: inst = 32'd136314880;
      12820: inst = 32'd268468224;
      12821: inst = 32'd201346149;
      12822: inst = 32'd203482872;
      12823: inst = 32'd136314880;
      12824: inst = 32'd268468224;
      12825: inst = 32'd201346150;
      12826: inst = 32'd203482840;
      12827: inst = 32'd136314880;
      12828: inst = 32'd268468224;
      12829: inst = 32'd201346151;
      12830: inst = 32'd203482808;
      12831: inst = 32'd136314880;
      12832: inst = 32'd268468224;
      12833: inst = 32'd201346152;
      12834: inst = 32'd203482840;
      12835: inst = 32'd136314880;
      12836: inst = 32'd268468224;
      12837: inst = 32'd201346153;
      12838: inst = 32'd203484889;
      12839: inst = 32'd136314880;
      12840: inst = 32'd268468224;
      12841: inst = 32'd201346154;
      12842: inst = 32'd203484889;
      12843: inst = 32'd136314880;
      12844: inst = 32'd268468224;
      12845: inst = 32'd201346155;
      12846: inst = 32'd203482841;
      12847: inst = 32'd136314880;
      12848: inst = 32'd268468224;
      12849: inst = 32'd201346156;
      12850: inst = 32'd203482840;
      12851: inst = 32'd136314880;
      12852: inst = 32'd268468224;
      12853: inst = 32'd201346157;
      12854: inst = 32'd203482872;
      12855: inst = 32'd136314880;
      12856: inst = 32'd268468224;
      12857: inst = 32'd201346158;
      12858: inst = 32'd203482872;
      12859: inst = 32'd136314880;
      12860: inst = 32'd268468224;
      12861: inst = 32'd201346159;
      12862: inst = 32'd203480824;
      12863: inst = 32'd136314880;
      12864: inst = 32'd268468224;
      12865: inst = 32'd201346160;
      12866: inst = 32'd203480824;
      12867: inst = 32'd136314880;
      12868: inst = 32'd268468224;
      12869: inst = 32'd201346161;
      12870: inst = 32'd203482872;
      12871: inst = 32'd136314880;
      12872: inst = 32'd268468224;
      12873: inst = 32'd201346162;
      12874: inst = 32'd203482872;
      12875: inst = 32'd136314880;
      12876: inst = 32'd268468224;
      12877: inst = 32'd201346163;
      12878: inst = 32'd203482840;
      12879: inst = 32'd136314880;
      12880: inst = 32'd268468224;
      12881: inst = 32'd201346164;
      12882: inst = 32'd203482841;
      12883: inst = 32'd136314880;
      12884: inst = 32'd268468224;
      12885: inst = 32'd201346165;
      12886: inst = 32'd203484889;
      12887: inst = 32'd136314880;
      12888: inst = 32'd268468224;
      12889: inst = 32'd201346166;
      12890: inst = 32'd203484889;
      12891: inst = 32'd136314880;
      12892: inst = 32'd268468224;
      12893: inst = 32'd201346167;
      12894: inst = 32'd203482840;
      12895: inst = 32'd136314880;
      12896: inst = 32'd268468224;
      12897: inst = 32'd201346168;
      12898: inst = 32'd203482808;
      12899: inst = 32'd136314880;
      12900: inst = 32'd268468224;
      12901: inst = 32'd201346169;
      12902: inst = 32'd203482840;
      12903: inst = 32'd136314880;
      12904: inst = 32'd268468224;
      12905: inst = 32'd201346170;
      12906: inst = 32'd203482872;
      12907: inst = 32'd136314880;
      12908: inst = 32'd268468224;
      12909: inst = 32'd201346171;
      12910: inst = 32'd203482872;
      12911: inst = 32'd136314880;
      12912: inst = 32'd268468224;
      12913: inst = 32'd201346172;
      12914: inst = 32'd203484920;
      12915: inst = 32'd136314880;
      12916: inst = 32'd268468224;
      12917: inst = 32'd201346173;
      12918: inst = 32'd203484889;
      12919: inst = 32'd136314880;
      12920: inst = 32'd268468224;
      12921: inst = 32'd201346174;
      12922: inst = 32'd203484857;
      12923: inst = 32'd136314880;
      12924: inst = 32'd268468224;
      12925: inst = 32'd201346175;
      12926: inst = 32'd203484824;
      12927: inst = 32'd136314880;
      12928: inst = 32'd268468224;
      12929: inst = 32'd201346176;
      12930: inst = 32'd203482840;
      12931: inst = 32'd136314880;
      12932: inst = 32'd268468224;
      12933: inst = 32'd201346177;
      12934: inst = 32'd203482807;
      12935: inst = 32'd136314880;
      12936: inst = 32'd268468224;
      12937: inst = 32'd201346178;
      12938: inst = 32'd203482807;
      12939: inst = 32'd136314880;
      12940: inst = 32'd268468224;
      12941: inst = 32'd201346179;
      12942: inst = 32'd203484888;
      12943: inst = 32'd136314880;
      12944: inst = 32'd268468224;
      12945: inst = 32'd201346180;
      12946: inst = 32'd203482775;
      12947: inst = 32'd136314880;
      12948: inst = 32'd268468224;
      12949: inst = 32'd201346181;
      12950: inst = 32'd203484823;
      12951: inst = 32'd136314880;
      12952: inst = 32'd268468224;
      12953: inst = 32'd201346182;
      12954: inst = 32'd203486935;
      12955: inst = 32'd136314880;
      12956: inst = 32'd268468224;
      12957: inst = 32'd201346183;
      12958: inst = 32'd203482774;
      12959: inst = 32'd136314880;
      12960: inst = 32'd268468224;
      12961: inst = 32'd201346184;
      12962: inst = 32'd203484887;
      12963: inst = 32'd136314880;
      12964: inst = 32'd268468224;
      12965: inst = 32'd201346185;
      12966: inst = 32'd203484854;
      12967: inst = 32'd136314880;
      12968: inst = 32'd268468224;
      12969: inst = 32'd201346186;
      12970: inst = 32'd203486901;
      12971: inst = 32'd136314880;
      12972: inst = 32'd268468224;
      12973: inst = 32'd201346187;
      12974: inst = 32'd203484854;
      12975: inst = 32'd136314880;
      12976: inst = 32'd268468224;
      12977: inst = 32'd201346188;
      12978: inst = 32'd203482840;
      12979: inst = 32'd136314880;
      12980: inst = 32'd268468224;
      12981: inst = 32'd201346189;
      12982: inst = 32'd203484855;
      12983: inst = 32'd136314880;
      12984: inst = 32'd268468224;
      12985: inst = 32'd201346190;
      12986: inst = 32'd203488884;
      12987: inst = 32'd136314880;
      12988: inst = 32'd268468224;
      12989: inst = 32'd201346191;
      12990: inst = 32'd203471619;
      12991: inst = 32'd136314880;
      12992: inst = 32'd268468224;
      12993: inst = 32'd201346192;
      12994: inst = 32'd203480005;
      12995: inst = 32'd136314880;
      12996: inst = 32'd268468224;
      12997: inst = 32'd201346193;
      12998: inst = 32'd203480005;
      12999: inst = 32'd136314880;
      13000: inst = 32'd268468224;
      13001: inst = 32'd201346194;
      13002: inst = 32'd203480005;
      13003: inst = 32'd136314880;
      13004: inst = 32'd268468224;
      13005: inst = 32'd201346195;
      13006: inst = 32'd203480005;
      13007: inst = 32'd136314880;
      13008: inst = 32'd268468224;
      13009: inst = 32'd201346196;
      13010: inst = 32'd203480006;
      13011: inst = 32'd136314880;
      13012: inst = 32'd268468224;
      13013: inst = 32'd201346197;
      13014: inst = 32'd203480006;
      13015: inst = 32'd136314880;
      13016: inst = 32'd268468224;
      13017: inst = 32'd201346198;
      13018: inst = 32'd203480006;
      13019: inst = 32'd136314880;
      13020: inst = 32'd268468224;
      13021: inst = 32'd201346199;
      13022: inst = 32'd203480006;
      13023: inst = 32'd136314880;
      13024: inst = 32'd268468224;
      13025: inst = 32'd201346200;
      13026: inst = 32'd203480039;
      13027: inst = 32'd136314880;
      13028: inst = 32'd268468224;
      13029: inst = 32'd201346201;
      13030: inst = 32'd203477958;
      13031: inst = 32'd136314880;
      13032: inst = 32'd268468224;
      13033: inst = 32'd201346202;
      13034: inst = 32'd203480039;
      13035: inst = 32'd136314880;
      13036: inst = 32'd268468224;
      13037: inst = 32'd201346203;
      13038: inst = 32'd203477927;
      13039: inst = 32'd136314880;
      13040: inst = 32'd268468224;
      13041: inst = 32'd201346204;
      13042: inst = 32'd203477991;
      13043: inst = 32'd136314880;
      13044: inst = 32'd268468224;
      13045: inst = 32'd201346205;
      13046: inst = 32'd203473765;
      13047: inst = 32'd136314880;
      13048: inst = 32'd268468224;
      13049: inst = 32'd201346206;
      13050: inst = 32'd203477992;
      13051: inst = 32'd136314880;
      13052: inst = 32'd268468224;
      13053: inst = 32'd201346207;
      13054: inst = 32'd203471652;
      13055: inst = 32'd136314880;
      13056: inst = 32'd268468224;
      13057: inst = 32'd201346208;
      13058: inst = 32'd203482742;
      13059: inst = 32'd136314880;
      13060: inst = 32'd268468224;
      13061: inst = 32'd201346209;
      13062: inst = 32'd203482807;
      13063: inst = 32'd136314880;
      13064: inst = 32'd268468224;
      13065: inst = 32'd201346210;
      13066: inst = 32'd203478549;
      13067: inst = 32'd136314880;
      13068: inst = 32'd268468224;
      13069: inst = 32'd201346211;
      13070: inst = 32'd203465936;
      13071: inst = 32'd136314880;
      13072: inst = 32'd268468224;
      13073: inst = 32'd201346212;
      13074: inst = 32'd203457452;
      13075: inst = 32'd136314880;
      13076: inst = 32'd268468224;
      13077: inst = 32'd201346213;
      13078: inst = 32'd203457485;
      13079: inst = 32'd136314880;
      13080: inst = 32'd268468224;
      13081: inst = 32'd201346214;
      13082: inst = 32'd203457550;
      13083: inst = 32'd136314880;
      13084: inst = 32'd268468224;
      13085: inst = 32'd201346215;
      13086: inst = 32'd203455438;
      13087: inst = 32'd136314880;
      13088: inst = 32'd268468224;
      13089: inst = 32'd201346216;
      13090: inst = 32'd203442760;
      13091: inst = 32'd136314880;
      13092: inst = 32'd268468224;
      13093: inst = 32'd201346217;
      13094: inst = 32'd203480794;
      13095: inst = 32'd136314880;
      13096: inst = 32'd268468224;
      13097: inst = 32'd201346218;
      13098: inst = 32'd203444874;
      13099: inst = 32'd136314880;
      13100: inst = 32'd268468224;
      13101: inst = 32'd201346219;
      13102: inst = 32'd203482908;
      13103: inst = 32'd136314880;
      13104: inst = 32'd268468224;
      13105: inst = 32'd201346220;
      13106: inst = 32'd203442761;
      13107: inst = 32'd136314880;
      13108: inst = 32'd268468224;
      13109: inst = 32'd201346221;
      13110: inst = 32'd203470197;
      13111: inst = 32'd136314880;
      13112: inst = 32'd268468224;
      13113: inst = 32'd201346222;
      13114: inst = 32'd203459600;
      13115: inst = 32'd136314880;
      13116: inst = 32'd268468224;
      13117: inst = 32'd201346223;
      13118: inst = 32'd203457552;
      13119: inst = 32'd136314880;
      13120: inst = 32'd268468224;
      13121: inst = 32'd201346224;
      13122: inst = 32'd203459535;
      13123: inst = 32'd136314880;
      13124: inst = 32'd268468224;
      13125: inst = 32'd201346225;
      13126: inst = 32'd203461647;
      13127: inst = 32'd136314880;
      13128: inst = 32'd268468224;
      13129: inst = 32'd201346226;
      13130: inst = 32'd203461646;
      13131: inst = 32'd136314880;
      13132: inst = 32'd268468224;
      13133: inst = 32'd201346227;
      13134: inst = 32'd203459598;
      13135: inst = 32'd136314880;
      13136: inst = 32'd268468224;
      13137: inst = 32'd201346228;
      13138: inst = 32'd203459566;
      13139: inst = 32'd136314880;
      13140: inst = 32'd268468224;
      13141: inst = 32'd201346229;
      13142: inst = 32'd203461679;
      13143: inst = 32'd136314880;
      13144: inst = 32'd268468224;
      13145: inst = 32'd201346230;
      13146: inst = 32'd203463791;
      13147: inst = 32'd136314880;
      13148: inst = 32'd268468224;
      13149: inst = 32'd201346231;
      13150: inst = 32'd203484919;
      13151: inst = 32'd136314880;
      13152: inst = 32'd268468224;
      13153: inst = 32'd201346232;
      13154: inst = 32'd203484886;
      13155: inst = 32'd136314880;
      13156: inst = 32'd268468224;
      13157: inst = 32'd201346233;
      13158: inst = 32'd203486968;
      13159: inst = 32'd136314880;
      13160: inst = 32'd268468224;
      13161: inst = 32'd201346234;
      13162: inst = 32'd203484856;
      13163: inst = 32'd136314880;
      13164: inst = 32'd268468224;
      13165: inst = 32'd201346235;
      13166: inst = 32'd203484888;
      13167: inst = 32'd136314880;
      13168: inst = 32'd268468224;
      13169: inst = 32'd201346236;
      13170: inst = 32'd203484919;
      13171: inst = 32'd136314880;
      13172: inst = 32'd268468224;
      13173: inst = 32'd201346237;
      13174: inst = 32'd203482806;
      13175: inst = 32'd136314880;
      13176: inst = 32'd268468224;
      13177: inst = 32'd201346238;
      13178: inst = 32'd203482807;
      13179: inst = 32'd136314880;
      13180: inst = 32'd268468224;
      13181: inst = 32'd201346239;
      13182: inst = 32'd203484888;
      13183: inst = 32'd136314880;
      13184: inst = 32'd268468224;
      13185: inst = 32'd201346240;
      13186: inst = 32'd203484823;
      13187: inst = 32'd136314880;
      13188: inst = 32'd268468224;
      13189: inst = 32'd201346241;
      13190: inst = 32'd203484823;
      13191: inst = 32'd136314880;
      13192: inst = 32'd268468224;
      13193: inst = 32'd201346242;
      13194: inst = 32'd203484822;
      13195: inst = 32'd136314880;
      13196: inst = 32'd268468224;
      13197: inst = 32'd201346243;
      13198: inst = 32'd203482774;
      13199: inst = 32'd136314880;
      13200: inst = 32'd268468224;
      13201: inst = 32'd201346244;
      13202: inst = 32'd203482806;
      13203: inst = 32'd136314880;
      13204: inst = 32'd268468224;
      13205: inst = 32'd201346245;
      13206: inst = 32'd203482806;
      13207: inst = 32'd136314880;
      13208: inst = 32'd268468224;
      13209: inst = 32'd201346246;
      13210: inst = 32'd203484887;
      13211: inst = 32'd136314880;
      13212: inst = 32'd268468224;
      13213: inst = 32'd201346247;
      13214: inst = 32'd203484919;
      13215: inst = 32'd136314880;
      13216: inst = 32'd268468224;
      13217: inst = 32'd201346248;
      13218: inst = 32'd203484855;
      13219: inst = 32'd136314880;
      13220: inst = 32'd268468224;
      13221: inst = 32'd201346249;
      13222: inst = 32'd203484823;
      13223: inst = 32'd136314880;
      13224: inst = 32'd268468224;
      13225: inst = 32'd201346250;
      13226: inst = 32'd203484823;
      13227: inst = 32'd136314880;
      13228: inst = 32'd268468224;
      13229: inst = 32'd201346251;
      13230: inst = 32'd203484823;
      13231: inst = 32'd136314880;
      13232: inst = 32'd268468224;
      13233: inst = 32'd201346252;
      13234: inst = 32'd203484855;
      13235: inst = 32'd136314880;
      13236: inst = 32'd268468224;
      13237: inst = 32'd201346253;
      13238: inst = 32'd203482806;
      13239: inst = 32'd136314880;
      13240: inst = 32'd268468224;
      13241: inst = 32'd201346254;
      13242: inst = 32'd203482806;
      13243: inst = 32'd136314880;
      13244: inst = 32'd268468224;
      13245: inst = 32'd201346255;
      13246: inst = 32'd203482806;
      13247: inst = 32'd136314880;
      13248: inst = 32'd268468224;
      13249: inst = 32'd201346256;
      13250: inst = 32'd203482806;
      13251: inst = 32'd136314880;
      13252: inst = 32'd268468224;
      13253: inst = 32'd201346257;
      13254: inst = 32'd203482806;
      13255: inst = 32'd136314880;
      13256: inst = 32'd268468224;
      13257: inst = 32'd201346258;
      13258: inst = 32'd203482806;
      13259: inst = 32'd136314880;
      13260: inst = 32'd268468224;
      13261: inst = 32'd201346259;
      13262: inst = 32'd203484855;
      13263: inst = 32'd136314880;
      13264: inst = 32'd268468224;
      13265: inst = 32'd201346260;
      13266: inst = 32'd203484823;
      13267: inst = 32'd136314880;
      13268: inst = 32'd268468224;
      13269: inst = 32'd201346261;
      13270: inst = 32'd203484823;
      13271: inst = 32'd136314880;
      13272: inst = 32'd268468224;
      13273: inst = 32'd201346262;
      13274: inst = 32'd203484823;
      13275: inst = 32'd136314880;
      13276: inst = 32'd268468224;
      13277: inst = 32'd201346263;
      13278: inst = 32'd203484855;
      13279: inst = 32'd136314880;
      13280: inst = 32'd268468224;
      13281: inst = 32'd201346264;
      13282: inst = 32'd203484919;
      13283: inst = 32'd136314880;
      13284: inst = 32'd268468224;
      13285: inst = 32'd201346265;
      13286: inst = 32'd203484887;
      13287: inst = 32'd136314880;
      13288: inst = 32'd268468224;
      13289: inst = 32'd201346266;
      13290: inst = 32'd203482806;
      13291: inst = 32'd136314880;
      13292: inst = 32'd268468224;
      13293: inst = 32'd201346267;
      13294: inst = 32'd203482806;
      13295: inst = 32'd136314880;
      13296: inst = 32'd268468224;
      13297: inst = 32'd201346268;
      13298: inst = 32'd203482774;
      13299: inst = 32'd136314880;
      13300: inst = 32'd268468224;
      13301: inst = 32'd201346269;
      13302: inst = 32'd203484822;
      13303: inst = 32'd136314880;
      13304: inst = 32'd268468224;
      13305: inst = 32'd201346270;
      13306: inst = 32'd203484823;
      13307: inst = 32'd136314880;
      13308: inst = 32'd268468224;
      13309: inst = 32'd201346271;
      13310: inst = 32'd203484823;
      13311: inst = 32'd136314880;
      13312: inst = 32'd268468224;
      13313: inst = 32'd201346272;
      13314: inst = 32'd203482872;
      13315: inst = 32'd136314880;
      13316: inst = 32'd268468224;
      13317: inst = 32'd201346273;
      13318: inst = 32'd203482807;
      13319: inst = 32'd136314880;
      13320: inst = 32'd268468224;
      13321: inst = 32'd201346274;
      13322: inst = 32'd203482775;
      13323: inst = 32'd136314880;
      13324: inst = 32'd268468224;
      13325: inst = 32'd201346275;
      13326: inst = 32'd203484920;
      13327: inst = 32'd136314880;
      13328: inst = 32'd268468224;
      13329: inst = 32'd201346276;
      13330: inst = 32'd203484888;
      13331: inst = 32'd136314880;
      13332: inst = 32'd268468224;
      13333: inst = 32'd201346277;
      13334: inst = 32'd203486935;
      13335: inst = 32'd136314880;
      13336: inst = 32'd268468224;
      13337: inst = 32'd201346278;
      13338: inst = 32'd203488983;
      13339: inst = 32'd136314880;
      13340: inst = 32'd268468224;
      13341: inst = 32'd201346279;
      13342: inst = 32'd203484854;
      13343: inst = 32'd136314880;
      13344: inst = 32'd268468224;
      13345: inst = 32'd201346280;
      13346: inst = 32'd203484887;
      13347: inst = 32'd136314880;
      13348: inst = 32'd268468224;
      13349: inst = 32'd201346281;
      13350: inst = 32'd203484854;
      13351: inst = 32'd136314880;
      13352: inst = 32'd268468224;
      13353: inst = 32'd201346282;
      13354: inst = 32'd203486901;
      13355: inst = 32'd136314880;
      13356: inst = 32'd268468224;
      13357: inst = 32'd201346283;
      13358: inst = 32'd203484854;
      13359: inst = 32'd136314880;
      13360: inst = 32'd268468224;
      13361: inst = 32'd201346284;
      13362: inst = 32'd203482840;
      13363: inst = 32'd136314880;
      13364: inst = 32'd268468224;
      13365: inst = 32'd201346285;
      13366: inst = 32'd203484855;
      13367: inst = 32'd136314880;
      13368: inst = 32'd268468224;
      13369: inst = 32'd201346286;
      13370: inst = 32'd203488884;
      13371: inst = 32'd136314880;
      13372: inst = 32'd268468224;
      13373: inst = 32'd201346287;
      13374: inst = 32'd203471619;
      13375: inst = 32'd136314880;
      13376: inst = 32'd268468224;
      13377: inst = 32'd201346288;
      13378: inst = 32'd203480005;
      13379: inst = 32'd136314880;
      13380: inst = 32'd268468224;
      13381: inst = 32'd201346289;
      13382: inst = 32'd203480005;
      13383: inst = 32'd136314880;
      13384: inst = 32'd268468224;
      13385: inst = 32'd201346290;
      13386: inst = 32'd203480005;
      13387: inst = 32'd136314880;
      13388: inst = 32'd268468224;
      13389: inst = 32'd201346291;
      13390: inst = 32'd203480005;
      13391: inst = 32'd136314880;
      13392: inst = 32'd268468224;
      13393: inst = 32'd201346292;
      13394: inst = 32'd203480006;
      13395: inst = 32'd136314880;
      13396: inst = 32'd268468224;
      13397: inst = 32'd201346293;
      13398: inst = 32'd203480006;
      13399: inst = 32'd136314880;
      13400: inst = 32'd268468224;
      13401: inst = 32'd201346294;
      13402: inst = 32'd203480006;
      13403: inst = 32'd136314880;
      13404: inst = 32'd268468224;
      13405: inst = 32'd201346295;
      13406: inst = 32'd203480006;
      13407: inst = 32'd136314880;
      13408: inst = 32'd268468224;
      13409: inst = 32'd201346296;
      13410: inst = 32'd203480039;
      13411: inst = 32'd136314880;
      13412: inst = 32'd268468224;
      13413: inst = 32'd201346297;
      13414: inst = 32'd203477926;
      13415: inst = 32'd136314880;
      13416: inst = 32'd268468224;
      13417: inst = 32'd201346298;
      13418: inst = 32'd203477958;
      13419: inst = 32'd136314880;
      13420: inst = 32'd268468224;
      13421: inst = 32'd201346299;
      13422: inst = 32'd203486411;
      13423: inst = 32'd136314880;
      13424: inst = 32'd268468224;
      13425: inst = 32'd201346300;
      13426: inst = 32'd203477926;
      13427: inst = 32'd136314880;
      13428: inst = 32'd268468224;
      13429: inst = 32'd201346301;
      13430: inst = 32'd203477927;
      13431: inst = 32'd136314880;
      13432: inst = 32'd268468224;
      13433: inst = 32'd201346302;
      13434: inst = 32'd203477959;
      13435: inst = 32'd136314880;
      13436: inst = 32'd268468224;
      13437: inst = 32'd201346303;
      13438: inst = 32'd203471620;
      13439: inst = 32'd136314880;
      13440: inst = 32'd268468224;
      13441: inst = 32'd201346304;
      13442: inst = 32'd203476469;
      13443: inst = 32'd136314880;
      13444: inst = 32'd268468224;
      13445: inst = 32'd201346305;
      13446: inst = 32'd203465937;
      13447: inst = 32'd136314880;
      13448: inst = 32'd268468224;
      13449: inst = 32'd201346306;
      13450: inst = 32'd203457485;
      13451: inst = 32'd136314880;
      13452: inst = 32'd268468224;
      13453: inst = 32'd201346307;
      13454: inst = 32'd203457485;
      13455: inst = 32'd136314880;
      13456: inst = 32'd268468224;
      13457: inst = 32'd201346308;
      13458: inst = 32'd203457486;
      13459: inst = 32'd136314880;
      13460: inst = 32'd268468224;
      13461: inst = 32'd201346309;
      13462: inst = 32'd203457486;
      13463: inst = 32'd136314880;
      13464: inst = 32'd268468224;
      13465: inst = 32'd201346310;
      13466: inst = 32'd203455471;
      13467: inst = 32'd136314880;
      13468: inst = 32'd268468224;
      13469: inst = 32'd201346311;
      13470: inst = 32'd203455438;
      13471: inst = 32'd136314880;
      13472: inst = 32'd268468224;
      13473: inst = 32'd201346312;
      13474: inst = 32'd203455471;
      13475: inst = 32'd136314880;
      13476: inst = 32'd268468224;
      13477: inst = 32'd201346313;
      13478: inst = 32'd203455471;
      13479: inst = 32'd136314880;
      13480: inst = 32'd268468224;
      13481: inst = 32'd201346314;
      13482: inst = 32'd203455472;
      13483: inst = 32'd136314880;
      13484: inst = 32'd268468224;
      13485: inst = 32'd201346315;
      13486: inst = 32'd203455439;
      13487: inst = 32'd136314880;
      13488: inst = 32'd268468224;
      13489: inst = 32'd201346316;
      13490: inst = 32'd203455439;
      13491: inst = 32'd136314880;
      13492: inst = 32'd268468224;
      13493: inst = 32'd201346317;
      13494: inst = 32'd203455439;
      13495: inst = 32'd136314880;
      13496: inst = 32'd268468224;
      13497: inst = 32'd201346318;
      13498: inst = 32'd203455406;
      13499: inst = 32'd136314880;
      13500: inst = 32'd268468224;
      13501: inst = 32'd201346319;
      13502: inst = 32'd203457519;
      13503: inst = 32'd136314880;
      13504: inst = 32'd268468224;
      13505: inst = 32'd201346320;
      13506: inst = 32'd203459569;
      13507: inst = 32'd136314880;
      13508: inst = 32'd268468224;
      13509: inst = 32'd201346321;
      13510: inst = 32'd203457488;
      13511: inst = 32'd136314880;
      13512: inst = 32'd268468224;
      13513: inst = 32'd201346322;
      13514: inst = 32'd203455406;
      13515: inst = 32'd136314880;
      13516: inst = 32'd268468224;
      13517: inst = 32'd201346323;
      13518: inst = 32'd203455406;
      13519: inst = 32'd136314880;
      13520: inst = 32'd268468224;
      13521: inst = 32'd201346324;
      13522: inst = 32'd203457519;
      13523: inst = 32'd136314880;
      13524: inst = 32'd268468224;
      13525: inst = 32'd201346325;
      13526: inst = 32'd203457519;
      13527: inst = 32'd136314880;
      13528: inst = 32'd268468224;
      13529: inst = 32'd201346326;
      13530: inst = 32'd203457452;
      13531: inst = 32'd136314880;
      13532: inst = 32'd268468224;
      13533: inst = 32'd201346327;
      13534: inst = 32'd203482806;
      13535: inst = 32'd136314880;
      13536: inst = 32'd268468224;
      13537: inst = 32'd201346328;
      13538: inst = 32'd203484886;
      13539: inst = 32'd136314880;
      13540: inst = 32'd268468224;
      13541: inst = 32'd201346329;
      13542: inst = 32'd203484854;
      13543: inst = 32'd136314880;
      13544: inst = 32'd268468224;
      13545: inst = 32'd201346330;
      13546: inst = 32'd203482742;
      13547: inst = 32'd136314880;
      13548: inst = 32'd268468224;
      13549: inst = 32'd201346331;
      13550: inst = 32'd203484822;
      13551: inst = 32'd136314880;
      13552: inst = 32'd268468224;
      13553: inst = 32'd201346332;
      13554: inst = 32'd203486933;
      13555: inst = 32'd136314880;
      13556: inst = 32'd268468224;
      13557: inst = 32'd201346333;
      13558: inst = 32'd203484852;
      13559: inst = 32'd136314880;
      13560: inst = 32'd268468224;
      13561: inst = 32'd201346334;
      13562: inst = 32'd203484885;
      13563: inst = 32'd136314880;
      13564: inst = 32'd268468224;
      13565: inst = 32'd201346335;
      13566: inst = 32'd203484854;
      13567: inst = 32'd136314880;
      13568: inst = 32'd268468224;
      13569: inst = 32'd201346336;
      13570: inst = 32'd203486902;
      13571: inst = 32'd136314880;
      13572: inst = 32'd268468224;
      13573: inst = 32'd201346337;
      13574: inst = 32'd203486902;
      13575: inst = 32'd136314880;
      13576: inst = 32'd268468224;
      13577: inst = 32'd201346338;
      13578: inst = 32'd203486901;
      13579: inst = 32'd136314880;
      13580: inst = 32'd268468224;
      13581: inst = 32'd201346339;
      13582: inst = 32'd203484885;
      13583: inst = 32'd136314880;
      13584: inst = 32'd268468224;
      13585: inst = 32'd201346340;
      13586: inst = 32'd203484885;
      13587: inst = 32'd136314880;
      13588: inst = 32'd268468224;
      13589: inst = 32'd201346341;
      13590: inst = 32'd203484853;
      13591: inst = 32'd136314880;
      13592: inst = 32'd268468224;
      13593: inst = 32'd201346342;
      13594: inst = 32'd203484821;
      13595: inst = 32'd136314880;
      13596: inst = 32'd268468224;
      13597: inst = 32'd201346343;
      13598: inst = 32'd203482741;
      13599: inst = 32'd136314880;
      13600: inst = 32'd268468224;
      13601: inst = 32'd201346344;
      13602: inst = 32'd203486902;
      13603: inst = 32'd136314880;
      13604: inst = 32'd268468224;
      13605: inst = 32'd201346345;
      13606: inst = 32'd203486902;
      13607: inst = 32'd136314880;
      13608: inst = 32'd268468224;
      13609: inst = 32'd201346346;
      13610: inst = 32'd203486902;
      13611: inst = 32'd136314880;
      13612: inst = 32'd268468224;
      13613: inst = 32'd201346347;
      13614: inst = 32'd203486902;
      13615: inst = 32'd136314880;
      13616: inst = 32'd268468224;
      13617: inst = 32'd201346348;
      13618: inst = 32'd203486902;
      13619: inst = 32'd136314880;
      13620: inst = 32'd268468224;
      13621: inst = 32'd201346349;
      13622: inst = 32'd203486902;
      13623: inst = 32'd136314880;
      13624: inst = 32'd268468224;
      13625: inst = 32'd201346350;
      13626: inst = 32'd203484854;
      13627: inst = 32'd136314880;
      13628: inst = 32'd268468224;
      13629: inst = 32'd201346351;
      13630: inst = 32'd203484886;
      13631: inst = 32'd136314880;
      13632: inst = 32'd268468224;
      13633: inst = 32'd201346352;
      13634: inst = 32'd203484886;
      13635: inst = 32'd136314880;
      13636: inst = 32'd268468224;
      13637: inst = 32'd201346353;
      13638: inst = 32'd203484854;
      13639: inst = 32'd136314880;
      13640: inst = 32'd268468224;
      13641: inst = 32'd201346354;
      13642: inst = 32'd203486902;
      13643: inst = 32'd136314880;
      13644: inst = 32'd268468224;
      13645: inst = 32'd201346355;
      13646: inst = 32'd203486902;
      13647: inst = 32'd136314880;
      13648: inst = 32'd268468224;
      13649: inst = 32'd201346356;
      13650: inst = 32'd203486902;
      13651: inst = 32'd136314880;
      13652: inst = 32'd268468224;
      13653: inst = 32'd201346357;
      13654: inst = 32'd203486902;
      13655: inst = 32'd136314880;
      13656: inst = 32'd268468224;
      13657: inst = 32'd201346358;
      13658: inst = 32'd203486902;
      13659: inst = 32'd136314880;
      13660: inst = 32'd268468224;
      13661: inst = 32'd201346359;
      13662: inst = 32'd203486902;
      13663: inst = 32'd136314880;
      13664: inst = 32'd268468224;
      13665: inst = 32'd201346360;
      13666: inst = 32'd203482741;
      13667: inst = 32'd136314880;
      13668: inst = 32'd268468224;
      13669: inst = 32'd201346361;
      13670: inst = 32'd203484821;
      13671: inst = 32'd136314880;
      13672: inst = 32'd268468224;
      13673: inst = 32'd201346362;
      13674: inst = 32'd203484853;
      13675: inst = 32'd136314880;
      13676: inst = 32'd268468224;
      13677: inst = 32'd201346363;
      13678: inst = 32'd203484885;
      13679: inst = 32'd136314880;
      13680: inst = 32'd268468224;
      13681: inst = 32'd201346364;
      13682: inst = 32'd203484885;
      13683: inst = 32'd136314880;
      13684: inst = 32'd268468224;
      13685: inst = 32'd201346365;
      13686: inst = 32'd203486901;
      13687: inst = 32'd136314880;
      13688: inst = 32'd268468224;
      13689: inst = 32'd201346366;
      13690: inst = 32'd203486902;
      13691: inst = 32'd136314880;
      13692: inst = 32'd268468224;
      13693: inst = 32'd201346367;
      13694: inst = 32'd203486902;
      13695: inst = 32'd136314880;
      13696: inst = 32'd268468224;
      13697: inst = 32'd201346368;
      13698: inst = 32'd203482840;
      13699: inst = 32'd136314880;
      13700: inst = 32'd268468224;
      13701: inst = 32'd201346369;
      13702: inst = 32'd203484887;
      13703: inst = 32'd136314880;
      13704: inst = 32'd268468224;
      13705: inst = 32'd201346370;
      13706: inst = 32'd203484854;
      13707: inst = 32'd136314880;
      13708: inst = 32'd268468224;
      13709: inst = 32'd201346371;
      13710: inst = 32'd203484887;
      13711: inst = 32'd136314880;
      13712: inst = 32'd268468224;
      13713: inst = 32'd201346372;
      13714: inst = 32'd203482807;
      13715: inst = 32'd136314880;
      13716: inst = 32'd268468224;
      13717: inst = 32'd201346373;
      13718: inst = 32'd203482742;
      13719: inst = 32'd136314880;
      13720: inst = 32'd268468224;
      13721: inst = 32'd201346374;
      13722: inst = 32'd203486870;
      13723: inst = 32'd136314880;
      13724: inst = 32'd268468224;
      13725: inst = 32'd201346375;
      13726: inst = 32'd203484854;
      13727: inst = 32'd136314880;
      13728: inst = 32'd268468224;
      13729: inst = 32'd201346376;
      13730: inst = 32'd203484887;
      13731: inst = 32'd136314880;
      13732: inst = 32'd268468224;
      13733: inst = 32'd201346377;
      13734: inst = 32'd203484854;
      13735: inst = 32'd136314880;
      13736: inst = 32'd268468224;
      13737: inst = 32'd201346378;
      13738: inst = 32'd203486901;
      13739: inst = 32'd136314880;
      13740: inst = 32'd268468224;
      13741: inst = 32'd201346379;
      13742: inst = 32'd203484854;
      13743: inst = 32'd136314880;
      13744: inst = 32'd268468224;
      13745: inst = 32'd201346380;
      13746: inst = 32'd203482840;
      13747: inst = 32'd136314880;
      13748: inst = 32'd268468224;
      13749: inst = 32'd201346381;
      13750: inst = 32'd203484855;
      13751: inst = 32'd136314880;
      13752: inst = 32'd268468224;
      13753: inst = 32'd201346382;
      13754: inst = 32'd203488884;
      13755: inst = 32'd136314880;
      13756: inst = 32'd268468224;
      13757: inst = 32'd201346383;
      13758: inst = 32'd203471619;
      13759: inst = 32'd136314880;
      13760: inst = 32'd268468224;
      13761: inst = 32'd201346384;
      13762: inst = 32'd203480005;
      13763: inst = 32'd136314880;
      13764: inst = 32'd268468224;
      13765: inst = 32'd201346385;
      13766: inst = 32'd203480005;
      13767: inst = 32'd136314880;
      13768: inst = 32'd268468224;
      13769: inst = 32'd201346386;
      13770: inst = 32'd203480005;
      13771: inst = 32'd136314880;
      13772: inst = 32'd268468224;
      13773: inst = 32'd201346387;
      13774: inst = 32'd203480005;
      13775: inst = 32'd136314880;
      13776: inst = 32'd268468224;
      13777: inst = 32'd201346388;
      13778: inst = 32'd203480006;
      13779: inst = 32'd136314880;
      13780: inst = 32'd268468224;
      13781: inst = 32'd201346389;
      13782: inst = 32'd203480006;
      13783: inst = 32'd136314880;
      13784: inst = 32'd268468224;
      13785: inst = 32'd201346390;
      13786: inst = 32'd203480006;
      13787: inst = 32'd136314880;
      13788: inst = 32'd268468224;
      13789: inst = 32'd201346391;
      13790: inst = 32'd203480006;
      13791: inst = 32'd136314880;
      13792: inst = 32'd268468224;
      13793: inst = 32'd201346392;
      13794: inst = 32'd203479974;
      13795: inst = 32'd136314880;
      13796: inst = 32'd268468224;
      13797: inst = 32'd201346393;
      13798: inst = 32'd203480006;
      13799: inst = 32'd136314880;
      13800: inst = 32'd268468224;
      13801: inst = 32'd201346394;
      13802: inst = 32'd203480006;
      13803: inst = 32'd136314880;
      13804: inst = 32'd268468224;
      13805: inst = 32'd201346395;
      13806: inst = 32'd203488556;
      13807: inst = 32'd136314880;
      13808: inst = 32'd268468224;
      13809: inst = 32'd201346396;
      13810: inst = 32'd203477958;
      13811: inst = 32'd136314880;
      13812: inst = 32'd268468224;
      13813: inst = 32'd201346397;
      13814: inst = 32'd203480071;
      13815: inst = 32'd136314880;
      13816: inst = 32'd268468224;
      13817: inst = 32'd201346398;
      13818: inst = 32'd203477926;
      13819: inst = 32'd136314880;
      13820: inst = 32'd268468224;
      13821: inst = 32'd201346399;
      13822: inst = 32'd203471587;
      13823: inst = 32'd136314880;
      13824: inst = 32'd268468224;
      13825: inst = 32'd201346400;
      13826: inst = 32'd203461744;
      13827: inst = 32'd136314880;
      13828: inst = 32'd268468224;
      13829: inst = 32'd201346401;
      13830: inst = 32'd203461712;
      13831: inst = 32'd136314880;
      13832: inst = 32'd268468224;
      13833: inst = 32'd201346402;
      13834: inst = 32'd203459664;
      13835: inst = 32'd136314880;
      13836: inst = 32'd268468224;
      13837: inst = 32'd201346403;
      13838: inst = 32'd203461777;
      13839: inst = 32'd136314880;
      13840: inst = 32'd268468224;
      13841: inst = 32'd201346404;
      13842: inst = 32'd203461745;
      13843: inst = 32'd136314880;
      13844: inst = 32'd268468224;
      13845: inst = 32'd201346405;
      13846: inst = 32'd203457584;
      13847: inst = 32'd136314880;
      13848: inst = 32'd268468224;
      13849: inst = 32'd201346406;
      13850: inst = 32'd203459697;
      13851: inst = 32'd136314880;
      13852: inst = 32'd268468224;
      13853: inst = 32'd201346407;
      13854: inst = 32'd203459730;
      13855: inst = 32'd136314880;
      13856: inst = 32'd268468224;
      13857: inst = 32'd201346408;
      13858: inst = 32'd203459730;
      13859: inst = 32'd136314880;
      13860: inst = 32'd268468224;
      13861: inst = 32'd201346409;
      13862: inst = 32'd203459698;
      13863: inst = 32'd136314880;
      13864: inst = 32'd268468224;
      13865: inst = 32'd201346410;
      13866: inst = 32'd203457617;
      13867: inst = 32'd136314880;
      13868: inst = 32'd268468224;
      13869: inst = 32'd201346411;
      13870: inst = 32'd203459698;
      13871: inst = 32'd136314880;
      13872: inst = 32'd268468224;
      13873: inst = 32'd201346412;
      13874: inst = 32'd203459698;
      13875: inst = 32'd136314880;
      13876: inst = 32'd268468224;
      13877: inst = 32'd201346413;
      13878: inst = 32'd203461810;
      13879: inst = 32'd136314880;
      13880: inst = 32'd268468224;
      13881: inst = 32'd201346414;
      13882: inst = 32'd203457585;
      13883: inst = 32'd136314880;
      13884: inst = 32'd268468224;
      13885: inst = 32'd201346415;
      13886: inst = 32'd203461778;
      13887: inst = 32'd136314880;
      13888: inst = 32'd268468224;
      13889: inst = 32'd201346416;
      13890: inst = 32'd203459635;
      13891: inst = 32'd136314880;
      13892: inst = 32'd268468224;
      13893: inst = 32'd201346417;
      13894: inst = 32'd203459634;
      13895: inst = 32'd136314880;
      13896: inst = 32'd268468224;
      13897: inst = 32'd201346418;
      13898: inst = 32'd203459665;
      13899: inst = 32'd136314880;
      13900: inst = 32'd268468224;
      13901: inst = 32'd201346419;
      13902: inst = 32'd203461778;
      13903: inst = 32'd136314880;
      13904: inst = 32'd268468224;
      13905: inst = 32'd201346420;
      13906: inst = 32'd203459666;
      13907: inst = 32'd136314880;
      13908: inst = 32'd268468224;
      13909: inst = 32'd201346421;
      13910: inst = 32'd203457487;
      13911: inst = 32'd136314880;
      13912: inst = 32'd268468224;
      13913: inst = 32'd201346422;
      13914: inst = 32'd203453259;
      13915: inst = 32'd136314880;
      13916: inst = 32'd268468224;
      13917: inst = 32'd201346423;
      13918: inst = 32'd203482807;
      13919: inst = 32'd136314880;
      13920: inst = 32'd268468224;
      13921: inst = 32'd201346424;
      13922: inst = 32'd203484886;
      13923: inst = 32'd136314880;
      13924: inst = 32'd268468224;
      13925: inst = 32'd201346425;
      13926: inst = 32'd203484854;
      13927: inst = 32'd136314880;
      13928: inst = 32'd268468224;
      13929: inst = 32'd201346426;
      13930: inst = 32'd203484822;
      13931: inst = 32'd136314880;
      13932: inst = 32'd268468224;
      13933: inst = 32'd201346427;
      13934: inst = 32'd203486934;
      13935: inst = 32'd136314880;
      13936: inst = 32'd268468224;
      13937: inst = 32'd201346428;
      13938: inst = 32'd203486965;
      13939: inst = 32'd136314880;
      13940: inst = 32'd268468224;
      13941: inst = 32'd201346429;
      13942: inst = 32'd203486932;
      13943: inst = 32'd136314880;
      13944: inst = 32'd268468224;
      13945: inst = 32'd201346430;
      13946: inst = 32'd203486933;
      13947: inst = 32'd136314880;
      13948: inst = 32'd268468224;
      13949: inst = 32'd201346431;
      13950: inst = 32'd203484822;
      13951: inst = 32'd136314880;
      13952: inst = 32'd268468224;
      13953: inst = 32'd201346432;
      13954: inst = 32'd203486901;
      13955: inst = 32'd136314880;
      13956: inst = 32'd268468224;
      13957: inst = 32'd201346433;
      13958: inst = 32'd203484821;
      13959: inst = 32'd136314880;
      13960: inst = 32'd268468224;
      13961: inst = 32'd201346434;
      13962: inst = 32'd203484853;
      13963: inst = 32'd136314880;
      13964: inst = 32'd268468224;
      13965: inst = 32'd201346435;
      13966: inst = 32'd203484853;
      13967: inst = 32'd136314880;
      13968: inst = 32'd268468224;
      13969: inst = 32'd201346436;
      13970: inst = 32'd203486934;
      13971: inst = 32'd136314880;
      13972: inst = 32'd268468224;
      13973: inst = 32'd201346437;
      13974: inst = 32'd203486966;
      13975: inst = 32'd136314880;
      13976: inst = 32'd268468224;
      13977: inst = 32'd201346438;
      13978: inst = 32'd203486934;
      13979: inst = 32'd136314880;
      13980: inst = 32'd268468224;
      13981: inst = 32'd201346439;
      13982: inst = 32'd203486934;
      13983: inst = 32'd136314880;
      13984: inst = 32'd268468224;
      13985: inst = 32'd201346440;
      13986: inst = 32'd203486869;
      13987: inst = 32'd136314880;
      13988: inst = 32'd268468224;
      13989: inst = 32'd201346441;
      13990: inst = 32'd203486869;
      13991: inst = 32'd136314880;
      13992: inst = 32'd268468224;
      13993: inst = 32'd201346442;
      13994: inst = 32'd203486869;
      13995: inst = 32'd136314880;
      13996: inst = 32'd268468224;
      13997: inst = 32'd201346443;
      13998: inst = 32'd203486869;
      13999: inst = 32'd136314880;
      14000: inst = 32'd268468224;
      14001: inst = 32'd201346444;
      14002: inst = 32'd203486869;
      14003: inst = 32'd136314880;
      14004: inst = 32'd268468224;
      14005: inst = 32'd201346445;
      14006: inst = 32'd203486869;
      14007: inst = 32'd136314880;
      14008: inst = 32'd268468224;
      14009: inst = 32'd201346446;
      14010: inst = 32'd203486901;
      14011: inst = 32'd136314880;
      14012: inst = 32'd268468224;
      14013: inst = 32'd201346447;
      14014: inst = 32'd203486901;
      14015: inst = 32'd136314880;
      14016: inst = 32'd268468224;
      14017: inst = 32'd201346448;
      14018: inst = 32'd203486901;
      14019: inst = 32'd136314880;
      14020: inst = 32'd268468224;
      14021: inst = 32'd201346449;
      14022: inst = 32'd203486901;
      14023: inst = 32'd136314880;
      14024: inst = 32'd268468224;
      14025: inst = 32'd201346450;
      14026: inst = 32'd203486869;
      14027: inst = 32'd136314880;
      14028: inst = 32'd268468224;
      14029: inst = 32'd201346451;
      14030: inst = 32'd203486869;
      14031: inst = 32'd136314880;
      14032: inst = 32'd268468224;
      14033: inst = 32'd201346452;
      14034: inst = 32'd203486869;
      14035: inst = 32'd136314880;
      14036: inst = 32'd268468224;
      14037: inst = 32'd201346453;
      14038: inst = 32'd203486869;
      14039: inst = 32'd136314880;
      14040: inst = 32'd268468224;
      14041: inst = 32'd201346454;
      14042: inst = 32'd203486869;
      14043: inst = 32'd136314880;
      14044: inst = 32'd268468224;
      14045: inst = 32'd201346455;
      14046: inst = 32'd203486869;
      14047: inst = 32'd136314880;
      14048: inst = 32'd268468224;
      14049: inst = 32'd201346456;
      14050: inst = 32'd203486934;
      14051: inst = 32'd136314880;
      14052: inst = 32'd268468224;
      14053: inst = 32'd201346457;
      14054: inst = 32'd203486934;
      14055: inst = 32'd136314880;
      14056: inst = 32'd268468224;
      14057: inst = 32'd201346458;
      14058: inst = 32'd203486966;
      14059: inst = 32'd136314880;
      14060: inst = 32'd268468224;
      14061: inst = 32'd201346459;
      14062: inst = 32'd203486934;
      14063: inst = 32'd136314880;
      14064: inst = 32'd268468224;
      14065: inst = 32'd201346460;
      14066: inst = 32'd203484853;
      14067: inst = 32'd136314880;
      14068: inst = 32'd268468224;
      14069: inst = 32'd201346461;
      14070: inst = 32'd203484853;
      14071: inst = 32'd136314880;
      14072: inst = 32'd268468224;
      14073: inst = 32'd201346462;
      14074: inst = 32'd203484821;
      14075: inst = 32'd136314880;
      14076: inst = 32'd268468224;
      14077: inst = 32'd201346463;
      14078: inst = 32'd203486901;
      14079: inst = 32'd136314880;
      14080: inst = 32'd268468224;
      14081: inst = 32'd201346464;
      14082: inst = 32'd203482807;
      14083: inst = 32'd136314880;
      14084: inst = 32'd268468224;
      14085: inst = 32'd201346465;
      14086: inst = 32'd203484887;
      14087: inst = 32'd136314880;
      14088: inst = 32'd268468224;
      14089: inst = 32'd201346466;
      14090: inst = 32'd203484855;
      14091: inst = 32'd136314880;
      14092: inst = 32'd268468224;
      14093: inst = 32'd201346467;
      14094: inst = 32'd203484888;
      14095: inst = 32'd136314880;
      14096: inst = 32'd268468224;
      14097: inst = 32'd201346468;
      14098: inst = 32'd203484888;
      14099: inst = 32'd136314880;
      14100: inst = 32'd268468224;
      14101: inst = 32'd201346469;
      14102: inst = 32'd203484822;
      14103: inst = 32'd136314880;
      14104: inst = 32'd268468224;
      14105: inst = 32'd201346470;
      14106: inst = 32'd203486902;
      14107: inst = 32'd136314880;
      14108: inst = 32'd268468224;
      14109: inst = 32'd201346471;
      14110: inst = 32'd203484854;
      14111: inst = 32'd136314880;
      14112: inst = 32'd268468224;
      14113: inst = 32'd201346472;
      14114: inst = 32'd203484887;
      14115: inst = 32'd136314880;
      14116: inst = 32'd268468224;
      14117: inst = 32'd201346473;
      14118: inst = 32'd203484854;
      14119: inst = 32'd136314880;
      14120: inst = 32'd268468224;
      14121: inst = 32'd201346474;
      14122: inst = 32'd203486901;
      14123: inst = 32'd136314880;
      14124: inst = 32'd268468224;
      14125: inst = 32'd201346475;
      14126: inst = 32'd203484854;
      14127: inst = 32'd136314880;
      14128: inst = 32'd268468224;
      14129: inst = 32'd201346476;
      14130: inst = 32'd203482840;
      14131: inst = 32'd136314880;
      14132: inst = 32'd268468224;
      14133: inst = 32'd201346477;
      14134: inst = 32'd203484856;
      14135: inst = 32'd136314880;
      14136: inst = 32'd268468224;
      14137: inst = 32'd201346478;
      14138: inst = 32'd203488884;
      14139: inst = 32'd136314880;
      14140: inst = 32'd268468224;
      14141: inst = 32'd201346479;
      14142: inst = 32'd203471619;
      14143: inst = 32'd136314880;
      14144: inst = 32'd268468224;
      14145: inst = 32'd201346480;
      14146: inst = 32'd203480005;
      14147: inst = 32'd136314880;
      14148: inst = 32'd268468224;
      14149: inst = 32'd201346481;
      14150: inst = 32'd203480005;
      14151: inst = 32'd136314880;
      14152: inst = 32'd268468224;
      14153: inst = 32'd201346482;
      14154: inst = 32'd203480005;
      14155: inst = 32'd136314880;
      14156: inst = 32'd268468224;
      14157: inst = 32'd201346483;
      14158: inst = 32'd203480005;
      14159: inst = 32'd136314880;
      14160: inst = 32'd268468224;
      14161: inst = 32'd201346484;
      14162: inst = 32'd203480006;
      14163: inst = 32'd136314880;
      14164: inst = 32'd268468224;
      14165: inst = 32'd201346485;
      14166: inst = 32'd203480006;
      14167: inst = 32'd136314880;
      14168: inst = 32'd268468224;
      14169: inst = 32'd201346486;
      14170: inst = 32'd203480006;
      14171: inst = 32'd136314880;
      14172: inst = 32'd268468224;
      14173: inst = 32'd201346487;
      14174: inst = 32'd203480006;
      14175: inst = 32'd136314880;
      14176: inst = 32'd268468224;
      14177: inst = 32'd201346488;
      14178: inst = 32'd203480006;
      14179: inst = 32'd136314880;
      14180: inst = 32'd268468224;
      14181: inst = 32'd201346489;
      14182: inst = 32'd203480006;
      14183: inst = 32'd136314880;
      14184: inst = 32'd268468224;
      14185: inst = 32'd201346490;
      14186: inst = 32'd203480039;
      14187: inst = 32'd136314880;
      14188: inst = 32'd268468224;
      14189: inst = 32'd201346491;
      14190: inst = 32'd203480039;
      14191: inst = 32'd136314880;
      14192: inst = 32'd268468224;
      14193: inst = 32'd201346492;
      14194: inst = 32'd203480039;
      14195: inst = 32'd136314880;
      14196: inst = 32'd268468224;
      14197: inst = 32'd201346493;
      14198: inst = 32'd203477893;
      14199: inst = 32'd136314880;
      14200: inst = 32'd268468224;
      14201: inst = 32'd201346494;
      14202: inst = 32'd203480039;
      14203: inst = 32'd136314880;
      14204: inst = 32'd268468224;
      14205: inst = 32'd201346495;
      14206: inst = 32'd203471587;
      14207: inst = 32'd136314880;
      14208: inst = 32'd268468224;
      14209: inst = 32'd201346496;
      14210: inst = 32'd203459665;
      14211: inst = 32'd136314880;
      14212: inst = 32'd268468224;
      14213: inst = 32'd201346497;
      14214: inst = 32'd203472342;
      14215: inst = 32'd136314880;
      14216: inst = 32'd268468224;
      14217: inst = 32'd201346498;
      14218: inst = 32'd203474455;
      14219: inst = 32'd136314880;
      14220: inst = 32'd268468224;
      14221: inst = 32'd201346499;
      14222: inst = 32'd203472343;
      14223: inst = 32'd136314880;
      14224: inst = 32'd268468224;
      14225: inst = 32'd201346500;
      14226: inst = 32'd203470295;
      14227: inst = 32'd136314880;
      14228: inst = 32'd268468224;
      14229: inst = 32'd201346501;
      14230: inst = 32'd203472375;
      14231: inst = 32'd136314880;
      14232: inst = 32'd268468224;
      14233: inst = 32'd201346502;
      14234: inst = 32'd203474489;
      14235: inst = 32'd136314880;
      14236: inst = 32'd268468224;
      14237: inst = 32'd201346503;
      14238: inst = 32'd203468215;
      14239: inst = 32'd136314880;
      14240: inst = 32'd268468224;
      14241: inst = 32'd201346504;
      14242: inst = 32'd203470295;
      14243: inst = 32'd136314880;
      14244: inst = 32'd268468224;
      14245: inst = 32'd201346505;
      14246: inst = 32'd203470295;
      14247: inst = 32'd136314880;
      14248: inst = 32'd268468224;
      14249: inst = 32'd201346506;
      14250: inst = 32'd203461811;
      14251: inst = 32'd136314880;
      14252: inst = 32'd268468224;
      14253: inst = 32'd201346507;
      14254: inst = 32'd203470263;
      14255: inst = 32'd136314880;
      14256: inst = 32'd268468224;
      14257: inst = 32'd201346508;
      14258: inst = 32'd203470295;
      14259: inst = 32'd136314880;
      14260: inst = 32'd268468224;
      14261: inst = 32'd201346509;
      14262: inst = 32'd203470263;
      14263: inst = 32'd136314880;
      14264: inst = 32'd268468224;
      14265: inst = 32'd201346510;
      14266: inst = 32'd203472343;
      14267: inst = 32'd136314880;
      14268: inst = 32'd268468224;
      14269: inst = 32'd201346511;
      14270: inst = 32'd203472375;
      14271: inst = 32'd136314880;
      14272: inst = 32'd268468224;
      14273: inst = 32'd201346512;
      14274: inst = 32'd203470265;
      14275: inst = 32'd136314880;
      14276: inst = 32'd268468224;
      14277: inst = 32'd201346513;
      14278: inst = 32'd203472377;
      14279: inst = 32'd136314880;
      14280: inst = 32'd268468224;
      14281: inst = 32'd201346514;
      14282: inst = 32'd203472408;
      14283: inst = 32'd136314880;
      14284: inst = 32'd268468224;
      14285: inst = 32'd201346515;
      14286: inst = 32'd203470263;
      14287: inst = 32'd136314880;
      14288: inst = 32'd268468224;
      14289: inst = 32'd201346516;
      14290: inst = 32'd203459666;
      14291: inst = 32'd136314880;
      14292: inst = 32'd268468224;
      14293: inst = 32'd201346517;
      14294: inst = 32'd203451213;
      14295: inst = 32'd136314880;
      14296: inst = 32'd268468224;
      14297: inst = 32'd201346518;
      14298: inst = 32'd203451147;
      14299: inst = 32'd136314880;
      14300: inst = 32'd268468224;
      14301: inst = 32'd201346519;
      14302: inst = 32'd203484952;
      14303: inst = 32'd136314880;
      14304: inst = 32'd268468224;
      14305: inst = 32'd201346520;
      14306: inst = 32'd203484886;
      14307: inst = 32'd136314880;
      14308: inst = 32'd268468224;
      14309: inst = 32'd201346521;
      14310: inst = 32'd203486935;
      14311: inst = 32'd136314880;
      14312: inst = 32'd268468224;
      14313: inst = 32'd201346522;
      14314: inst = 32'd203486903;
      14315: inst = 32'd136314880;
      14316: inst = 32'd268468224;
      14317: inst = 32'd201346523;
      14318: inst = 32'd203486902;
      14319: inst = 32'd136314880;
      14320: inst = 32'd268468224;
      14321: inst = 32'd201346524;
      14322: inst = 32'd203484820;
      14323: inst = 32'd136314880;
      14324: inst = 32'd268468224;
      14325: inst = 32'd201346525;
      14326: inst = 32'd203484820;
      14327: inst = 32'd136314880;
      14328: inst = 32'd268468224;
      14329: inst = 32'd201346526;
      14330: inst = 32'd203486934;
      14331: inst = 32'd136314880;
      14332: inst = 32'd268468224;
      14333: inst = 32'd201346527;
      14334: inst = 32'd203484822;
      14335: inst = 32'd136314880;
      14336: inst = 32'd268468224;
      14337: inst = 32'd201346528;
      14338: inst = 32'd203484886;
      14339: inst = 32'd136314880;
      14340: inst = 32'd268468224;
      14341: inst = 32'd201346529;
      14342: inst = 32'd203484854;
      14343: inst = 32'd136314880;
      14344: inst = 32'd268468224;
      14345: inst = 32'd201346530;
      14346: inst = 32'd203484854;
      14347: inst = 32'd136314880;
      14348: inst = 32'd268468224;
      14349: inst = 32'd201346531;
      14350: inst = 32'd203482806;
      14351: inst = 32'd136314880;
      14352: inst = 32'd268468224;
      14353: inst = 32'd201346532;
      14354: inst = 32'd203482806;
      14355: inst = 32'd136314880;
      14356: inst = 32'd268468224;
      14357: inst = 32'd201346533;
      14358: inst = 32'd203482806;
      14359: inst = 32'd136314880;
      14360: inst = 32'd268468224;
      14361: inst = 32'd201346534;
      14362: inst = 32'd203484854;
      14363: inst = 32'd136314880;
      14364: inst = 32'd268468224;
      14365: inst = 32'd201346535;
      14366: inst = 32'd203484854;
      14367: inst = 32'd136314880;
      14368: inst = 32'd268468224;
      14369: inst = 32'd201346536;
      14370: inst = 32'd203486902;
      14371: inst = 32'd136314880;
      14372: inst = 32'd268468224;
      14373: inst = 32'd201346537;
      14374: inst = 32'd203486902;
      14375: inst = 32'd136314880;
      14376: inst = 32'd268468224;
      14377: inst = 32'd201346538;
      14378: inst = 32'd203486902;
      14379: inst = 32'd136314880;
      14380: inst = 32'd268468224;
      14381: inst = 32'd201346539;
      14382: inst = 32'd203486902;
      14383: inst = 32'd136314880;
      14384: inst = 32'd268468224;
      14385: inst = 32'd201346540;
      14386: inst = 32'd203486902;
      14387: inst = 32'd136314880;
      14388: inst = 32'd268468224;
      14389: inst = 32'd201346541;
      14390: inst = 32'd203486902;
      14391: inst = 32'd136314880;
      14392: inst = 32'd268468224;
      14393: inst = 32'd201346542;
      14394: inst = 32'd203486902;
      14395: inst = 32'd136314880;
      14396: inst = 32'd268468224;
      14397: inst = 32'd201346543;
      14398: inst = 32'd203486902;
      14399: inst = 32'd136314880;
      14400: inst = 32'd268468224;
      14401: inst = 32'd201346544;
      14402: inst = 32'd203486902;
      14403: inst = 32'd136314880;
      14404: inst = 32'd268468224;
      14405: inst = 32'd201346545;
      14406: inst = 32'd203486902;
      14407: inst = 32'd136314880;
      14408: inst = 32'd268468224;
      14409: inst = 32'd201346546;
      14410: inst = 32'd203486902;
      14411: inst = 32'd136314880;
      14412: inst = 32'd268468224;
      14413: inst = 32'd201346547;
      14414: inst = 32'd203486902;
      14415: inst = 32'd136314880;
      14416: inst = 32'd268468224;
      14417: inst = 32'd201346548;
      14418: inst = 32'd203486902;
      14419: inst = 32'd136314880;
      14420: inst = 32'd268468224;
      14421: inst = 32'd201346549;
      14422: inst = 32'd203486902;
      14423: inst = 32'd136314880;
      14424: inst = 32'd268468224;
      14425: inst = 32'd201346550;
      14426: inst = 32'd203486902;
      14427: inst = 32'd136314880;
      14428: inst = 32'd268468224;
      14429: inst = 32'd201346551;
      14430: inst = 32'd203486902;
      14431: inst = 32'd136314880;
      14432: inst = 32'd268468224;
      14433: inst = 32'd201346552;
      14434: inst = 32'd203484854;
      14435: inst = 32'd136314880;
      14436: inst = 32'd268468224;
      14437: inst = 32'd201346553;
      14438: inst = 32'd203484854;
      14439: inst = 32'd136314880;
      14440: inst = 32'd268468224;
      14441: inst = 32'd201346554;
      14442: inst = 32'd203482806;
      14443: inst = 32'd136314880;
      14444: inst = 32'd268468224;
      14445: inst = 32'd201346555;
      14446: inst = 32'd203482806;
      14447: inst = 32'd136314880;
      14448: inst = 32'd268468224;
      14449: inst = 32'd201346556;
      14450: inst = 32'd203482806;
      14451: inst = 32'd136314880;
      14452: inst = 32'd268468224;
      14453: inst = 32'd201346557;
      14454: inst = 32'd203484854;
      14455: inst = 32'd136314880;
      14456: inst = 32'd268468224;
      14457: inst = 32'd201346558;
      14458: inst = 32'd203484854;
      14459: inst = 32'd136314880;
      14460: inst = 32'd268468224;
      14461: inst = 32'd201346559;
      14462: inst = 32'd203484886;
      14463: inst = 32'd136314880;
      14464: inst = 32'd268468224;
      14465: inst = 32'd201346560;
      14466: inst = 32'd203482807;
      14467: inst = 32'd136314880;
      14468: inst = 32'd268468224;
      14469: inst = 32'd201346561;
      14470: inst = 32'd203484887;
      14471: inst = 32'd136314880;
      14472: inst = 32'd268468224;
      14473: inst = 32'd201346562;
      14474: inst = 32'd203484822;
      14475: inst = 32'd136314880;
      14476: inst = 32'd268468224;
      14477: inst = 32'd201346563;
      14478: inst = 32'd203484823;
      14479: inst = 32'd136314880;
      14480: inst = 32'd268468224;
      14481: inst = 32'd201346564;
      14482: inst = 32'd203484887;
      14483: inst = 32'd136314880;
      14484: inst = 32'd268468224;
      14485: inst = 32'd201346565;
      14486: inst = 32'd203486902;
      14487: inst = 32'd136314880;
      14488: inst = 32'd268468224;
      14489: inst = 32'd201346566;
      14490: inst = 32'd203486902;
      14491: inst = 32'd136314880;
      14492: inst = 32'd268468224;
      14493: inst = 32'd201346567;
      14494: inst = 32'd203486934;
      14495: inst = 32'd136314880;
      14496: inst = 32'd268468224;
      14497: inst = 32'd201346568;
      14498: inst = 32'd203484887;
      14499: inst = 32'd136314880;
      14500: inst = 32'd268468224;
      14501: inst = 32'd201346569;
      14502: inst = 32'd203484854;
      14503: inst = 32'd136314880;
      14504: inst = 32'd268468224;
      14505: inst = 32'd201346570;
      14506: inst = 32'd203486901;
      14507: inst = 32'd136314880;
      14508: inst = 32'd268468224;
      14509: inst = 32'd201346571;
      14510: inst = 32'd203484854;
      14511: inst = 32'd136314880;
      14512: inst = 32'd268468224;
      14513: inst = 32'd201346572;
      14514: inst = 32'd203482840;
      14515: inst = 32'd136314880;
      14516: inst = 32'd268468224;
      14517: inst = 32'd201346573;
      14518: inst = 32'd203484856;
      14519: inst = 32'd136314880;
      14520: inst = 32'd268468224;
      14521: inst = 32'd201346574;
      14522: inst = 32'd203488884;
      14523: inst = 32'd136314880;
      14524: inst = 32'd268468224;
      14525: inst = 32'd201346575;
      14526: inst = 32'd203471619;
      14527: inst = 32'd136314880;
      14528: inst = 32'd268468224;
      14529: inst = 32'd201346576;
      14530: inst = 32'd203480005;
      14531: inst = 32'd136314880;
      14532: inst = 32'd268468224;
      14533: inst = 32'd201346577;
      14534: inst = 32'd203480005;
      14535: inst = 32'd136314880;
      14536: inst = 32'd268468224;
      14537: inst = 32'd201346578;
      14538: inst = 32'd203480005;
      14539: inst = 32'd136314880;
      14540: inst = 32'd268468224;
      14541: inst = 32'd201346579;
      14542: inst = 32'd203480005;
      14543: inst = 32'd136314880;
      14544: inst = 32'd268468224;
      14545: inst = 32'd201346580;
      14546: inst = 32'd203480006;
      14547: inst = 32'd136314880;
      14548: inst = 32'd268468224;
      14549: inst = 32'd201346581;
      14550: inst = 32'd203480006;
      14551: inst = 32'd136314880;
      14552: inst = 32'd268468224;
      14553: inst = 32'd201346582;
      14554: inst = 32'd203480006;
      14555: inst = 32'd136314880;
      14556: inst = 32'd268468224;
      14557: inst = 32'd201346583;
      14558: inst = 32'd203480006;
      14559: inst = 32'd136314880;
      14560: inst = 32'd268468224;
      14561: inst = 32'd201346584;
      14562: inst = 32'd203479973;
      14563: inst = 32'd136314880;
      14564: inst = 32'd268468224;
      14565: inst = 32'd201346585;
      14566: inst = 32'd203480038;
      14567: inst = 32'd136314880;
      14568: inst = 32'd268468224;
      14569: inst = 32'd201346586;
      14570: inst = 32'd203479974;
      14571: inst = 32'd136314880;
      14572: inst = 32'd268468224;
      14573: inst = 32'd201346587;
      14574: inst = 32'd203477893;
      14575: inst = 32'd136314880;
      14576: inst = 32'd268468224;
      14577: inst = 32'd201346588;
      14578: inst = 32'd203480006;
      14579: inst = 32'd136314880;
      14580: inst = 32'd268468224;
      14581: inst = 32'd201346589;
      14582: inst = 32'd203479973;
      14583: inst = 32'd136314880;
      14584: inst = 32'd268468224;
      14585: inst = 32'd201346590;
      14586: inst = 32'd203480038;
      14587: inst = 32'd136314880;
      14588: inst = 32'd268468224;
      14589: inst = 32'd201346591;
      14590: inst = 32'd203473667;
      14591: inst = 32'd136314880;
      14592: inst = 32'd268468224;
      14593: inst = 32'd201346592;
      14594: inst = 32'd203461778;
      14595: inst = 32'd136314880;
      14596: inst = 32'd268468224;
      14597: inst = 32'd201346593;
      14598: inst = 32'd203472343;
      14599: inst = 32'd136314880;
      14600: inst = 32'd268468224;
      14601: inst = 32'd201346594;
      14602: inst = 32'd203472343;
      14603: inst = 32'd136314880;
      14604: inst = 32'd268468224;
      14605: inst = 32'd201346595;
      14606: inst = 32'd203472376;
      14607: inst = 32'd136314880;
      14608: inst = 32'd268468224;
      14609: inst = 32'd201346596;
      14610: inst = 32'd203472408;
      14611: inst = 32'd136314880;
      14612: inst = 32'd268468224;
      14613: inst = 32'd201346597;
      14614: inst = 32'd203470263;
      14615: inst = 32'd136314880;
      14616: inst = 32'd268468224;
      14617: inst = 32'd201346598;
      14618: inst = 32'd203470328;
      14619: inst = 32'd136314880;
      14620: inst = 32'd268468224;
      14621: inst = 32'd201346599;
      14622: inst = 32'd203472376;
      14623: inst = 32'd136314880;
      14624: inst = 32'd268468224;
      14625: inst = 32'd201346600;
      14626: inst = 32'd203472376;
      14627: inst = 32'd136314880;
      14628: inst = 32'd268468224;
      14629: inst = 32'd201346601;
      14630: inst = 32'd203470295;
      14631: inst = 32'd136314880;
      14632: inst = 32'd268468224;
      14633: inst = 32'd201346602;
      14634: inst = 32'd203457585;
      14635: inst = 32'd136314880;
      14636: inst = 32'd268468224;
      14637: inst = 32'd201346603;
      14638: inst = 32'd203474488;
      14639: inst = 32'd136314880;
      14640: inst = 32'd268468224;
      14641: inst = 32'd201346604;
      14642: inst = 32'd203472343;
      14643: inst = 32'd136314880;
      14644: inst = 32'd268468224;
      14645: inst = 32'd201346605;
      14646: inst = 32'd203472408;
      14647: inst = 32'd136314880;
      14648: inst = 32'd268468224;
      14649: inst = 32'd201346606;
      14650: inst = 32'd203470262;
      14651: inst = 32'd136314880;
      14652: inst = 32'd268468224;
      14653: inst = 32'd201346607;
      14654: inst = 32'd203472343;
      14655: inst = 32'd136314880;
      14656: inst = 32'd268468224;
      14657: inst = 32'd201346608;
      14658: inst = 32'd203470296;
      14659: inst = 32'd136314880;
      14660: inst = 32'd268468224;
      14661: inst = 32'd201346609;
      14662: inst = 32'd203470295;
      14663: inst = 32'd136314880;
      14664: inst = 32'd268468224;
      14665: inst = 32'd201346610;
      14666: inst = 32'd203470326;
      14667: inst = 32'd136314880;
      14668: inst = 32'd268468224;
      14669: inst = 32'd201346611;
      14670: inst = 32'd203472375;
      14671: inst = 32'd136314880;
      14672: inst = 32'd268468224;
      14673: inst = 32'd201346612;
      14674: inst = 32'd203459730;
      14675: inst = 32'd136314880;
      14676: inst = 32'd268468224;
      14677: inst = 32'd201346613;
      14678: inst = 32'd203453359;
      14679: inst = 32'd136314880;
      14680: inst = 32'd268468224;
      14681: inst = 32'd201346614;
      14682: inst = 32'd203453292;
      14683: inst = 32'd136314880;
      14684: inst = 32'd268468224;
      14685: inst = 32'd201346615;
      14686: inst = 32'd203482839;
      14687: inst = 32'd136314880;
      14688: inst = 32'd268468224;
      14689: inst = 32'd201346616;
      14690: inst = 32'd203482806;
      14691: inst = 32'd136314880;
      14692: inst = 32'd268468224;
      14693: inst = 32'd201346617;
      14694: inst = 32'd203484854;
      14695: inst = 32'd136314880;
      14696: inst = 32'd268468224;
      14697: inst = 32'd201346618;
      14698: inst = 32'd203484823;
      14699: inst = 32'd136314880;
      14700: inst = 32'd268468224;
      14701: inst = 32'd201346619;
      14702: inst = 32'd203486870;
      14703: inst = 32'd136314880;
      14704: inst = 32'd268468224;
      14705: inst = 32'd201346620;
      14706: inst = 32'd203484821;
      14707: inst = 32'd136314880;
      14708: inst = 32'd268468224;
      14709: inst = 32'd201346621;
      14710: inst = 32'd203486902;
      14711: inst = 32'd136314880;
      14712: inst = 32'd268468224;
      14713: inst = 32'd201346622;
      14714: inst = 32'd203489016;
      14715: inst = 32'd136314880;
      14716: inst = 32'd268468224;
      14717: inst = 32'd201346623;
      14718: inst = 32'd203484791;
      14719: inst = 32'd136314880;
      14720: inst = 32'd268468224;
      14721: inst = 32'd201346624;
      14722: inst = 32'd203482807;
      14723: inst = 32'd136314880;
      14724: inst = 32'd268468224;
      14725: inst = 32'd201346625;
      14726: inst = 32'd203482840;
      14727: inst = 32'd136314880;
      14728: inst = 32'd268468224;
      14729: inst = 32'd201346626;
      14730: inst = 32'd203482872;
      14731: inst = 32'd136314880;
      14732: inst = 32'd268468224;
      14733: inst = 32'd201346627;
      14734: inst = 32'd203482872;
      14735: inst = 32'd136314880;
      14736: inst = 32'd268468224;
      14737: inst = 32'd201346628;
      14738: inst = 32'd203482840;
      14739: inst = 32'd136314880;
      14740: inst = 32'd268468224;
      14741: inst = 32'd201346629;
      14742: inst = 32'd203480791;
      14743: inst = 32'd136314880;
      14744: inst = 32'd268468224;
      14745: inst = 32'd201346630;
      14746: inst = 32'd203482840;
      14747: inst = 32'd136314880;
      14748: inst = 32'd268468224;
      14749: inst = 32'd201346631;
      14750: inst = 32'd203484920;
      14751: inst = 32'd136314880;
      14752: inst = 32'd268468224;
      14753: inst = 32'd201346632;
      14754: inst = 32'd203484855;
      14755: inst = 32'd136314880;
      14756: inst = 32'd268468224;
      14757: inst = 32'd201346633;
      14758: inst = 32'd203484855;
      14759: inst = 32'd136314880;
      14760: inst = 32'd268468224;
      14761: inst = 32'd201346634;
      14762: inst = 32'd203484855;
      14763: inst = 32'd136314880;
      14764: inst = 32'd268468224;
      14765: inst = 32'd201346635;
      14766: inst = 32'd203486903;
      14767: inst = 32'd136314880;
      14768: inst = 32'd268468224;
      14769: inst = 32'd201346636;
      14770: inst = 32'd203484854;
      14771: inst = 32'd136314880;
      14772: inst = 32'd268468224;
      14773: inst = 32'd201346637;
      14774: inst = 32'd203484854;
      14775: inst = 32'd136314880;
      14776: inst = 32'd268468224;
      14777: inst = 32'd201346638;
      14778: inst = 32'd203484855;
      14779: inst = 32'd136314880;
      14780: inst = 32'd268468224;
      14781: inst = 32'd201346639;
      14782: inst = 32'd203484855;
      14783: inst = 32'd136314880;
      14784: inst = 32'd268468224;
      14785: inst = 32'd201346640;
      14786: inst = 32'd203484855;
      14787: inst = 32'd136314880;
      14788: inst = 32'd268468224;
      14789: inst = 32'd201346641;
      14790: inst = 32'd203484855;
      14791: inst = 32'd136314880;
      14792: inst = 32'd268468224;
      14793: inst = 32'd201346642;
      14794: inst = 32'd203484854;
      14795: inst = 32'd136314880;
      14796: inst = 32'd268468224;
      14797: inst = 32'd201346643;
      14798: inst = 32'd203484854;
      14799: inst = 32'd136314880;
      14800: inst = 32'd268468224;
      14801: inst = 32'd201346644;
      14802: inst = 32'd203486903;
      14803: inst = 32'd136314880;
      14804: inst = 32'd268468224;
      14805: inst = 32'd201346645;
      14806: inst = 32'd203484855;
      14807: inst = 32'd136314880;
      14808: inst = 32'd268468224;
      14809: inst = 32'd201346646;
      14810: inst = 32'd203484855;
      14811: inst = 32'd136314880;
      14812: inst = 32'd268468224;
      14813: inst = 32'd201346647;
      14814: inst = 32'd203484855;
      14815: inst = 32'd136314880;
      14816: inst = 32'd268468224;
      14817: inst = 32'd201346648;
      14818: inst = 32'd203484920;
      14819: inst = 32'd136314880;
      14820: inst = 32'd268468224;
      14821: inst = 32'd201346649;
      14822: inst = 32'd203482840;
      14823: inst = 32'd136314880;
      14824: inst = 32'd268468224;
      14825: inst = 32'd201346650;
      14826: inst = 32'd203480791;
      14827: inst = 32'd136314880;
      14828: inst = 32'd268468224;
      14829: inst = 32'd201346651;
      14830: inst = 32'd203482840;
      14831: inst = 32'd136314880;
      14832: inst = 32'd268468224;
      14833: inst = 32'd201346652;
      14834: inst = 32'd203482872;
      14835: inst = 32'd136314880;
      14836: inst = 32'd268468224;
      14837: inst = 32'd201346653;
      14838: inst = 32'd203482872;
      14839: inst = 32'd136314880;
      14840: inst = 32'd268468224;
      14841: inst = 32'd201346654;
      14842: inst = 32'd203482840;
      14843: inst = 32'd136314880;
      14844: inst = 32'd268468224;
      14845: inst = 32'd201346655;
      14846: inst = 32'd203482807;
      14847: inst = 32'd136314880;
      14848: inst = 32'd268468224;
      14849: inst = 32'd201346656;
      14850: inst = 32'd203482807;
      14851: inst = 32'd136314880;
      14852: inst = 32'd268468224;
      14853: inst = 32'd201346657;
      14854: inst = 32'd203487000;
      14855: inst = 32'd136314880;
      14856: inst = 32'd268468224;
      14857: inst = 32'd201346658;
      14858: inst = 32'd203486903;
      14859: inst = 32'd136314880;
      14860: inst = 32'd268468224;
      14861: inst = 32'd201346659;
      14862: inst = 32'd203484822;
      14863: inst = 32'd136314880;
      14864: inst = 32'd268468224;
      14865: inst = 32'd201346660;
      14866: inst = 32'd203484855;
      14867: inst = 32'd136314880;
      14868: inst = 32'd268468224;
      14869: inst = 32'd201346661;
      14870: inst = 32'd203484822;
      14871: inst = 32'd136314880;
      14872: inst = 32'd268468224;
      14873: inst = 32'd201346662;
      14874: inst = 32'd203486901;
      14875: inst = 32'd136314880;
      14876: inst = 32'd268468224;
      14877: inst = 32'd201346663;
      14878: inst = 32'd203484854;
      14879: inst = 32'd136314880;
      14880: inst = 32'd268468224;
      14881: inst = 32'd201346664;
      14882: inst = 32'd203484887;
      14883: inst = 32'd136314880;
      14884: inst = 32'd268468224;
      14885: inst = 32'd201346665;
      14886: inst = 32'd203484854;
      14887: inst = 32'd136314880;
      14888: inst = 32'd268468224;
      14889: inst = 32'd201346666;
      14890: inst = 32'd203486901;
      14891: inst = 32'd136314880;
      14892: inst = 32'd268468224;
      14893: inst = 32'd201346667;
      14894: inst = 32'd203484854;
      14895: inst = 32'd136314880;
      14896: inst = 32'd268468224;
      14897: inst = 32'd201346668;
      14898: inst = 32'd203482840;
      14899: inst = 32'd136314880;
      14900: inst = 32'd268468224;
      14901: inst = 32'd201346669;
      14902: inst = 32'd203484856;
      14903: inst = 32'd136314880;
      14904: inst = 32'd268468224;
      14905: inst = 32'd201346670;
      14906: inst = 32'd203488884;
      14907: inst = 32'd136314880;
      14908: inst = 32'd268468224;
      14909: inst = 32'd201346671;
      14910: inst = 32'd203469571;
      14911: inst = 32'd136314880;
      14912: inst = 32'd268468224;
      14913: inst = 32'd201346672;
      14914: inst = 32'd203480005;
      14915: inst = 32'd136314880;
      14916: inst = 32'd268468224;
      14917: inst = 32'd201346673;
      14918: inst = 32'd203480005;
      14919: inst = 32'd136314880;
      14920: inst = 32'd268468224;
      14921: inst = 32'd201346674;
      14922: inst = 32'd203480006;
      14923: inst = 32'd136314880;
      14924: inst = 32'd268468224;
      14925: inst = 32'd201346675;
      14926: inst = 32'd203480006;
      14927: inst = 32'd136314880;
      14928: inst = 32'd268468224;
      14929: inst = 32'd201346676;
      14930: inst = 32'd203480006;
      14931: inst = 32'd136314880;
      14932: inst = 32'd268468224;
      14933: inst = 32'd201346677;
      14934: inst = 32'd203480006;
      14935: inst = 32'd136314880;
      14936: inst = 32'd268468224;
      14937: inst = 32'd201346678;
      14938: inst = 32'd203480006;
      14939: inst = 32'd136314880;
      14940: inst = 32'd268468224;
      14941: inst = 32'd201346679;
      14942: inst = 32'd203480006;
      14943: inst = 32'd136314880;
      14944: inst = 32'd268468224;
      14945: inst = 32'd201346680;
      14946: inst = 32'd203479973;
      14947: inst = 32'd136314880;
      14948: inst = 32'd268468224;
      14949: inst = 32'd201346681;
      14950: inst = 32'd203482086;
      14951: inst = 32'd136314880;
      14952: inst = 32'd268468224;
      14953: inst = 32'd201346682;
      14954: inst = 32'd203479941;
      14955: inst = 32'd136314880;
      14956: inst = 32'd268468224;
      14957: inst = 32'd201346683;
      14958: inst = 32'd203482086;
      14959: inst = 32'd136314880;
      14960: inst = 32'd268468224;
      14961: inst = 32'd201346684;
      14962: inst = 32'd203479973;
      14963: inst = 32'd136314880;
      14964: inst = 32'd268468224;
      14965: inst = 32'd201346685;
      14966: inst = 32'd203482086;
      14967: inst = 32'd136314880;
      14968: inst = 32'd268468224;
      14969: inst = 32'd201346686;
      14970: inst = 32'd203480006;
      14971: inst = 32'd136314880;
      14972: inst = 32'd268468224;
      14973: inst = 32'd201346687;
      14974: inst = 32'd203473634;
      14975: inst = 32'd136314880;
      14976: inst = 32'd268468224;
      14977: inst = 32'd201346688;
      14978: inst = 32'd203459698;
      14979: inst = 32'd136314880;
      14980: inst = 32'd268468224;
      14981: inst = 32'd201346689;
      14982: inst = 32'd203472376;
      14983: inst = 32'd136314880;
      14984: inst = 32'd268468224;
      14985: inst = 32'd201346690;
      14986: inst = 32'd203472343;
      14987: inst = 32'd136314880;
      14988: inst = 32'd268468224;
      14989: inst = 32'd201346691;
      14990: inst = 32'd203470263;
      14991: inst = 32'd136314880;
      14992: inst = 32'd268468224;
      14993: inst = 32'd201346692;
      14994: inst = 32'd203472408;
      14995: inst = 32'd136314880;
      14996: inst = 32'd268468224;
      14997: inst = 32'd201346693;
      14998: inst = 32'd203470295;
      14999: inst = 32'd136314880;
      15000: inst = 32'd268468224;
      15001: inst = 32'd201346694;
      15002: inst = 32'd203470328;
      15003: inst = 32'd136314880;
      15004: inst = 32'd268468224;
      15005: inst = 32'd201346695;
      15006: inst = 32'd203470295;
      15007: inst = 32'd136314880;
      15008: inst = 32'd268468224;
      15009: inst = 32'd201346696;
      15010: inst = 32'd203470263;
      15011: inst = 32'd136314880;
      15012: inst = 32'd268468224;
      15013: inst = 32'd201346697;
      15014: inst = 32'd203472408;
      15015: inst = 32'd136314880;
      15016: inst = 32'd268468224;
      15017: inst = 32'd201346698;
      15018: inst = 32'd203457617;
      15019: inst = 32'd136314880;
      15020: inst = 32'd268468224;
      15021: inst = 32'd201346699;
      15022: inst = 32'd203472376;
      15023: inst = 32'd136314880;
      15024: inst = 32'd268468224;
      15025: inst = 32'd201346700;
      15026: inst = 32'd203470262;
      15027: inst = 32'd136314880;
      15028: inst = 32'd268468224;
      15029: inst = 32'd201346701;
      15030: inst = 32'd203472343;
      15031: inst = 32'd136314880;
      15032: inst = 32'd268468224;
      15033: inst = 32'd201346702;
      15034: inst = 32'd203474456;
      15035: inst = 32'd136314880;
      15036: inst = 32'd268468224;
      15037: inst = 32'd201346703;
      15038: inst = 32'd203472343;
      15039: inst = 32'd136314880;
      15040: inst = 32'd268468224;
      15041: inst = 32'd201346704;
      15042: inst = 32'd203472376;
      15043: inst = 32'd136314880;
      15044: inst = 32'd268468224;
      15045: inst = 32'd201346705;
      15046: inst = 32'd203470327;
      15047: inst = 32'd136314880;
      15048: inst = 32'd268468224;
      15049: inst = 32'd201346706;
      15050: inst = 32'd203470326;
      15051: inst = 32'd136314880;
      15052: inst = 32'd268468224;
      15053: inst = 32'd201346707;
      15054: inst = 32'd203472407;
      15055: inst = 32'd136314880;
      15056: inst = 32'd268468224;
      15057: inst = 32'd201346708;
      15058: inst = 32'd203457585;
      15059: inst = 32'd136314880;
      15060: inst = 32'd268468224;
      15061: inst = 32'd201346709;
      15062: inst = 32'd203451245;
      15063: inst = 32'd136314880;
      15064: inst = 32'd268468224;
      15065: inst = 32'd201346710;
      15066: inst = 32'd203455372;
      15067: inst = 32'd136314880;
      15068: inst = 32'd268468224;
      15069: inst = 32'd201346711;
      15070: inst = 32'd203482839;
      15071: inst = 32'd136314880;
      15072: inst = 32'd268468224;
      15073: inst = 32'd201346712;
      15074: inst = 32'd203484919;
      15075: inst = 32'd136314880;
      15076: inst = 32'd268468224;
      15077: inst = 32'd201346713;
      15078: inst = 32'd203484887;
      15079: inst = 32'd136314880;
      15080: inst = 32'd268468224;
      15081: inst = 32'd201346714;
      15082: inst = 32'd203484823;
      15083: inst = 32'd136314880;
      15084: inst = 32'd268468224;
      15085: inst = 32'd201346715;
      15086: inst = 32'd203486903;
      15087: inst = 32'd136314880;
      15088: inst = 32'd268468224;
      15089: inst = 32'd201346716;
      15090: inst = 32'd203484854;
      15091: inst = 32'd136314880;
      15092: inst = 32'd268468224;
      15093: inst = 32'd201346717;
      15094: inst = 32'd203484854;
      15095: inst = 32'd136314880;
      15096: inst = 32'd268468224;
      15097: inst = 32'd201346718;
      15098: inst = 32'd203482743;
      15099: inst = 32'd136314880;
      15100: inst = 32'd268468224;
      15101: inst = 32'd201346719;
      15102: inst = 32'd203474260;
      15103: inst = 32'd136314880;
      15104: inst = 32'd268468224;
      15105: inst = 32'd201346720;
      15106: inst = 32'd203449099;
      15107: inst = 32'd136314880;
      15108: inst = 32'd268468224;
      15109: inst = 32'd201346721;
      15110: inst = 32'd203449099;
      15111: inst = 32'd136314880;
      15112: inst = 32'd268468224;
      15113: inst = 32'd201346722;
      15114: inst = 32'd203447018;
      15115: inst = 32'd136314880;
      15116: inst = 32'd268468224;
      15117: inst = 32'd201346723;
      15118: inst = 32'd203447018;
      15119: inst = 32'd136314880;
      15120: inst = 32'd268468224;
      15121: inst = 32'd201346724;
      15122: inst = 32'd203449131;
      15123: inst = 32'd136314880;
      15124: inst = 32'd268468224;
      15125: inst = 32'd201346725;
      15126: inst = 32'd203457550;
      15127: inst = 32'd136314880;
      15128: inst = 32'd268468224;
      15129: inst = 32'd201346726;
      15130: inst = 32'd203468115;
      15131: inst = 32'd136314880;
      15132: inst = 32'd268468224;
      15133: inst = 32'd201346727;
      15134: inst = 32'd203476566;
      15135: inst = 32'd136314880;
      15136: inst = 32'd268468224;
      15137: inst = 32'd201346728;
      15138: inst = 32'd203482808;
      15139: inst = 32'd136314880;
      15140: inst = 32'd268468224;
      15141: inst = 32'd201346729;
      15142: inst = 32'd203482807;
      15143: inst = 32'd136314880;
      15144: inst = 32'd268468224;
      15145: inst = 32'd201346730;
      15146: inst = 32'd203484855;
      15147: inst = 32'd136314880;
      15148: inst = 32'd268468224;
      15149: inst = 32'd201346731;
      15150: inst = 32'd203484855;
      15151: inst = 32'd136314880;
      15152: inst = 32'd268468224;
      15153: inst = 32'd201346732;
      15154: inst = 32'd203484855;
      15155: inst = 32'd136314880;
      15156: inst = 32'd268468224;
      15157: inst = 32'd201346733;
      15158: inst = 32'd203484855;
      15159: inst = 32'd136314880;
      15160: inst = 32'd268468224;
      15161: inst = 32'd201346734;
      15162: inst = 32'd203484855;
      15163: inst = 32'd136314880;
      15164: inst = 32'd268468224;
      15165: inst = 32'd201346735;
      15166: inst = 32'd203484855;
      15167: inst = 32'd136314880;
      15168: inst = 32'd268468224;
      15169: inst = 32'd201346736;
      15170: inst = 32'd203484855;
      15171: inst = 32'd136314880;
      15172: inst = 32'd268468224;
      15173: inst = 32'd201346737;
      15174: inst = 32'd203484855;
      15175: inst = 32'd136314880;
      15176: inst = 32'd268468224;
      15177: inst = 32'd201346738;
      15178: inst = 32'd203484855;
      15179: inst = 32'd136314880;
      15180: inst = 32'd268468224;
      15181: inst = 32'd201346739;
      15182: inst = 32'd203484855;
      15183: inst = 32'd136314880;
      15184: inst = 32'd268468224;
      15185: inst = 32'd201346740;
      15186: inst = 32'd203484855;
      15187: inst = 32'd136314880;
      15188: inst = 32'd268468224;
      15189: inst = 32'd201346741;
      15190: inst = 32'd203484855;
      15191: inst = 32'd136314880;
      15192: inst = 32'd268468224;
      15193: inst = 32'd201346742;
      15194: inst = 32'd203482807;
      15195: inst = 32'd136314880;
      15196: inst = 32'd268468224;
      15197: inst = 32'd201346743;
      15198: inst = 32'd203482808;
      15199: inst = 32'd136314880;
      15200: inst = 32'd268468224;
      15201: inst = 32'd201346744;
      15202: inst = 32'd203476566;
      15203: inst = 32'd136314880;
      15204: inst = 32'd268468224;
      15205: inst = 32'd201346745;
      15206: inst = 32'd203468115;
      15207: inst = 32'd136314880;
      15208: inst = 32'd268468224;
      15209: inst = 32'd201346746;
      15210: inst = 32'd203457550;
      15211: inst = 32'd136314880;
      15212: inst = 32'd268468224;
      15213: inst = 32'd201346747;
      15214: inst = 32'd203449131;
      15215: inst = 32'd136314880;
      15216: inst = 32'd268468224;
      15217: inst = 32'd201346748;
      15218: inst = 32'd203447018;
      15219: inst = 32'd136314880;
      15220: inst = 32'd268468224;
      15221: inst = 32'd201346749;
      15222: inst = 32'd203447018;
      15223: inst = 32'd136314880;
      15224: inst = 32'd268468224;
      15225: inst = 32'd201346750;
      15226: inst = 32'd203449099;
      15227: inst = 32'd136314880;
      15228: inst = 32'd268468224;
      15229: inst = 32'd201346751;
      15230: inst = 32'd203449099;
      15231: inst = 32'd136314880;
      15232: inst = 32'd268468224;
      15233: inst = 32'd201346752;
      15234: inst = 32'd203474322;
      15235: inst = 32'd136314880;
      15236: inst = 32'd268468224;
      15237: inst = 32'd201346753;
      15238: inst = 32'd203482741;
      15239: inst = 32'd136314880;
      15240: inst = 32'd268468224;
      15241: inst = 32'd201346754;
      15242: inst = 32'd203486902;
      15243: inst = 32'd136314880;
      15244: inst = 32'd268468224;
      15245: inst = 32'd201346755;
      15246: inst = 32'd203484855;
      15247: inst = 32'd136314880;
      15248: inst = 32'd268468224;
      15249: inst = 32'd201346756;
      15250: inst = 32'd203484887;
      15251: inst = 32'd136314880;
      15252: inst = 32'd268468224;
      15253: inst = 32'd201346757;
      15254: inst = 32'd203486870;
      15255: inst = 32'd136314880;
      15256: inst = 32'd268468224;
      15257: inst = 32'd201346758;
      15258: inst = 32'd203486902;
      15259: inst = 32'd136314880;
      15260: inst = 32'd268468224;
      15261: inst = 32'd201346759;
      15262: inst = 32'd203486934;
      15263: inst = 32'd136314880;
      15264: inst = 32'd268468224;
      15265: inst = 32'd201346760;
      15266: inst = 32'd203484887;
      15267: inst = 32'd136314880;
      15268: inst = 32'd268468224;
      15269: inst = 32'd201346761;
      15270: inst = 32'd203484854;
      15271: inst = 32'd136314880;
      15272: inst = 32'd268468224;
      15273: inst = 32'd201346762;
      15274: inst = 32'd203486901;
      15275: inst = 32'd136314880;
      15276: inst = 32'd268468224;
      15277: inst = 32'd201346763;
      15278: inst = 32'd203484854;
      15279: inst = 32'd136314880;
      15280: inst = 32'd268468224;
      15281: inst = 32'd201346764;
      15282: inst = 32'd203482840;
      15283: inst = 32'd136314880;
      15284: inst = 32'd268468224;
      15285: inst = 32'd201346765;
      15286: inst = 32'd203484856;
      15287: inst = 32'd136314880;
      15288: inst = 32'd268468224;
      15289: inst = 32'd201346766;
      15290: inst = 32'd203488884;
      15291: inst = 32'd136314880;
      15292: inst = 32'd268468224;
      15293: inst = 32'd201346767;
      15294: inst = 32'd203469571;
      15295: inst = 32'd136314880;
      15296: inst = 32'd268468224;
      15297: inst = 32'd201346768;
      15298: inst = 32'd203480006;
      15299: inst = 32'd136314880;
      15300: inst = 32'd268468224;
      15301: inst = 32'd201346769;
      15302: inst = 32'd203480006;
      15303: inst = 32'd136314880;
      15304: inst = 32'd268468224;
      15305: inst = 32'd201346770;
      15306: inst = 32'd203480006;
      15307: inst = 32'd136314880;
      15308: inst = 32'd268468224;
      15309: inst = 32'd201346771;
      15310: inst = 32'd203480006;
      15311: inst = 32'd136314880;
      15312: inst = 32'd268468224;
      15313: inst = 32'd201346772;
      15314: inst = 32'd203480005;
      15315: inst = 32'd136314880;
      15316: inst = 32'd268468224;
      15317: inst = 32'd201346773;
      15318: inst = 32'd203480005;
      15319: inst = 32'd136314880;
      15320: inst = 32'd268468224;
      15321: inst = 32'd201346774;
      15322: inst = 32'd203480005;
      15323: inst = 32'd136314880;
      15324: inst = 32'd268468224;
      15325: inst = 32'd201346775;
      15326: inst = 32'd203480005;
      15327: inst = 32'd136314880;
      15328: inst = 32'd268468224;
      15329: inst = 32'd201346776;
      15330: inst = 32'd203480005;
      15331: inst = 32'd136314880;
      15332: inst = 32'd268468224;
      15333: inst = 32'd201346777;
      15334: inst = 32'd203479973;
      15335: inst = 32'd136314880;
      15336: inst = 32'd268468224;
      15337: inst = 32'd201346778;
      15338: inst = 32'd203482054;
      15339: inst = 32'd136314880;
      15340: inst = 32'd268468224;
      15341: inst = 32'd201346779;
      15342: inst = 32'd203482054;
      15343: inst = 32'd136314880;
      15344: inst = 32'd268468224;
      15345: inst = 32'd201346780;
      15346: inst = 32'd203480005;
      15347: inst = 32'd136314880;
      15348: inst = 32'd268468224;
      15349: inst = 32'd201346781;
      15350: inst = 32'd203479973;
      15351: inst = 32'd136314880;
      15352: inst = 32'd268468224;
      15353: inst = 32'd201346782;
      15354: inst = 32'd203482086;
      15355: inst = 32'd136314880;
      15356: inst = 32'd268468224;
      15357: inst = 32'd201346783;
      15358: inst = 32'd203473634;
      15359: inst = 32'd136314880;
      15360: inst = 32'd268468224;
      15361: inst = 32'd201346784;
      15362: inst = 32'd203459698;
      15363: inst = 32'd136314880;
      15364: inst = 32'd268468224;
      15365: inst = 32'd201346785;
      15366: inst = 32'd203472376;
      15367: inst = 32'd136314880;
      15368: inst = 32'd268468224;
      15369: inst = 32'd201346786;
      15370: inst = 32'd203472344;
      15371: inst = 32'd136314880;
      15372: inst = 32'd268468224;
      15373: inst = 32'd201346787;
      15374: inst = 32'd203472344;
      15375: inst = 32'd136314880;
      15376: inst = 32'd268468224;
      15377: inst = 32'd201346788;
      15378: inst = 32'd203472344;
      15379: inst = 32'd136314880;
      15380: inst = 32'd268468224;
      15381: inst = 32'd201346789;
      15382: inst = 32'd203472376;
      15383: inst = 32'd136314880;
      15384: inst = 32'd268468224;
      15385: inst = 32'd201346790;
      15386: inst = 32'd203472344;
      15387: inst = 32'd136314880;
      15388: inst = 32'd268468224;
      15389: inst = 32'd201346791;
      15390: inst = 32'd203472376;
      15391: inst = 32'd136314880;
      15392: inst = 32'd268468224;
      15393: inst = 32'd201346792;
      15394: inst = 32'd203470263;
      15395: inst = 32'd136314880;
      15396: inst = 32'd268468224;
      15397: inst = 32'd201346793;
      15398: inst = 32'd203472408;
      15399: inst = 32'd136314880;
      15400: inst = 32'd268468224;
      15401: inst = 32'd201346794;
      15402: inst = 32'd203459665;
      15403: inst = 32'd136314880;
      15404: inst = 32'd268468224;
      15405: inst = 32'd201346795;
      15406: inst = 32'd203470262;
      15407: inst = 32'd136314880;
      15408: inst = 32'd268468224;
      15409: inst = 32'd201346796;
      15410: inst = 32'd203474456;
      15411: inst = 32'd136314880;
      15412: inst = 32'd268468224;
      15413: inst = 32'd201346797;
      15414: inst = 32'd203472375;
      15415: inst = 32'd136314880;
      15416: inst = 32'd268468224;
      15417: inst = 32'd201346798;
      15418: inst = 32'd203472310;
      15419: inst = 32'd136314880;
      15420: inst = 32'd268468224;
      15421: inst = 32'd201346799;
      15422: inst = 32'd203472375;
      15423: inst = 32'd136314880;
      15424: inst = 32'd268468224;
      15425: inst = 32'd201346800;
      15426: inst = 32'd203470295;
      15427: inst = 32'd136314880;
      15428: inst = 32'd268468224;
      15429: inst = 32'd201346801;
      15430: inst = 32'd203472375;
      15431: inst = 32'd136314880;
      15432: inst = 32'd268468224;
      15433: inst = 32'd201346802;
      15434: inst = 32'd203470325;
      15435: inst = 32'd136314880;
      15436: inst = 32'd268468224;
      15437: inst = 32'd201346803;
      15438: inst = 32'd203472374;
      15439: inst = 32'd136314880;
      15440: inst = 32'd268468224;
      15441: inst = 32'd201346804;
      15442: inst = 32'd203459697;
      15443: inst = 32'd136314880;
      15444: inst = 32'd268468224;
      15445: inst = 32'd201346805;
      15446: inst = 32'd203453293;
      15447: inst = 32'd136314880;
      15448: inst = 32'd268468224;
      15449: inst = 32'd201346806;
      15450: inst = 32'd203453292;
      15451: inst = 32'd136314880;
      15452: inst = 32'd268468224;
      15453: inst = 32'd201346807;
      15454: inst = 32'd203482839;
      15455: inst = 32'd136314880;
      15456: inst = 32'd268468224;
      15457: inst = 32'd201346808;
      15458: inst = 32'd203482838;
      15459: inst = 32'd136314880;
      15460: inst = 32'd268468224;
      15461: inst = 32'd201346809;
      15462: inst = 32'd203484887;
      15463: inst = 32'd136314880;
      15464: inst = 32'd268468224;
      15465: inst = 32'd201346810;
      15466: inst = 32'd203486936;
      15467: inst = 32'd136314880;
      15468: inst = 32'd268468224;
      15469: inst = 32'd201346811;
      15470: inst = 32'd203482742;
      15471: inst = 32'd136314880;
      15472: inst = 32'd268468224;
      15473: inst = 32'd201346812;
      15474: inst = 32'd203486935;
      15475: inst = 32'd136314880;
      15476: inst = 32'd268468224;
      15477: inst = 32'd201346813;
      15478: inst = 32'd203484855;
      15479: inst = 32'd136314880;
      15480: inst = 32'd268468224;
      15481: inst = 32'd201346814;
      15482: inst = 32'd203482776;
      15483: inst = 32'd136314880;
      15484: inst = 32'd268468224;
      15485: inst = 32'd201346815;
      15486: inst = 32'd203467954;
      15487: inst = 32'd136314880;
      15488: inst = 32'd268468224;
      15489: inst = 32'd201346816;
      15490: inst = 32'd203447020;
      15491: inst = 32'd136314880;
      15492: inst = 32'd268468224;
      15493: inst = 32'd201346817;
      15494: inst = 32'd203449100;
      15495: inst = 32'd136314880;
      15496: inst = 32'd268468224;
      15497: inst = 32'd201346818;
      15498: inst = 32'd203447052;
      15499: inst = 32'd136314880;
      15500: inst = 32'd268468224;
      15501: inst = 32'd201346819;
      15502: inst = 32'd203447020;
      15503: inst = 32'd136314880;
      15504: inst = 32'd268468224;
      15505: inst = 32'd201346820;
      15506: inst = 32'd203449133;
      15507: inst = 32'd136314880;
      15508: inst = 32'd268468224;
      15509: inst = 32'd201346821;
      15510: inst = 32'd203447019;
      15511: inst = 32'd136314880;
      15512: inst = 32'd268468224;
      15513: inst = 32'd201346822;
      15514: inst = 32'd203449099;
      15515: inst = 32'd136314880;
      15516: inst = 32'd268468224;
      15517: inst = 32'd201346823;
      15518: inst = 32'd203461711;
      15519: inst = 32'd136314880;
      15520: inst = 32'd268468224;
      15521: inst = 32'd201346824;
      15522: inst = 32'd203480728;
      15523: inst = 32'd136314880;
      15524: inst = 32'd268468224;
      15525: inst = 32'd201346825;
      15526: inst = 32'd203482808;
      15527: inst = 32'd136314880;
      15528: inst = 32'd268468224;
      15529: inst = 32'd201346826;
      15530: inst = 32'd203484888;
      15531: inst = 32'd136314880;
      15532: inst = 32'd268468224;
      15533: inst = 32'd201346827;
      15534: inst = 32'd203484855;
      15535: inst = 32'd136314880;
      15536: inst = 32'd268468224;
      15537: inst = 32'd201346828;
      15538: inst = 32'd203484855;
      15539: inst = 32'd136314880;
      15540: inst = 32'd268468224;
      15541: inst = 32'd201346829;
      15542: inst = 32'd203484887;
      15543: inst = 32'd136314880;
      15544: inst = 32'd268468224;
      15545: inst = 32'd201346830;
      15546: inst = 32'd203482774;
      15547: inst = 32'd136314880;
      15548: inst = 32'd268468224;
      15549: inst = 32'd201346831;
      15550: inst = 32'd203484920;
      15551: inst = 32'd136314880;
      15552: inst = 32'd268468224;
      15553: inst = 32'd201346832;
      15554: inst = 32'd203484920;
      15555: inst = 32'd136314880;
      15556: inst = 32'd268468224;
      15557: inst = 32'd201346833;
      15558: inst = 32'd203482774;
      15559: inst = 32'd136314880;
      15560: inst = 32'd268468224;
      15561: inst = 32'd201346834;
      15562: inst = 32'd203484887;
      15563: inst = 32'd136314880;
      15564: inst = 32'd268468224;
      15565: inst = 32'd201346835;
      15566: inst = 32'd203484855;
      15567: inst = 32'd136314880;
      15568: inst = 32'd268468224;
      15569: inst = 32'd201346836;
      15570: inst = 32'd203484855;
      15571: inst = 32'd136314880;
      15572: inst = 32'd268468224;
      15573: inst = 32'd201346837;
      15574: inst = 32'd203484888;
      15575: inst = 32'd136314880;
      15576: inst = 32'd268468224;
      15577: inst = 32'd201346838;
      15578: inst = 32'd203482808;
      15579: inst = 32'd136314880;
      15580: inst = 32'd268468224;
      15581: inst = 32'd201346839;
      15582: inst = 32'd203480728;
      15583: inst = 32'd136314880;
      15584: inst = 32'd268468224;
      15585: inst = 32'd201346840;
      15586: inst = 32'd203461712;
      15587: inst = 32'd136314880;
      15588: inst = 32'd268468224;
      15589: inst = 32'd201346841;
      15590: inst = 32'd203449099;
      15591: inst = 32'd136314880;
      15592: inst = 32'd268468224;
      15593: inst = 32'd201346842;
      15594: inst = 32'd203447019;
      15595: inst = 32'd136314880;
      15596: inst = 32'd268468224;
      15597: inst = 32'd201346843;
      15598: inst = 32'd203449133;
      15599: inst = 32'd136314880;
      15600: inst = 32'd268468224;
      15601: inst = 32'd201346844;
      15602: inst = 32'd203447020;
      15603: inst = 32'd136314880;
      15604: inst = 32'd268468224;
      15605: inst = 32'd201346845;
      15606: inst = 32'd203447052;
      15607: inst = 32'd136314880;
      15608: inst = 32'd268468224;
      15609: inst = 32'd201346846;
      15610: inst = 32'd203449100;
      15611: inst = 32'd136314880;
      15612: inst = 32'd268468224;
      15613: inst = 32'd201346847;
      15614: inst = 32'd203447020;
      15615: inst = 32'd136314880;
      15616: inst = 32'd268468224;
      15617: inst = 32'd201346848;
      15618: inst = 32'd203467983;
      15619: inst = 32'd136314880;
      15620: inst = 32'd268468224;
      15621: inst = 32'd201346849;
      15622: inst = 32'd203484822;
      15623: inst = 32'd136314880;
      15624: inst = 32'd268468224;
      15625: inst = 32'd201346850;
      15626: inst = 32'd203484822;
      15627: inst = 32'd136314880;
      15628: inst = 32'd268468224;
      15629: inst = 32'd201346851;
      15630: inst = 32'd203486935;
      15631: inst = 32'd136314880;
      15632: inst = 32'd268468224;
      15633: inst = 32'd201346852;
      15634: inst = 32'd203482742;
      15635: inst = 32'd136314880;
      15636: inst = 32'd268468224;
      15637: inst = 32'd201346853;
      15638: inst = 32'd203486902;
      15639: inst = 32'd136314880;
      15640: inst = 32'd268468224;
      15641: inst = 32'd201346854;
      15642: inst = 32'd203486901;
      15643: inst = 32'd136314880;
      15644: inst = 32'd268468224;
      15645: inst = 32'd201346855;
      15646: inst = 32'd203484854;
      15647: inst = 32'd136314880;
      15648: inst = 32'd268468224;
      15649: inst = 32'd201346856;
      15650: inst = 32'd203484887;
      15651: inst = 32'd136314880;
      15652: inst = 32'd268468224;
      15653: inst = 32'd201346857;
      15654: inst = 32'd203484854;
      15655: inst = 32'd136314880;
      15656: inst = 32'd268468224;
      15657: inst = 32'd201346858;
      15658: inst = 32'd203486901;
      15659: inst = 32'd136314880;
      15660: inst = 32'd268468224;
      15661: inst = 32'd201346859;
      15662: inst = 32'd203484854;
      15663: inst = 32'd136314880;
      15664: inst = 32'd268468224;
      15665: inst = 32'd201346860;
      15666: inst = 32'd203482840;
      15667: inst = 32'd136314880;
      15668: inst = 32'd268468224;
      15669: inst = 32'd201346861;
      15670: inst = 32'd203484856;
      15671: inst = 32'd136314880;
      15672: inst = 32'd268468224;
      15673: inst = 32'd201346862;
      15674: inst = 32'd203488884;
      15675: inst = 32'd136314880;
      15676: inst = 32'd268468224;
      15677: inst = 32'd201346863;
      15678: inst = 32'd203469571;
      15679: inst = 32'd136314880;
      15680: inst = 32'd268468224;
      15681: inst = 32'd201346864;
      15682: inst = 32'd203480006;
      15683: inst = 32'd136314880;
      15684: inst = 32'd268468224;
      15685: inst = 32'd201346865;
      15686: inst = 32'd203480006;
      15687: inst = 32'd136314880;
      15688: inst = 32'd268468224;
      15689: inst = 32'd201346866;
      15690: inst = 32'd203480006;
      15691: inst = 32'd136314880;
      15692: inst = 32'd268468224;
      15693: inst = 32'd201346867;
      15694: inst = 32'd203480006;
      15695: inst = 32'd136314880;
      15696: inst = 32'd268468224;
      15697: inst = 32'd201346868;
      15698: inst = 32'd203480005;
      15699: inst = 32'd136314880;
      15700: inst = 32'd268468224;
      15701: inst = 32'd201346869;
      15702: inst = 32'd203480005;
      15703: inst = 32'd136314880;
      15704: inst = 32'd268468224;
      15705: inst = 32'd201346870;
      15706: inst = 32'd203480005;
      15707: inst = 32'd136314880;
      15708: inst = 32'd268468224;
      15709: inst = 32'd201346871;
      15710: inst = 32'd203480005;
      15711: inst = 32'd136314880;
      15712: inst = 32'd268468224;
      15713: inst = 32'd201346872;
      15714: inst = 32'd203480005;
      15715: inst = 32'd136314880;
      15716: inst = 32'd268468224;
      15717: inst = 32'd201346873;
      15718: inst = 32'd203482053;
      15719: inst = 32'd136314880;
      15720: inst = 32'd268468224;
      15721: inst = 32'd201346874;
      15722: inst = 32'd203479973;
      15723: inst = 32'd136314880;
      15724: inst = 32'd268468224;
      15725: inst = 32'd201346875;
      15726: inst = 32'd203482053;
      15727: inst = 32'd136314880;
      15728: inst = 32'd268468224;
      15729: inst = 32'd201346876;
      15730: inst = 32'd203479973;
      15731: inst = 32'd136314880;
      15732: inst = 32'd268468224;
      15733: inst = 32'd201346877;
      15734: inst = 32'd203482053;
      15735: inst = 32'd136314880;
      15736: inst = 32'd268468224;
      15737: inst = 32'd201346878;
      15738: inst = 32'd203479973;
      15739: inst = 32'd136314880;
      15740: inst = 32'd268468224;
      15741: inst = 32'd201346879;
      15742: inst = 32'd203473634;
      15743: inst = 32'd136314880;
      15744: inst = 32'd268468224;
      15745: inst = 32'd201346880;
      15746: inst = 32'd203459698;
      15747: inst = 32'd136314880;
      15748: inst = 32'd268468224;
      15749: inst = 32'd201346881;
      15750: inst = 32'd203472376;
      15751: inst = 32'd136314880;
      15752: inst = 32'd268468224;
      15753: inst = 32'd201346882;
      15754: inst = 32'd203472343;
      15755: inst = 32'd136314880;
      15756: inst = 32'd268468224;
      15757: inst = 32'd201346883;
      15758: inst = 32'd203472343;
      15759: inst = 32'd136314880;
      15760: inst = 32'd268468224;
      15761: inst = 32'd201346884;
      15762: inst = 32'd203472343;
      15763: inst = 32'd136314880;
      15764: inst = 32'd268468224;
      15765: inst = 32'd201346885;
      15766: inst = 32'd203472376;
      15767: inst = 32'd136314880;
      15768: inst = 32'd268468224;
      15769: inst = 32'd201346886;
      15770: inst = 32'd203472343;
      15771: inst = 32'd136314880;
      15772: inst = 32'd268468224;
      15773: inst = 32'd201346887;
      15774: inst = 32'd203472375;
      15775: inst = 32'd136314880;
      15776: inst = 32'd268468224;
      15777: inst = 32'd201346888;
      15778: inst = 32'd203474456;
      15779: inst = 32'd136314880;
      15780: inst = 32'd268468224;
      15781: inst = 32'd201346889;
      15782: inst = 32'd203472343;
      15783: inst = 32'd136314880;
      15784: inst = 32'd268468224;
      15785: inst = 32'd201346890;
      15786: inst = 32'd203459697;
      15787: inst = 32'd136314880;
      15788: inst = 32'd268468224;
      15789: inst = 32'd201346891;
      15790: inst = 32'd203474455;
      15791: inst = 32'd136314880;
      15792: inst = 32'd268468224;
      15793: inst = 32'd201346892;
      15794: inst = 32'd203472375;
      15795: inst = 32'd136314880;
      15796: inst = 32'd268468224;
      15797: inst = 32'd201346893;
      15798: inst = 32'd203472310;
      15799: inst = 32'd136314880;
      15800: inst = 32'd268468224;
      15801: inst = 32'd201346894;
      15802: inst = 32'd203472343;
      15803: inst = 32'd136314880;
      15804: inst = 32'd268468224;
      15805: inst = 32'd201346895;
      15806: inst = 32'd203472342;
      15807: inst = 32'd136314880;
      15808: inst = 32'd268468224;
      15809: inst = 32'd201346896;
      15810: inst = 32'd203472343;
      15811: inst = 32'd136314880;
      15812: inst = 32'd268468224;
      15813: inst = 32'd201346897;
      15814: inst = 32'd203472375;
      15815: inst = 32'd136314880;
      15816: inst = 32'd268468224;
      15817: inst = 32'd201346898;
      15818: inst = 32'd203472374;
      15819: inst = 32'd136314880;
      15820: inst = 32'd268468224;
      15821: inst = 32'd201346899;
      15822: inst = 32'd203472375;
      15823: inst = 32'd136314880;
      15824: inst = 32'd268468224;
      15825: inst = 32'd201346900;
      15826: inst = 32'd203459698;
      15827: inst = 32'd136314880;
      15828: inst = 32'd268468224;
      15829: inst = 32'd201346901;
      15830: inst = 32'd203453294;
      15831: inst = 32'd136314880;
      15832: inst = 32'd268468224;
      15833: inst = 32'd201346902;
      15834: inst = 32'd203453260;
      15835: inst = 32'd136314880;
      15836: inst = 32'd268468224;
      15837: inst = 32'd201346903;
      15838: inst = 32'd203482839;
      15839: inst = 32'd136314880;
      15840: inst = 32'd268468224;
      15841: inst = 32'd201346904;
      15842: inst = 32'd203484886;
      15843: inst = 32'd136314880;
      15844: inst = 32'd268468224;
      15845: inst = 32'd201346905;
      15846: inst = 32'd203484887;
      15847: inst = 32'd136314880;
      15848: inst = 32'd268468224;
      15849: inst = 32'd201346906;
      15850: inst = 32'd203484855;
      15851: inst = 32'd136314880;
      15852: inst = 32'd268468224;
      15853: inst = 32'd201346907;
      15854: inst = 32'd203482774;
      15855: inst = 32'd136314880;
      15856: inst = 32'd268468224;
      15857: inst = 32'd201346908;
      15858: inst = 32'd203484887;
      15859: inst = 32'd136314880;
      15860: inst = 32'd268468224;
      15861: inst = 32'd201346909;
      15862: inst = 32'd203482806;
      15863: inst = 32'd136314880;
      15864: inst = 32'd268468224;
      15865: inst = 32'd201346910;
      15866: inst = 32'd203484889;
      15867: inst = 32'd136314880;
      15868: inst = 32'd268468224;
      15869: inst = 32'd201346911;
      15870: inst = 32'd203467954;
      15871: inst = 32'd136314880;
      15872: inst = 32'd268468224;
      15873: inst = 32'd201346912;
      15874: inst = 32'd203447021;
      15875: inst = 32'd136314880;
      15876: inst = 32'd268468224;
      15877: inst = 32'd201346913;
      15878: inst = 32'd203449101;
      15879: inst = 32'd136314880;
      15880: inst = 32'd268468224;
      15881: inst = 32'd201346914;
      15882: inst = 32'd203447021;
      15883: inst = 32'd136314880;
      15884: inst = 32'd268468224;
      15885: inst = 32'd201346915;
      15886: inst = 32'd203446988;
      15887: inst = 32'd136314880;
      15888: inst = 32'd268468224;
      15889: inst = 32'd201346916;
      15890: inst = 32'd203447053;
      15891: inst = 32'd136314880;
      15892: inst = 32'd268468224;
      15893: inst = 32'd201346917;
      15894: inst = 32'd203449101;
      15895: inst = 32'd136314880;
      15896: inst = 32'd268468224;
      15897: inst = 32'd201346918;
      15898: inst = 32'd203446987;
      15899: inst = 32'd136314880;
      15900: inst = 32'd268468224;
      15901: inst = 32'd201346919;
      15902: inst = 32'd203451180;
      15903: inst = 32'd136314880;
      15904: inst = 32'd268468224;
      15905: inst = 32'd201346920;
      15906: inst = 32'd203482841;
      15907: inst = 32'd136314880;
      15908: inst = 32'd268468224;
      15909: inst = 32'd201346921;
      15910: inst = 32'd203484888;
      15911: inst = 32'd136314880;
      15912: inst = 32'd268468224;
      15913: inst = 32'd201346922;
      15914: inst = 32'd203484887;
      15915: inst = 32'd136314880;
      15916: inst = 32'd268468224;
      15917: inst = 32'd201346923;
      15918: inst = 32'd203484855;
      15919: inst = 32'd136314880;
      15920: inst = 32'd268468224;
      15921: inst = 32'd201346924;
      15922: inst = 32'd203484887;
      15923: inst = 32'd136314880;
      15924: inst = 32'd268468224;
      15925: inst = 32'd201346925;
      15926: inst = 32'd203484887;
      15927: inst = 32'd136314880;
      15928: inst = 32'd268468224;
      15929: inst = 32'd201346926;
      15930: inst = 32'd203484854;
      15931: inst = 32'd136314880;
      15932: inst = 32'd268468224;
      15933: inst = 32'd201346927;
      15934: inst = 32'd203484854;
      15935: inst = 32'd136314880;
      15936: inst = 32'd268468224;
      15937: inst = 32'd201346928;
      15938: inst = 32'd203484854;
      15939: inst = 32'd136314880;
      15940: inst = 32'd268468224;
      15941: inst = 32'd201346929;
      15942: inst = 32'd203484854;
      15943: inst = 32'd136314880;
      15944: inst = 32'd268468224;
      15945: inst = 32'd201346930;
      15946: inst = 32'd203484887;
      15947: inst = 32'd136314880;
      15948: inst = 32'd268468224;
      15949: inst = 32'd201346931;
      15950: inst = 32'd203484887;
      15951: inst = 32'd136314880;
      15952: inst = 32'd268468224;
      15953: inst = 32'd201346932;
      15954: inst = 32'd203484855;
      15955: inst = 32'd136314880;
      15956: inst = 32'd268468224;
      15957: inst = 32'd201346933;
      15958: inst = 32'd203484887;
      15959: inst = 32'd136314880;
      15960: inst = 32'd268468224;
      15961: inst = 32'd201346934;
      15962: inst = 32'd203484888;
      15963: inst = 32'd136314880;
      15964: inst = 32'd268468224;
      15965: inst = 32'd201346935;
      15966: inst = 32'd203482841;
      15967: inst = 32'd136314880;
      15968: inst = 32'd268468224;
      15969: inst = 32'd201346936;
      15970: inst = 32'd203451179;
      15971: inst = 32'd136314880;
      15972: inst = 32'd268468224;
      15973: inst = 32'd201346937;
      15974: inst = 32'd203446987;
      15975: inst = 32'd136314880;
      15976: inst = 32'd268468224;
      15977: inst = 32'd201346938;
      15978: inst = 32'd203449101;
      15979: inst = 32'd136314880;
      15980: inst = 32'd268468224;
      15981: inst = 32'd201346939;
      15982: inst = 32'd203447053;
      15983: inst = 32'd136314880;
      15984: inst = 32'd268468224;
      15985: inst = 32'd201346940;
      15986: inst = 32'd203446988;
      15987: inst = 32'd136314880;
      15988: inst = 32'd268468224;
      15989: inst = 32'd201346941;
      15990: inst = 32'd203447021;
      15991: inst = 32'd136314880;
      15992: inst = 32'd268468224;
      15993: inst = 32'd201346942;
      15994: inst = 32'd203449101;
      15995: inst = 32'd136314880;
      15996: inst = 32'd268468224;
      15997: inst = 32'd201346943;
      15998: inst = 32'd203447021;
      15999: inst = 32'd136314880;
      16000: inst = 32'd268468224;
      16001: inst = 32'd201346944;
      16002: inst = 32'd203467984;
      16003: inst = 32'd136314880;
      16004: inst = 32'd268468224;
      16005: inst = 32'd201346945;
      16006: inst = 32'd203486935;
      16007: inst = 32'd136314880;
      16008: inst = 32'd268468224;
      16009: inst = 32'd201346946;
      16010: inst = 32'd203484822;
      16011: inst = 32'd136314880;
      16012: inst = 32'd268468224;
      16013: inst = 32'd201346947;
      16014: inst = 32'd203486935;
      16015: inst = 32'd136314880;
      16016: inst = 32'd268468224;
      16017: inst = 32'd201346948;
      16018: inst = 32'd203482774;
      16019: inst = 32'd136314880;
      16020: inst = 32'd268468224;
      16021: inst = 32'd201346949;
      16022: inst = 32'd203486870;
      16023: inst = 32'd136314880;
      16024: inst = 32'd268468224;
      16025: inst = 32'd201346950;
      16026: inst = 32'd203486901;
      16027: inst = 32'd136314880;
      16028: inst = 32'd268468224;
      16029: inst = 32'd201346951;
      16030: inst = 32'd203484854;
      16031: inst = 32'd136314880;
      16032: inst = 32'd268468224;
      16033: inst = 32'd201346952;
      16034: inst = 32'd203484887;
      16035: inst = 32'd136314880;
      16036: inst = 32'd268468224;
      16037: inst = 32'd201346953;
      16038: inst = 32'd203484854;
      16039: inst = 32'd136314880;
      16040: inst = 32'd268468224;
      16041: inst = 32'd201346954;
      16042: inst = 32'd203486901;
      16043: inst = 32'd136314880;
      16044: inst = 32'd268468224;
      16045: inst = 32'd201346955;
      16046: inst = 32'd203484854;
      16047: inst = 32'd136314880;
      16048: inst = 32'd268468224;
      16049: inst = 32'd201346956;
      16050: inst = 32'd203482840;
      16051: inst = 32'd136314880;
      16052: inst = 32'd268468224;
      16053: inst = 32'd201346957;
      16054: inst = 32'd203484856;
      16055: inst = 32'd136314880;
      16056: inst = 32'd268468224;
      16057: inst = 32'd201346958;
      16058: inst = 32'd203488884;
      16059: inst = 32'd136314880;
      16060: inst = 32'd268468224;
      16061: inst = 32'd201346959;
      16062: inst = 32'd203469571;
      16063: inst = 32'd136314880;
      16064: inst = 32'd268468224;
      16065: inst = 32'd201346960;
      16066: inst = 32'd203480006;
      16067: inst = 32'd136314880;
      16068: inst = 32'd268468224;
      16069: inst = 32'd201346961;
      16070: inst = 32'd203480006;
      16071: inst = 32'd136314880;
      16072: inst = 32'd268468224;
      16073: inst = 32'd201346962;
      16074: inst = 32'd203480006;
      16075: inst = 32'd136314880;
      16076: inst = 32'd268468224;
      16077: inst = 32'd201346963;
      16078: inst = 32'd203480006;
      16079: inst = 32'd136314880;
      16080: inst = 32'd268468224;
      16081: inst = 32'd201346964;
      16082: inst = 32'd203480005;
      16083: inst = 32'd136314880;
      16084: inst = 32'd268468224;
      16085: inst = 32'd201346965;
      16086: inst = 32'd203480005;
      16087: inst = 32'd136314880;
      16088: inst = 32'd268468224;
      16089: inst = 32'd201346966;
      16090: inst = 32'd203480005;
      16091: inst = 32'd136314880;
      16092: inst = 32'd268468224;
      16093: inst = 32'd201346967;
      16094: inst = 32'd203480005;
      16095: inst = 32'd136314880;
      16096: inst = 32'd268468224;
      16097: inst = 32'd201346968;
      16098: inst = 32'd203482053;
      16099: inst = 32'd136314880;
      16100: inst = 32'd268468224;
      16101: inst = 32'd201346969;
      16102: inst = 32'd203482053;
      16103: inst = 32'd136314880;
      16104: inst = 32'd268468224;
      16105: inst = 32'd201346970;
      16106: inst = 32'd203479973;
      16107: inst = 32'd136314880;
      16108: inst = 32'd268468224;
      16109: inst = 32'd201346971;
      16110: inst = 32'd203482053;
      16111: inst = 32'd136314880;
      16112: inst = 32'd268468224;
      16113: inst = 32'd201346972;
      16114: inst = 32'd203479973;
      16115: inst = 32'd136314880;
      16116: inst = 32'd268468224;
      16117: inst = 32'd201346973;
      16118: inst = 32'd203482053;
      16119: inst = 32'd136314880;
      16120: inst = 32'd268468224;
      16121: inst = 32'd201346974;
      16122: inst = 32'd203482021;
      16123: inst = 32'd136314880;
      16124: inst = 32'd268468224;
      16125: inst = 32'd201346975;
      16126: inst = 32'd203475682;
      16127: inst = 32'd136314880;
      16128: inst = 32'd268468224;
      16129: inst = 32'd201346976;
      16130: inst = 32'd203459697;
      16131: inst = 32'd136314880;
      16132: inst = 32'd268468224;
      16133: inst = 32'd201346977;
      16134: inst = 32'd203472375;
      16135: inst = 32'd136314880;
      16136: inst = 32'd268468224;
      16137: inst = 32'd201346978;
      16138: inst = 32'd203472343;
      16139: inst = 32'd136314880;
      16140: inst = 32'd268468224;
      16141: inst = 32'd201346979;
      16142: inst = 32'd203472343;
      16143: inst = 32'd136314880;
      16144: inst = 32'd268468224;
      16145: inst = 32'd201346980;
      16146: inst = 32'd203472343;
      16147: inst = 32'd136314880;
      16148: inst = 32'd268468224;
      16149: inst = 32'd201346981;
      16150: inst = 32'd203472375;
      16151: inst = 32'd136314880;
      16152: inst = 32'd268468224;
      16153: inst = 32'd201346982;
      16154: inst = 32'd203472343;
      16155: inst = 32'd136314880;
      16156: inst = 32'd268468224;
      16157: inst = 32'd201346983;
      16158: inst = 32'd203472375;
      16159: inst = 32'd136314880;
      16160: inst = 32'd268468224;
      16161: inst = 32'd201346984;
      16162: inst = 32'd203440647;
      16163: inst = 32'd136314880;
      16164: inst = 32'd268468224;
      16165: inst = 32'd201346985;
      16166: inst = 32'd203472342;
      16167: inst = 32'd136314880;
      16168: inst = 32'd268468224;
      16169: inst = 32'd201346986;
      16170: inst = 32'd203459697;
      16171: inst = 32'd136314880;
      16172: inst = 32'd268468224;
      16173: inst = 32'd201346987;
      16174: inst = 32'd203472342;
      16175: inst = 32'd136314880;
      16176: inst = 32'd268468224;
      16177: inst = 32'd201346988;
      16178: inst = 32'd203440647;
      16179: inst = 32'd136314880;
      16180: inst = 32'd268468224;
      16181: inst = 32'd201346989;
      16182: inst = 32'd203472342;
      16183: inst = 32'd136314880;
      16184: inst = 32'd268468224;
      16185: inst = 32'd201346990;
      16186: inst = 32'd203474423;
      16187: inst = 32'd136314880;
      16188: inst = 32'd268468224;
      16189: inst = 32'd201346991;
      16190: inst = 32'd203472342;
      16191: inst = 32'd136314880;
      16192: inst = 32'd268468224;
      16193: inst = 32'd201346992;
      16194: inst = 32'd203472344;
      16195: inst = 32'd136314880;
      16196: inst = 32'd268468224;
      16197: inst = 32'd201346993;
      16198: inst = 32'd203472375;
      16199: inst = 32'd136314880;
      16200: inst = 32'd268468224;
      16201: inst = 32'd201346994;
      16202: inst = 32'd203472342;
      16203: inst = 32'd136314880;
      16204: inst = 32'd268468224;
      16205: inst = 32'd201346995;
      16206: inst = 32'd203472343;
      16207: inst = 32'd136314880;
      16208: inst = 32'd268468224;
      16209: inst = 32'd201346996;
      16210: inst = 32'd203461714;
      16211: inst = 32'd136314880;
      16212: inst = 32'd268468224;
      16213: inst = 32'd201346997;
      16214: inst = 32'd203453262;
      16215: inst = 32'd136314880;
      16216: inst = 32'd268468224;
      16217: inst = 32'd201346998;
      16218: inst = 32'd203453260;
      16219: inst = 32'd136314880;
      16220: inst = 32'd268468224;
      16221: inst = 32'd201346999;
      16222: inst = 32'd203482839;
      16223: inst = 32'd136314880;
      16224: inst = 32'd268468224;
      16225: inst = 32'd201347000;
      16226: inst = 32'd203484886;
      16227: inst = 32'd136314880;
      16228: inst = 32'd268468224;
      16229: inst = 32'd201347001;
      16230: inst = 32'd203484886;
      16231: inst = 32'd136314880;
      16232: inst = 32'd268468224;
      16233: inst = 32'd201347002;
      16234: inst = 32'd203484822;
      16235: inst = 32'd136314880;
      16236: inst = 32'd268468224;
      16237: inst = 32'd201347003;
      16238: inst = 32'd203484886;
      16239: inst = 32'd136314880;
      16240: inst = 32'd268468224;
      16241: inst = 32'd201347004;
      16242: inst = 32'd203484918;
      16243: inst = 32'd136314880;
      16244: inst = 32'd268468224;
      16245: inst = 32'd201347005;
      16246: inst = 32'd203482806;
      16247: inst = 32'd136314880;
      16248: inst = 32'd268468224;
      16249: inst = 32'd201347006;
      16250: inst = 32'd203484921;
      16251: inst = 32'd136314880;
      16252: inst = 32'd268468224;
      16253: inst = 32'd201347007;
      16254: inst = 32'd203461712;
      16255: inst = 32'd136314880;
      16256: inst = 32'd268468224;
      16257: inst = 32'd201347008;
      16258: inst = 32'd203449069;
      16259: inst = 32'd136314880;
      16260: inst = 32'd268468224;
      16261: inst = 32'd201347009;
      16262: inst = 32'd203449069;
      16263: inst = 32'd136314880;
      16264: inst = 32'd268468224;
      16265: inst = 32'd201347010;
      16266: inst = 32'd203447021;
      16267: inst = 32'd136314880;
      16268: inst = 32'd268468224;
      16269: inst = 32'd201347011;
      16270: inst = 32'd203447021;
      16271: inst = 32'd136314880;
      16272: inst = 32'd268468224;
      16273: inst = 32'd201347012;
      16274: inst = 32'd203449069;
      16275: inst = 32'd136314880;
      16276: inst = 32'd268468224;
      16277: inst = 32'd201347013;
      16278: inst = 32'd203449068;
      16279: inst = 32'd136314880;
      16280: inst = 32'd268468224;
      16281: inst = 32'd201347014;
      16282: inst = 32'd203449035;
      16283: inst = 32'd136314880;
      16284: inst = 32'd268468224;
      16285: inst = 32'd201347015;
      16286: inst = 32'd203449002;
      16287: inst = 32'd136314880;
      16288: inst = 32'd268468224;
      16289: inst = 32'd201347016;
      16290: inst = 32'd203482808;
      16291: inst = 32'd136314880;
      16292: inst = 32'd268468224;
      16293: inst = 32'd201347017;
      16294: inst = 32'd203484855;
      16295: inst = 32'd136314880;
      16296: inst = 32'd268468224;
      16297: inst = 32'd201347018;
      16298: inst = 32'd203482741;
      16299: inst = 32'd136314880;
      16300: inst = 32'd268468224;
      16301: inst = 32'd201347019;
      16302: inst = 32'd203484821;
      16303: inst = 32'd136314880;
      16304: inst = 32'd268468224;
      16305: inst = 32'd201347020;
      16306: inst = 32'd203484853;
      16307: inst = 32'd136314880;
      16308: inst = 32'd268468224;
      16309: inst = 32'd201347021;
      16310: inst = 32'd203484853;
      16311: inst = 32'd136314880;
      16312: inst = 32'd268468224;
      16313: inst = 32'd201347022;
      16314: inst = 32'd203486934;
      16315: inst = 32'd136314880;
      16316: inst = 32'd268468224;
      16317: inst = 32'd201347023;
      16318: inst = 32'd203484854;
      16319: inst = 32'd136314880;
      16320: inst = 32'd268468224;
      16321: inst = 32'd201347024;
      16322: inst = 32'd203484854;
      16323: inst = 32'd136314880;
      16324: inst = 32'd268468224;
      16325: inst = 32'd201347025;
      16326: inst = 32'd203486934;
      16327: inst = 32'd136314880;
      16328: inst = 32'd268468224;
      16329: inst = 32'd201347026;
      16330: inst = 32'd203484853;
      16331: inst = 32'd136314880;
      16332: inst = 32'd268468224;
      16333: inst = 32'd201347027;
      16334: inst = 32'd203484853;
      16335: inst = 32'd136314880;
      16336: inst = 32'd268468224;
      16337: inst = 32'd201347028;
      16338: inst = 32'd203484821;
      16339: inst = 32'd136314880;
      16340: inst = 32'd268468224;
      16341: inst = 32'd201347029;
      16342: inst = 32'd203482741;
      16343: inst = 32'd136314880;
      16344: inst = 32'd268468224;
      16345: inst = 32'd201347030;
      16346: inst = 32'd203484855;
      16347: inst = 32'd136314880;
      16348: inst = 32'd268468224;
      16349: inst = 32'd201347031;
      16350: inst = 32'd203482808;
      16351: inst = 32'd136314880;
      16352: inst = 32'd268468224;
      16353: inst = 32'd201347032;
      16354: inst = 32'd203449002;
      16355: inst = 32'd136314880;
      16356: inst = 32'd268468224;
      16357: inst = 32'd201347033;
      16358: inst = 32'd203449035;
      16359: inst = 32'd136314880;
      16360: inst = 32'd268468224;
      16361: inst = 32'd201347034;
      16362: inst = 32'd203449068;
      16363: inst = 32'd136314880;
      16364: inst = 32'd268468224;
      16365: inst = 32'd201347035;
      16366: inst = 32'd203449069;
      16367: inst = 32'd136314880;
      16368: inst = 32'd268468224;
      16369: inst = 32'd201347036;
      16370: inst = 32'd203447021;
      16371: inst = 32'd136314880;
      16372: inst = 32'd268468224;
      16373: inst = 32'd201347037;
      16374: inst = 32'd203447021;
      16375: inst = 32'd136314880;
      16376: inst = 32'd268468224;
      16377: inst = 32'd201347038;
      16378: inst = 32'd203449069;
      16379: inst = 32'd136314880;
      16380: inst = 32'd268468224;
      16381: inst = 32'd201347039;
      16382: inst = 32'd203449069;
      16383: inst = 32'd136314880;
      16384: inst = 32'd268468224;
      16385: inst = 32'd201347040;
      16386: inst = 32'd203463758;
      16387: inst = 32'd136314880;
      16388: inst = 32'd268468224;
      16389: inst = 32'd201347041;
      16390: inst = 32'd203486967;
      16391: inst = 32'd136314880;
      16392: inst = 32'd268468224;
      16393: inst = 32'd201347042;
      16394: inst = 32'd203484822;
      16395: inst = 32'd136314880;
      16396: inst = 32'd268468224;
      16397: inst = 32'd201347043;
      16398: inst = 32'd203484887;
      16399: inst = 32'd136314880;
      16400: inst = 32'd268468224;
      16401: inst = 32'd201347044;
      16402: inst = 32'd203484855;
      16403: inst = 32'd136314880;
      16404: inst = 32'd268468224;
      16405: inst = 32'd201347045;
      16406: inst = 32'd203484822;
      16407: inst = 32'd136314880;
      16408: inst = 32'd268468224;
      16409: inst = 32'd201347046;
      16410: inst = 32'd203486901;
      16411: inst = 32'd136314880;
      16412: inst = 32'd268468224;
      16413: inst = 32'd201347047;
      16414: inst = 32'd203484854;
      16415: inst = 32'd136314880;
      16416: inst = 32'd268468224;
      16417: inst = 32'd201347048;
      16418: inst = 32'd203484887;
      16419: inst = 32'd136314880;
      16420: inst = 32'd268468224;
      16421: inst = 32'd201347049;
      16422: inst = 32'd203484854;
      16423: inst = 32'd136314880;
      16424: inst = 32'd268468224;
      16425: inst = 32'd201347050;
      16426: inst = 32'd203486901;
      16427: inst = 32'd136314880;
      16428: inst = 32'd268468224;
      16429: inst = 32'd201347051;
      16430: inst = 32'd203484854;
      16431: inst = 32'd136314880;
      16432: inst = 32'd268468224;
      16433: inst = 32'd201347052;
      16434: inst = 32'd203482840;
      16435: inst = 32'd136314880;
      16436: inst = 32'd268468224;
      16437: inst = 32'd201347053;
      16438: inst = 32'd203484856;
      16439: inst = 32'd136314880;
      16440: inst = 32'd268468224;
      16441: inst = 32'd201347054;
      16442: inst = 32'd203488884;
      16443: inst = 32'd136314880;
      16444: inst = 32'd268468224;
      16445: inst = 32'd201347055;
      16446: inst = 32'd203471619;
      16447: inst = 32'd136314880;
      16448: inst = 32'd268468224;
      16449: inst = 32'd201347056;
      16450: inst = 32'd203480006;
      16451: inst = 32'd136314880;
      16452: inst = 32'd268468224;
      16453: inst = 32'd201347057;
      16454: inst = 32'd203480006;
      16455: inst = 32'd136314880;
      16456: inst = 32'd268468224;
      16457: inst = 32'd201347058;
      16458: inst = 32'd203480006;
      16459: inst = 32'd136314880;
      16460: inst = 32'd268468224;
      16461: inst = 32'd201347059;
      16462: inst = 32'd203480006;
      16463: inst = 32'd136314880;
      16464: inst = 32'd268468224;
      16465: inst = 32'd201347060;
      16466: inst = 32'd203480005;
      16467: inst = 32'd136314880;
      16468: inst = 32'd268468224;
      16469: inst = 32'd201347061;
      16470: inst = 32'd203480005;
      16471: inst = 32'd136314880;
      16472: inst = 32'd268468224;
      16473: inst = 32'd201347062;
      16474: inst = 32'd203480005;
      16475: inst = 32'd136314880;
      16476: inst = 32'd268468224;
      16477: inst = 32'd201347063;
      16478: inst = 32'd203480005;
      16479: inst = 32'd136314880;
      16480: inst = 32'd268468224;
      16481: inst = 32'd201347064;
      16482: inst = 32'd203482053;
      16483: inst = 32'd136314880;
      16484: inst = 32'd268468224;
      16485: inst = 32'd201347065;
      16486: inst = 32'd203482053;
      16487: inst = 32'd136314880;
      16488: inst = 32'd268468224;
      16489: inst = 32'd201347066;
      16490: inst = 32'd203479973;
      16491: inst = 32'd136314880;
      16492: inst = 32'd268468224;
      16493: inst = 32'd201347067;
      16494: inst = 32'd203482053;
      16495: inst = 32'd136314880;
      16496: inst = 32'd268468224;
      16497: inst = 32'd201347068;
      16498: inst = 32'd203479973;
      16499: inst = 32'd136314880;
      16500: inst = 32'd268468224;
      16501: inst = 32'd201347069;
      16502: inst = 32'd203482053;
      16503: inst = 32'd136314880;
      16504: inst = 32'd268468224;
      16505: inst = 32'd201347070;
      16506: inst = 32'd203482021;
      16507: inst = 32'd136314880;
      16508: inst = 32'd268468224;
      16509: inst = 32'd201347071;
      16510: inst = 32'd203475682;
      16511: inst = 32'd136314880;
      16512: inst = 32'd268468224;
      16513: inst = 32'd201347072;
      16514: inst = 32'd203459697;
      16515: inst = 32'd136314880;
      16516: inst = 32'd268468224;
      16517: inst = 32'd201347073;
      16518: inst = 32'd203472375;
      16519: inst = 32'd136314880;
      16520: inst = 32'd268468224;
      16521: inst = 32'd201347074;
      16522: inst = 32'd203472343;
      16523: inst = 32'd136314880;
      16524: inst = 32'd268468224;
      16525: inst = 32'd201347075;
      16526: inst = 32'd203472343;
      16527: inst = 32'd136314880;
      16528: inst = 32'd268468224;
      16529: inst = 32'd201347076;
      16530: inst = 32'd203472343;
      16531: inst = 32'd136314880;
      16532: inst = 32'd268468224;
      16533: inst = 32'd201347077;
      16534: inst = 32'd203472375;
      16535: inst = 32'd136314880;
      16536: inst = 32'd268468224;
      16537: inst = 32'd201347078;
      16538: inst = 32'd203472343;
      16539: inst = 32'd136314880;
      16540: inst = 32'd268468224;
      16541: inst = 32'd201347079;
      16542: inst = 32'd203472375;
      16543: inst = 32'd136314880;
      16544: inst = 32'd268468224;
      16545: inst = 32'd201347080;
      16546: inst = 32'd203442793;
      16547: inst = 32'd136314880;
      16548: inst = 32'd268468224;
      16549: inst = 32'd201347081;
      16550: inst = 32'd203472310;
      16551: inst = 32'd136314880;
      16552: inst = 32'd268468224;
      16553: inst = 32'd201347082;
      16554: inst = 32'd203459697;
      16555: inst = 32'd136314880;
      16556: inst = 32'd268468224;
      16557: inst = 32'd201347083;
      16558: inst = 32'd203472342;
      16559: inst = 32'd136314880;
      16560: inst = 32'd268468224;
      16561: inst = 32'd201347084;
      16562: inst = 32'd203444873;
      16563: inst = 32'd136314880;
      16564: inst = 32'd268468224;
      16565: inst = 32'd201347085;
      16566: inst = 32'd203472310;
      16567: inst = 32'd136314880;
      16568: inst = 32'd268468224;
      16569: inst = 32'd201347086;
      16570: inst = 32'd203474423;
      16571: inst = 32'd136314880;
      16572: inst = 32'd268468224;
      16573: inst = 32'd201347087;
      16574: inst = 32'd203472342;
      16575: inst = 32'd136314880;
      16576: inst = 32'd268468224;
      16577: inst = 32'd201347088;
      16578: inst = 32'd203472312;
      16579: inst = 32'd136314880;
      16580: inst = 32'd268468224;
      16581: inst = 32'd201347089;
      16582: inst = 32'd203472344;
      16583: inst = 32'd136314880;
      16584: inst = 32'd268468224;
      16585: inst = 32'd201347090;
      16586: inst = 32'd203472343;
      16587: inst = 32'd136314880;
      16588: inst = 32'd268468224;
      16589: inst = 32'd201347091;
      16590: inst = 32'd203472344;
      16591: inst = 32'd136314880;
      16592: inst = 32'd268468224;
      16593: inst = 32'd201347092;
      16594: inst = 32'd203461715;
      16595: inst = 32'd136314880;
      16596: inst = 32'd268468224;
      16597: inst = 32'd201347093;
      16598: inst = 32'd203453263;
      16599: inst = 32'd136314880;
      16600: inst = 32'd268468224;
      16601: inst = 32'd201347094;
      16602: inst = 32'd203453260;
      16603: inst = 32'd136314880;
      16604: inst = 32'd268468224;
      16605: inst = 32'd201347095;
      16606: inst = 32'd203482839;
      16607: inst = 32'd136314880;
      16608: inst = 32'd268468224;
      16609: inst = 32'd201347096;
      16610: inst = 32'd203482838;
      16611: inst = 32'd136314880;
      16612: inst = 32'd268468224;
      16613: inst = 32'd201347097;
      16614: inst = 32'd203484886;
      16615: inst = 32'd136314880;
      16616: inst = 32'd268468224;
      16617: inst = 32'd201347098;
      16618: inst = 32'd203484854;
      16619: inst = 32'd136314880;
      16620: inst = 32'd268468224;
      16621: inst = 32'd201347099;
      16622: inst = 32'd203484886;
      16623: inst = 32'd136314880;
      16624: inst = 32'd268468224;
      16625: inst = 32'd201347100;
      16626: inst = 32'd203484917;
      16627: inst = 32'd136314880;
      16628: inst = 32'd268468224;
      16629: inst = 32'd201347101;
      16630: inst = 32'd203480725;
      16631: inst = 32'd136314880;
      16632: inst = 32'd268468224;
      16633: inst = 32'd201347102;
      16634: inst = 32'd203482839;
      16635: inst = 32'd136314880;
      16636: inst = 32'd268468224;
      16637: inst = 32'd201347103;
      16638: inst = 32'd203453292;
      16639: inst = 32'd136314880;
      16640: inst = 32'd268468224;
      16641: inst = 32'd201347104;
      16642: inst = 32'd203449100;
      16643: inst = 32'd136314880;
      16644: inst = 32'd268468224;
      16645: inst = 32'd201347105;
      16646: inst = 32'd203449036;
      16647: inst = 32'd136314880;
      16648: inst = 32'd268468224;
      16649: inst = 32'd201347106;
      16650: inst = 32'd203449069;
      16651: inst = 32'd136314880;
      16652: inst = 32'd268468224;
      16653: inst = 32'd201347107;
      16654: inst = 32'd203449102;
      16655: inst = 32'd136314880;
      16656: inst = 32'd268468224;
      16657: inst = 32'd201347108;
      16658: inst = 32'd203446956;
      16659: inst = 32'd136314880;
      16660: inst = 32'd268468224;
      16661: inst = 32'd201347109;
      16662: inst = 32'd203444842;
      16663: inst = 32'd136314880;
      16664: inst = 32'd268468224;
      16665: inst = 32'd201347110;
      16666: inst = 32'd203449035;
      16667: inst = 32'd136314880;
      16668: inst = 32'd268468224;
      16669: inst = 32'd201347111;
      16670: inst = 32'd203453195;
      16671: inst = 32'd136314880;
      16672: inst = 32'd268468224;
      16673: inst = 32'd201347112;
      16674: inst = 32'd203484856;
      16675: inst = 32'd136314880;
      16676: inst = 32'd268468224;
      16677: inst = 32'd201347113;
      16678: inst = 32'd203486935;
      16679: inst = 32'd136314880;
      16680: inst = 32'd268468224;
      16681: inst = 32'd201347114;
      16682: inst = 32'd203486902;
      16683: inst = 32'd136314880;
      16684: inst = 32'd268468224;
      16685: inst = 32'd201347115;
      16686: inst = 32'd203486934;
      16687: inst = 32'd136314880;
      16688: inst = 32'd268468224;
      16689: inst = 32'd201347116;
      16690: inst = 32'd203486869;
      16691: inst = 32'd136314880;
      16692: inst = 32'd268468224;
      16693: inst = 32'd201347117;
      16694: inst = 32'd203484788;
      16695: inst = 32'd136314880;
      16696: inst = 32'd268468224;
      16697: inst = 32'd201347118;
      16698: inst = 32'd203486902;
      16699: inst = 32'd136314880;
      16700: inst = 32'd268468224;
      16701: inst = 32'd201347119;
      16702: inst = 32'd203484821;
      16703: inst = 32'd136314880;
      16704: inst = 32'd268468224;
      16705: inst = 32'd201347120;
      16706: inst = 32'd203484821;
      16707: inst = 32'd136314880;
      16708: inst = 32'd268468224;
      16709: inst = 32'd201347121;
      16710: inst = 32'd203486902;
      16711: inst = 32'd136314880;
      16712: inst = 32'd268468224;
      16713: inst = 32'd201347122;
      16714: inst = 32'd203484788;
      16715: inst = 32'd136314880;
      16716: inst = 32'd268468224;
      16717: inst = 32'd201347123;
      16718: inst = 32'd203486869;
      16719: inst = 32'd136314880;
      16720: inst = 32'd268468224;
      16721: inst = 32'd201347124;
      16722: inst = 32'd203486934;
      16723: inst = 32'd136314880;
      16724: inst = 32'd268468224;
      16725: inst = 32'd201347125;
      16726: inst = 32'd203486902;
      16727: inst = 32'd136314880;
      16728: inst = 32'd268468224;
      16729: inst = 32'd201347126;
      16730: inst = 32'd203486935;
      16731: inst = 32'd136314880;
      16732: inst = 32'd268468224;
      16733: inst = 32'd201347127;
      16734: inst = 32'd203484856;
      16735: inst = 32'd136314880;
      16736: inst = 32'd268468224;
      16737: inst = 32'd201347128;
      16738: inst = 32'd203453195;
      16739: inst = 32'd136314880;
      16740: inst = 32'd268468224;
      16741: inst = 32'd201347129;
      16742: inst = 32'd203449035;
      16743: inst = 32'd136314880;
      16744: inst = 32'd268468224;
      16745: inst = 32'd201347130;
      16746: inst = 32'd203444842;
      16747: inst = 32'd136314880;
      16748: inst = 32'd268468224;
      16749: inst = 32'd201347131;
      16750: inst = 32'd203446956;
      16751: inst = 32'd136314880;
      16752: inst = 32'd268468224;
      16753: inst = 32'd201347132;
      16754: inst = 32'd203449102;
      16755: inst = 32'd136314880;
      16756: inst = 32'd268468224;
      16757: inst = 32'd201347133;
      16758: inst = 32'd203449069;
      16759: inst = 32'd136314880;
      16760: inst = 32'd268468224;
      16761: inst = 32'd201347134;
      16762: inst = 32'd203449036;
      16763: inst = 32'd136314880;
      16764: inst = 32'd268468224;
      16765: inst = 32'd201347135;
      16766: inst = 32'd203449100;
      16767: inst = 32'd136314880;
      16768: inst = 32'd268468224;
      16769: inst = 32'd201347136;
      16770: inst = 32'd203455338;
      16771: inst = 32'd136314880;
      16772: inst = 32'd268468224;
      16773: inst = 32'd201347137;
      16774: inst = 32'd203484855;
      16775: inst = 32'd136314880;
      16776: inst = 32'd268468224;
      16777: inst = 32'd201347138;
      16778: inst = 32'd203482742;
      16779: inst = 32'd136314880;
      16780: inst = 32'd268468224;
      16781: inst = 32'd201347139;
      16782: inst = 32'd203484887;
      16783: inst = 32'd136314880;
      16784: inst = 32'd268468224;
      16785: inst = 32'd201347140;
      16786: inst = 32'd203484888;
      16787: inst = 32'd136314880;
      16788: inst = 32'd268468224;
      16789: inst = 32'd201347141;
      16790: inst = 32'd203484822;
      16791: inst = 32'd136314880;
      16792: inst = 32'd268468224;
      16793: inst = 32'd201347142;
      16794: inst = 32'd203486901;
      16795: inst = 32'd136314880;
      16796: inst = 32'd268468224;
      16797: inst = 32'd201347143;
      16798: inst = 32'd203484854;
      16799: inst = 32'd136314880;
      16800: inst = 32'd268468224;
      16801: inst = 32'd201347144;
      16802: inst = 32'd203484887;
      16803: inst = 32'd136314880;
      16804: inst = 32'd268468224;
      16805: inst = 32'd201347145;
      16806: inst = 32'd203484854;
      16807: inst = 32'd136314880;
      16808: inst = 32'd268468224;
      16809: inst = 32'd201347146;
      16810: inst = 32'd203486901;
      16811: inst = 32'd136314880;
      16812: inst = 32'd268468224;
      16813: inst = 32'd201347147;
      16814: inst = 32'd203484853;
      16815: inst = 32'd136314880;
      16816: inst = 32'd268468224;
      16817: inst = 32'd201347148;
      16818: inst = 32'd203482840;
      16819: inst = 32'd136314880;
      16820: inst = 32'd268468224;
      16821: inst = 32'd201347149;
      16822: inst = 32'd203484856;
      16823: inst = 32'd136314880;
      16824: inst = 32'd268468224;
      16825: inst = 32'd201347150;
      16826: inst = 32'd203488884;
      16827: inst = 32'd136314880;
      16828: inst = 32'd268468224;
      16829: inst = 32'd201347151;
      16830: inst = 32'd203471619;
      16831: inst = 32'd136314880;
      16832: inst = 32'd268468224;
      16833: inst = 32'd201347152;
      16834: inst = 32'd203480006;
      16835: inst = 32'd136314880;
      16836: inst = 32'd268468224;
      16837: inst = 32'd201347153;
      16838: inst = 32'd203480006;
      16839: inst = 32'd136314880;
      16840: inst = 32'd268468224;
      16841: inst = 32'd201347154;
      16842: inst = 32'd203480006;
      16843: inst = 32'd136314880;
      16844: inst = 32'd268468224;
      16845: inst = 32'd201347155;
      16846: inst = 32'd203480005;
      16847: inst = 32'd136314880;
      16848: inst = 32'd268468224;
      16849: inst = 32'd201347156;
      16850: inst = 32'd203480005;
      16851: inst = 32'd136314880;
      16852: inst = 32'd268468224;
      16853: inst = 32'd201347157;
      16854: inst = 32'd203480005;
      16855: inst = 32'd136314880;
      16856: inst = 32'd268468224;
      16857: inst = 32'd201347158;
      16858: inst = 32'd203480005;
      16859: inst = 32'd136314880;
      16860: inst = 32'd268468224;
      16861: inst = 32'd201347159;
      16862: inst = 32'd203480005;
      16863: inst = 32'd136314880;
      16864: inst = 32'd268468224;
      16865: inst = 32'd201347160;
      16866: inst = 32'd203480005;
      16867: inst = 32'd136314880;
      16868: inst = 32'd268468224;
      16869: inst = 32'd201347161;
      16870: inst = 32'd203482053;
      16871: inst = 32'd136314880;
      16872: inst = 32'd268468224;
      16873: inst = 32'd201347162;
      16874: inst = 32'd203479973;
      16875: inst = 32'd136314880;
      16876: inst = 32'd268468224;
      16877: inst = 32'd201347163;
      16878: inst = 32'd203482053;
      16879: inst = 32'd136314880;
      16880: inst = 32'd268468224;
      16881: inst = 32'd201347164;
      16882: inst = 32'd203479973;
      16883: inst = 32'd136314880;
      16884: inst = 32'd268468224;
      16885: inst = 32'd201347165;
      16886: inst = 32'd203482053;
      16887: inst = 32'd136314880;
      16888: inst = 32'd268468224;
      16889: inst = 32'd201347166;
      16890: inst = 32'd203479973;
      16891: inst = 32'd136314880;
      16892: inst = 32'd268468224;
      16893: inst = 32'd201347167;
      16894: inst = 32'd203473634;
      16895: inst = 32'd136314880;
      16896: inst = 32'd268468224;
      16897: inst = 32'd201347168;
      16898: inst = 32'd203459697;
      16899: inst = 32'd136314880;
      16900: inst = 32'd268468224;
      16901: inst = 32'd201347169;
      16902: inst = 32'd203472375;
      16903: inst = 32'd136314880;
      16904: inst = 32'd268468224;
      16905: inst = 32'd201347170;
      16906: inst = 32'd203472343;
      16907: inst = 32'd136314880;
      16908: inst = 32'd268468224;
      16909: inst = 32'd201347171;
      16910: inst = 32'd203472343;
      16911: inst = 32'd136314880;
      16912: inst = 32'd268468224;
      16913: inst = 32'd201347172;
      16914: inst = 32'd203472343;
      16915: inst = 32'd136314880;
      16916: inst = 32'd268468224;
      16917: inst = 32'd201347173;
      16918: inst = 32'd203472375;
      16919: inst = 32'd136314880;
      16920: inst = 32'd268468224;
      16921: inst = 32'd201347174;
      16922: inst = 32'd203472343;
      16923: inst = 32'd136314880;
      16924: inst = 32'd268468224;
      16925: inst = 32'd201347175;
      16926: inst = 32'd203472375;
      16927: inst = 32'd136314880;
      16928: inst = 32'd268468224;
      16929: inst = 32'd201347176;
      16930: inst = 32'd203472342;
      16931: inst = 32'd136314880;
      16932: inst = 32'd268468224;
      16933: inst = 32'd201347177;
      16934: inst = 32'd203472343;
      16935: inst = 32'd136314880;
      16936: inst = 32'd268468224;
      16937: inst = 32'd201347178;
      16938: inst = 32'd203459697;
      16939: inst = 32'd136314880;
      16940: inst = 32'd268468224;
      16941: inst = 32'd201347179;
      16942: inst = 32'd203474455;
      16943: inst = 32'd136314880;
      16944: inst = 32'd268468224;
      16945: inst = 32'd201347180;
      16946: inst = 32'd203470262;
      16947: inst = 32'd136314880;
      16948: inst = 32'd268468224;
      16949: inst = 32'd201347181;
      16950: inst = 32'd203472342;
      16951: inst = 32'd136314880;
      16952: inst = 32'd268468224;
      16953: inst = 32'd201347182;
      16954: inst = 32'd203472375;
      16955: inst = 32'd136314880;
      16956: inst = 32'd268468224;
      16957: inst = 32'd201347183;
      16958: inst = 32'd203472343;
      16959: inst = 32'd136314880;
      16960: inst = 32'd268468224;
      16961: inst = 32'd201347184;
      16962: inst = 32'd203472344;
      16963: inst = 32'd136314880;
      16964: inst = 32'd268468224;
      16965: inst = 32'd201347185;
      16966: inst = 32'd203472376;
      16967: inst = 32'd136314880;
      16968: inst = 32'd268468224;
      16969: inst = 32'd201347186;
      16970: inst = 32'd203472343;
      16971: inst = 32'd136314880;
      16972: inst = 32'd268468224;
      16973: inst = 32'd201347187;
      16974: inst = 32'd203472344;
      16975: inst = 32'd136314880;
      16976: inst = 32'd268468224;
      16977: inst = 32'd201347188;
      16978: inst = 32'd203461715;
      16979: inst = 32'd136314880;
      16980: inst = 32'd268468224;
      16981: inst = 32'd201347189;
      16982: inst = 32'd203453263;
      16983: inst = 32'd136314880;
      16984: inst = 32'd268468224;
      16985: inst = 32'd201347190;
      16986: inst = 32'd203453260;
      16987: inst = 32'd136314880;
      16988: inst = 32'd268468224;
      16989: inst = 32'd201347191;
      16990: inst = 32'd203482839;
      16991: inst = 32'd136314880;
      16992: inst = 32'd268468224;
      16993: inst = 32'd201347192;
      16994: inst = 32'd203482805;
      16995: inst = 32'd136314880;
      16996: inst = 32'd268468224;
      16997: inst = 32'd201347193;
      16998: inst = 32'd203484886;
      16999: inst = 32'd136314880;
      17000: inst = 32'd268468224;
      17001: inst = 32'd201347194;
      17002: inst = 32'd203484854;
      17003: inst = 32'd136314880;
      17004: inst = 32'd268468224;
      17005: inst = 32'd201347195;
      17006: inst = 32'd203484885;
      17007: inst = 32'd136314880;
      17008: inst = 32'd268468224;
      17009: inst = 32'd201347196;
      17010: inst = 32'd203484885;
      17011: inst = 32'd136314880;
      17012: inst = 32'd268468224;
      17013: inst = 32'd201347197;
      17014: inst = 32'd203482837;
      17015: inst = 32'd136314880;
      17016: inst = 32'd268468224;
      17017: inst = 32'd201347198;
      17018: inst = 32'd203482840;
      17019: inst = 32'd136314880;
      17020: inst = 32'd268468224;
      17021: inst = 32'd201347199;
      17022: inst = 32'd203449034;
      17023: inst = 32'd136314880;
      17024: inst = 32'd268468224;
      17025: inst = 32'd201347200;
      17026: inst = 32'd203449100;
      17027: inst = 32'd136314880;
      17028: inst = 32'd268468224;
      17029: inst = 32'd201347201;
      17030: inst = 32'd203449068;
      17031: inst = 32'd136314880;
      17032: inst = 32'd268468224;
      17033: inst = 32'd201347202;
      17034: inst = 32'd203449068;
      17035: inst = 32'd136314880;
      17036: inst = 32'd268468224;
      17037: inst = 32'd201347203;
      17038: inst = 32'd203449101;
      17039: inst = 32'd136314880;
      17040: inst = 32'd268468224;
      17041: inst = 32'd201347204;
      17042: inst = 32'd203444810;
      17043: inst = 32'd136314880;
      17044: inst = 32'd268468224;
      17045: inst = 32'd201347205;
      17046: inst = 32'd203442697;
      17047: inst = 32'd136314880;
      17048: inst = 32'd268468224;
      17049: inst = 32'd201347206;
      17050: inst = 32'd203449035;
      17051: inst = 32'd136314880;
      17052: inst = 32'd268468224;
      17053: inst = 32'd201347207;
      17054: inst = 32'd203453195;
      17055: inst = 32'd136314880;
      17056: inst = 32'd268468224;
      17057: inst = 32'd201347208;
      17058: inst = 32'd203482775;
      17059: inst = 32'd136314880;
      17060: inst = 32'd268468224;
      17061: inst = 32'd201347209;
      17062: inst = 32'd203484822;
      17063: inst = 32'd136314880;
      17064: inst = 32'd268468224;
      17065: inst = 32'd201347210;
      17066: inst = 32'd203486901;
      17067: inst = 32'd136314880;
      17068: inst = 32'd268468224;
      17069: inst = 32'd201347211;
      17070: inst = 32'd203486934;
      17071: inst = 32'd136314880;
      17072: inst = 32'd268468224;
      17073: inst = 32'd201347212;
      17074: inst = 32'd203486901;
      17075: inst = 32'd136314880;
      17076: inst = 32'd268468224;
      17077: inst = 32'd201347213;
      17078: inst = 32'd203486869;
      17079: inst = 32'd136314880;
      17080: inst = 32'd268468224;
      17081: inst = 32'd201347214;
      17082: inst = 32'd203486902;
      17083: inst = 32'd136314880;
      17084: inst = 32'd268468224;
      17085: inst = 32'd201347215;
      17086: inst = 32'd203484821;
      17087: inst = 32'd136314880;
      17088: inst = 32'd268468224;
      17089: inst = 32'd201347216;
      17090: inst = 32'd203484821;
      17091: inst = 32'd136314880;
      17092: inst = 32'd268468224;
      17093: inst = 32'd201347217;
      17094: inst = 32'd203486902;
      17095: inst = 32'd136314880;
      17096: inst = 32'd268468224;
      17097: inst = 32'd201347218;
      17098: inst = 32'd203486869;
      17099: inst = 32'd136314880;
      17100: inst = 32'd268468224;
      17101: inst = 32'd201347219;
      17102: inst = 32'd203486901;
      17103: inst = 32'd136314880;
      17104: inst = 32'd268468224;
      17105: inst = 32'd201347220;
      17106: inst = 32'd203486934;
      17107: inst = 32'd136314880;
      17108: inst = 32'd268468224;
      17109: inst = 32'd201347221;
      17110: inst = 32'd203486901;
      17111: inst = 32'd136314880;
      17112: inst = 32'd268468224;
      17113: inst = 32'd201347222;
      17114: inst = 32'd203484822;
      17115: inst = 32'd136314880;
      17116: inst = 32'd268468224;
      17117: inst = 32'd201347223;
      17118: inst = 32'd203482775;
      17119: inst = 32'd136314880;
      17120: inst = 32'd268468224;
      17121: inst = 32'd201347224;
      17122: inst = 32'd203453195;
      17123: inst = 32'd136314880;
      17124: inst = 32'd268468224;
      17125: inst = 32'd201347225;
      17126: inst = 32'd203449035;
      17127: inst = 32'd136314880;
      17128: inst = 32'd268468224;
      17129: inst = 32'd201347226;
      17130: inst = 32'd203442729;
      17131: inst = 32'd136314880;
      17132: inst = 32'd268468224;
      17133: inst = 32'd201347227;
      17134: inst = 32'd203444843;
      17135: inst = 32'd136314880;
      17136: inst = 32'd268468224;
      17137: inst = 32'd201347228;
      17138: inst = 32'd203449101;
      17139: inst = 32'd136314880;
      17140: inst = 32'd268468224;
      17141: inst = 32'd201347229;
      17142: inst = 32'd203449068;
      17143: inst = 32'd136314880;
      17144: inst = 32'd268468224;
      17145: inst = 32'd201347230;
      17146: inst = 32'd203449068;
      17147: inst = 32'd136314880;
      17148: inst = 32'd268468224;
      17149: inst = 32'd201347231;
      17150: inst = 32'd203449100;
      17151: inst = 32'd136314880;
      17152: inst = 32'd268468224;
      17153: inst = 32'd201347232;
      17154: inst = 32'd203449033;
      17155: inst = 32'd136314880;
      17156: inst = 32'd268468224;
      17157: inst = 32'd201347233;
      17158: inst = 32'd203484855;
      17159: inst = 32'd136314880;
      17160: inst = 32'd268468224;
      17161: inst = 32'd201347234;
      17162: inst = 32'd203484855;
      17163: inst = 32'd136314880;
      17164: inst = 32'd268468224;
      17165: inst = 32'd201347235;
      17166: inst = 32'd203484855;
      17167: inst = 32'd136314880;
      17168: inst = 32'd268468224;
      17169: inst = 32'd201347236;
      17170: inst = 32'd203484855;
      17171: inst = 32'd136314880;
      17172: inst = 32'd268468224;
      17173: inst = 32'd201347237;
      17174: inst = 32'd203484822;
      17175: inst = 32'd136314880;
      17176: inst = 32'd268468224;
      17177: inst = 32'd201347238;
      17178: inst = 32'd203486902;
      17179: inst = 32'd136314880;
      17180: inst = 32'd268468224;
      17181: inst = 32'd201347239;
      17182: inst = 32'd203484854;
      17183: inst = 32'd136314880;
      17184: inst = 32'd268468224;
      17185: inst = 32'd201347240;
      17186: inst = 32'd203484887;
      17187: inst = 32'd136314880;
      17188: inst = 32'd268468224;
      17189: inst = 32'd201347241;
      17190: inst = 32'd203484854;
      17191: inst = 32'd136314880;
      17192: inst = 32'd268468224;
      17193: inst = 32'd201347242;
      17194: inst = 32'd203486901;
      17195: inst = 32'd136314880;
      17196: inst = 32'd268468224;
      17197: inst = 32'd201347243;
      17198: inst = 32'd203484853;
      17199: inst = 32'd136314880;
      17200: inst = 32'd268468224;
      17201: inst = 32'd201347244;
      17202: inst = 32'd203482840;
      17203: inst = 32'd136314880;
      17204: inst = 32'd268468224;
      17205: inst = 32'd201347245;
      17206: inst = 32'd203484856;
      17207: inst = 32'd136314880;
      17208: inst = 32'd268468224;
      17209: inst = 32'd201347246;
      17210: inst = 32'd203488884;
      17211: inst = 32'd136314880;
      17212: inst = 32'd268468224;
      17213: inst = 32'd201347247;
      17214: inst = 32'd203471619;
      17215: inst = 32'd136314880;
      17216: inst = 32'd268468224;
      17217: inst = 32'd201347248;
      17218: inst = 32'd203480006;
      17219: inst = 32'd136314880;
      17220: inst = 32'd268468224;
      17221: inst = 32'd201347249;
      17222: inst = 32'd203480006;
      17223: inst = 32'd136314880;
      17224: inst = 32'd268468224;
      17225: inst = 32'd201347250;
      17226: inst = 32'd203480005;
      17227: inst = 32'd136314880;
      17228: inst = 32'd268468224;
      17229: inst = 32'd201347251;
      17230: inst = 32'd203480005;
      17231: inst = 32'd136314880;
      17232: inst = 32'd268468224;
      17233: inst = 32'd201347252;
      17234: inst = 32'd203480005;
      17235: inst = 32'd136314880;
      17236: inst = 32'd268468224;
      17237: inst = 32'd201347253;
      17238: inst = 32'd203480005;
      17239: inst = 32'd136314880;
      17240: inst = 32'd268468224;
      17241: inst = 32'd201347254;
      17242: inst = 32'd203480005;
      17243: inst = 32'd136314880;
      17244: inst = 32'd268468224;
      17245: inst = 32'd201347255;
      17246: inst = 32'd203480005;
      17247: inst = 32'd136314880;
      17248: inst = 32'd268468224;
      17249: inst = 32'd201347256;
      17250: inst = 32'd203480005;
      17251: inst = 32'd136314880;
      17252: inst = 32'd268468224;
      17253: inst = 32'd201347257;
      17254: inst = 32'd203480005;
      17255: inst = 32'd136314880;
      17256: inst = 32'd268468224;
      17257: inst = 32'd201347258;
      17258: inst = 32'd203479973;
      17259: inst = 32'd136314880;
      17260: inst = 32'd268468224;
      17261: inst = 32'd201347259;
      17262: inst = 32'd203482053;
      17263: inst = 32'd136314880;
      17264: inst = 32'd268468224;
      17265: inst = 32'd201347260;
      17266: inst = 32'd203479973;
      17267: inst = 32'd136314880;
      17268: inst = 32'd268468224;
      17269: inst = 32'd201347261;
      17270: inst = 32'd203482053;
      17271: inst = 32'd136314880;
      17272: inst = 32'd268468224;
      17273: inst = 32'd201347262;
      17274: inst = 32'd203479973;
      17275: inst = 32'd136314880;
      17276: inst = 32'd268468224;
      17277: inst = 32'd201347263;
      17278: inst = 32'd203473634;
      17279: inst = 32'd136314880;
      17280: inst = 32'd268468224;
      17281: inst = 32'd201347264;
      17282: inst = 32'd203459697;
      17283: inst = 32'd136314880;
      17284: inst = 32'd268468224;
      17285: inst = 32'd201347265;
      17286: inst = 32'd203472375;
      17287: inst = 32'd136314880;
      17288: inst = 32'd268468224;
      17289: inst = 32'd201347266;
      17290: inst = 32'd203472375;
      17291: inst = 32'd136314880;
      17292: inst = 32'd268468224;
      17293: inst = 32'd201347267;
      17294: inst = 32'd203472375;
      17295: inst = 32'd136314880;
      17296: inst = 32'd268468224;
      17297: inst = 32'd201347268;
      17298: inst = 32'd203472375;
      17299: inst = 32'd136314880;
      17300: inst = 32'd268468224;
      17301: inst = 32'd201347269;
      17302: inst = 32'd203472375;
      17303: inst = 32'd136314880;
      17304: inst = 32'd268468224;
      17305: inst = 32'd201347270;
      17306: inst = 32'd203472343;
      17307: inst = 32'd136314880;
      17308: inst = 32'd268468224;
      17309: inst = 32'd201347271;
      17310: inst = 32'd203472375;
      17311: inst = 32'd136314880;
      17312: inst = 32'd268468224;
      17313: inst = 32'd201347272;
      17314: inst = 32'd203472343;
      17315: inst = 32'd136314880;
      17316: inst = 32'd268468224;
      17317: inst = 32'd201347273;
      17318: inst = 32'd203472375;
      17319: inst = 32'd136314880;
      17320: inst = 32'd268468224;
      17321: inst = 32'd201347274;
      17322: inst = 32'd203459665;
      17323: inst = 32'd136314880;
      17324: inst = 32'd268468224;
      17325: inst = 32'd201347275;
      17326: inst = 32'd203472343;
      17327: inst = 32'd136314880;
      17328: inst = 32'd268468224;
      17329: inst = 32'd201347276;
      17330: inst = 32'd203472375;
      17331: inst = 32'd136314880;
      17332: inst = 32'd268468224;
      17333: inst = 32'd201347277;
      17334: inst = 32'd203472375;
      17335: inst = 32'd136314880;
      17336: inst = 32'd268468224;
      17337: inst = 32'd201347278;
      17338: inst = 32'd203472343;
      17339: inst = 32'd136314880;
      17340: inst = 32'd268468224;
      17341: inst = 32'd201347279;
      17342: inst = 32'd203472375;
      17343: inst = 32'd136314880;
      17344: inst = 32'd268468224;
      17345: inst = 32'd201347280;
      17346: inst = 32'd203472343;
      17347: inst = 32'd136314880;
      17348: inst = 32'd268468224;
      17349: inst = 32'd201347281;
      17350: inst = 32'd203472375;
      17351: inst = 32'd136314880;
      17352: inst = 32'd268468224;
      17353: inst = 32'd201347282;
      17354: inst = 32'd203472342;
      17355: inst = 32'd136314880;
      17356: inst = 32'd268468224;
      17357: inst = 32'd201347283;
      17358: inst = 32'd203472375;
      17359: inst = 32'd136314880;
      17360: inst = 32'd268468224;
      17361: inst = 32'd201347284;
      17362: inst = 32'd203461714;
      17363: inst = 32'd136314880;
      17364: inst = 32'd268468224;
      17365: inst = 32'd201347285;
      17366: inst = 32'd203453262;
      17367: inst = 32'd136314880;
      17368: inst = 32'd268468224;
      17369: inst = 32'd201347286;
      17370: inst = 32'd203453260;
      17371: inst = 32'd136314880;
      17372: inst = 32'd268468224;
      17373: inst = 32'd201347287;
      17374: inst = 32'd203482839;
      17375: inst = 32'd136314880;
      17376: inst = 32'd268468224;
      17377: inst = 32'd201347288;
      17378: inst = 32'd203484853;
      17379: inst = 32'd136314880;
      17380: inst = 32'd268468224;
      17381: inst = 32'd201347289;
      17382: inst = 32'd203484886;
      17383: inst = 32'd136314880;
      17384: inst = 32'd268468224;
      17385: inst = 32'd201347290;
      17386: inst = 32'd203484854;
      17387: inst = 32'd136314880;
      17388: inst = 32'd268468224;
      17389: inst = 32'd201347291;
      17390: inst = 32'd203484821;
      17391: inst = 32'd136314880;
      17392: inst = 32'd268468224;
      17393: inst = 32'd201347292;
      17394: inst = 32'd203484853;
      17395: inst = 32'd136314880;
      17396: inst = 32'd268468224;
      17397: inst = 32'd201347293;
      17398: inst = 32'd203484919;
      17399: inst = 32'd136314880;
      17400: inst = 32'd268468224;
      17401: inst = 32'd201347294;
      17402: inst = 32'd203484888;
      17403: inst = 32'd136314880;
      17404: inst = 32'd268468224;
      17405: inst = 32'd201347295;
      17406: inst = 32'd203451083;
      17407: inst = 32'd136314880;
      17408: inst = 32'd268468224;
      17409: inst = 32'd201347296;
      17410: inst = 32'd203447019;
      17411: inst = 32'd136314880;
      17412: inst = 32'd268468224;
      17413: inst = 32'd201347297;
      17414: inst = 32'd203449132;
      17415: inst = 32'd136314880;
      17416: inst = 32'd268468224;
      17417: inst = 32'd201347298;
      17418: inst = 32'd203447020;
      17419: inst = 32'd136314880;
      17420: inst = 32'd268468224;
      17421: inst = 32'd201347299;
      17422: inst = 32'd203444907;
      17423: inst = 32'd136314880;
      17424: inst = 32'd268468224;
      17425: inst = 32'd201347300;
      17426: inst = 32'd203442762;
      17427: inst = 32'd136314880;
      17428: inst = 32'd268468224;
      17429: inst = 32'd201347301;
      17430: inst = 32'd203442794;
      17431: inst = 32'd136314880;
      17432: inst = 32'd268468224;
      17433: inst = 32'd201347302;
      17434: inst = 32'd203451148;
      17435: inst = 32'd136314880;
      17436: inst = 32'd268468224;
      17437: inst = 32'd201347303;
      17438: inst = 32'd203449034;
      17439: inst = 32'd136314880;
      17440: inst = 32'd268468224;
      17441: inst = 32'd201347304;
      17442: inst = 32'd203487001;
      17443: inst = 32'd136314880;
      17444: inst = 32'd268468224;
      17445: inst = 32'd201347305;
      17446: inst = 32'd203482774;
      17447: inst = 32'd136314880;
      17448: inst = 32'd268468224;
      17449: inst = 32'd201347306;
      17450: inst = 32'd203484854;
      17451: inst = 32'd136314880;
      17452: inst = 32'd268468224;
      17453: inst = 32'd201347307;
      17454: inst = 32'd203484853;
      17455: inst = 32'd136314880;
      17456: inst = 32'd268468224;
      17457: inst = 32'd201347308;
      17458: inst = 32'd203484821;
      17459: inst = 32'd136314880;
      17460: inst = 32'd268468224;
      17461: inst = 32'd201347309;
      17462: inst = 32'd203486935;
      17463: inst = 32'd136314880;
      17464: inst = 32'd268468224;
      17465: inst = 32'd201347310;
      17466: inst = 32'd203486903;
      17467: inst = 32'd136314880;
      17468: inst = 32'd268468224;
      17469: inst = 32'd201347311;
      17470: inst = 32'd203484823;
      17471: inst = 32'd136314880;
      17472: inst = 32'd268468224;
      17473: inst = 32'd201347312;
      17474: inst = 32'd203484823;
      17475: inst = 32'd136314880;
      17476: inst = 32'd268468224;
      17477: inst = 32'd201347313;
      17478: inst = 32'd203486903;
      17479: inst = 32'd136314880;
      17480: inst = 32'd268468224;
      17481: inst = 32'd201347314;
      17482: inst = 32'd203486935;
      17483: inst = 32'd136314880;
      17484: inst = 32'd268468224;
      17485: inst = 32'd201347315;
      17486: inst = 32'd203484821;
      17487: inst = 32'd136314880;
      17488: inst = 32'd268468224;
      17489: inst = 32'd201347316;
      17490: inst = 32'd203484853;
      17491: inst = 32'd136314880;
      17492: inst = 32'd268468224;
      17493: inst = 32'd201347317;
      17494: inst = 32'd203484854;
      17495: inst = 32'd136314880;
      17496: inst = 32'd268468224;
      17497: inst = 32'd201347318;
      17498: inst = 32'd203482774;
      17499: inst = 32'd136314880;
      17500: inst = 32'd268468224;
      17501: inst = 32'd201347319;
      17502: inst = 32'd203487001;
      17503: inst = 32'd136314880;
      17504: inst = 32'd268468224;
      17505: inst = 32'd201347320;
      17506: inst = 32'd203449034;
      17507: inst = 32'd136314880;
      17508: inst = 32'd268468224;
      17509: inst = 32'd201347321;
      17510: inst = 32'd203451148;
      17511: inst = 32'd136314880;
      17512: inst = 32'd268468224;
      17513: inst = 32'd201347322;
      17514: inst = 32'd203444842;
      17515: inst = 32'd136314880;
      17516: inst = 32'd268468224;
      17517: inst = 32'd201347323;
      17518: inst = 32'd203442762;
      17519: inst = 32'd136314880;
      17520: inst = 32'd268468224;
      17521: inst = 32'd201347324;
      17522: inst = 32'd203444907;
      17523: inst = 32'd136314880;
      17524: inst = 32'd268468224;
      17525: inst = 32'd201347325;
      17526: inst = 32'd203446988;
      17527: inst = 32'd136314880;
      17528: inst = 32'd268468224;
      17529: inst = 32'd201347326;
      17530: inst = 32'd203449132;
      17531: inst = 32'd136314880;
      17532: inst = 32'd268468224;
      17533: inst = 32'd201347327;
      17534: inst = 32'd203447019;
      17535: inst = 32'd136314880;
      17536: inst = 32'd268468224;
      17537: inst = 32'd201347328;
      17538: inst = 32'd203449065;
      17539: inst = 32'd136314880;
      17540: inst = 32'd268468224;
      17541: inst = 32'd201347329;
      17542: inst = 32'd203484888;
      17543: inst = 32'd136314880;
      17544: inst = 32'd268468224;
      17545: inst = 32'd201347330;
      17546: inst = 32'd203484888;
      17547: inst = 32'd136314880;
      17548: inst = 32'd268468224;
      17549: inst = 32'd201347331;
      17550: inst = 32'd203482807;
      17551: inst = 32'd136314880;
      17552: inst = 32'd268468224;
      17553: inst = 32'd201347332;
      17554: inst = 32'd203482775;
      17555: inst = 32'd136314880;
      17556: inst = 32'd268468224;
      17557: inst = 32'd201347333;
      17558: inst = 32'd203484854;
      17559: inst = 32'd136314880;
      17560: inst = 32'd268468224;
      17561: inst = 32'd201347334;
      17562: inst = 32'd203486902;
      17563: inst = 32'd136314880;
      17564: inst = 32'd268468224;
      17565: inst = 32'd201347335;
      17566: inst = 32'd203484854;
      17567: inst = 32'd136314880;
      17568: inst = 32'd268468224;
      17569: inst = 32'd201347336;
      17570: inst = 32'd203484887;
      17571: inst = 32'd136314880;
      17572: inst = 32'd268468224;
      17573: inst = 32'd201347337;
      17574: inst = 32'd203484854;
      17575: inst = 32'd136314880;
      17576: inst = 32'd268468224;
      17577: inst = 32'd201347338;
      17578: inst = 32'd203486901;
      17579: inst = 32'd136314880;
      17580: inst = 32'd268468224;
      17581: inst = 32'd201347339;
      17582: inst = 32'd203484853;
      17583: inst = 32'd136314880;
      17584: inst = 32'd268468224;
      17585: inst = 32'd201347340;
      17586: inst = 32'd203482840;
      17587: inst = 32'd136314880;
      17588: inst = 32'd268468224;
      17589: inst = 32'd201347341;
      17590: inst = 32'd203484856;
      17591: inst = 32'd136314880;
      17592: inst = 32'd268468224;
      17593: inst = 32'd201347342;
      17594: inst = 32'd203488884;
      17595: inst = 32'd136314880;
      17596: inst = 32'd268468224;
      17597: inst = 32'd201347343;
      17598: inst = 32'd203471619;
      17599: inst = 32'd136314880;
      17600: inst = 32'd268468224;
      17601: inst = 32'd201347344;
      17602: inst = 32'd203480005;
      17603: inst = 32'd136314880;
      17604: inst = 32'd268468224;
      17605: inst = 32'd201347345;
      17606: inst = 32'd203480005;
      17607: inst = 32'd136314880;
      17608: inst = 32'd268468224;
      17609: inst = 32'd201347346;
      17610: inst = 32'd203480005;
      17611: inst = 32'd136314880;
      17612: inst = 32'd268468224;
      17613: inst = 32'd201347347;
      17614: inst = 32'd203480005;
      17615: inst = 32'd136314880;
      17616: inst = 32'd268468224;
      17617: inst = 32'd201347348;
      17618: inst = 32'd203480005;
      17619: inst = 32'd136314880;
      17620: inst = 32'd268468224;
      17621: inst = 32'd201347349;
      17622: inst = 32'd203480005;
      17623: inst = 32'd136314880;
      17624: inst = 32'd268468224;
      17625: inst = 32'd201347350;
      17626: inst = 32'd203480005;
      17627: inst = 32'd136314880;
      17628: inst = 32'd268468224;
      17629: inst = 32'd201347351;
      17630: inst = 32'd203480005;
      17631: inst = 32'd136314880;
      17632: inst = 32'd268468224;
      17633: inst = 32'd201347352;
      17634: inst = 32'd203480005;
      17635: inst = 32'd136314880;
      17636: inst = 32'd268468224;
      17637: inst = 32'd201347353;
      17638: inst = 32'd203480005;
      17639: inst = 32'd136314880;
      17640: inst = 32'd268468224;
      17641: inst = 32'd201347354;
      17642: inst = 32'd203479973;
      17643: inst = 32'd136314880;
      17644: inst = 32'd268468224;
      17645: inst = 32'd201347355;
      17646: inst = 32'd203480005;
      17647: inst = 32'd136314880;
      17648: inst = 32'd268468224;
      17649: inst = 32'd201347356;
      17650: inst = 32'd203479973;
      17651: inst = 32'd136314880;
      17652: inst = 32'd268468224;
      17653: inst = 32'd201347357;
      17654: inst = 32'd203480005;
      17655: inst = 32'd136314880;
      17656: inst = 32'd268468224;
      17657: inst = 32'd201347358;
      17658: inst = 32'd203479973;
      17659: inst = 32'd136314880;
      17660: inst = 32'd268468224;
      17661: inst = 32'd201347359;
      17662: inst = 32'd203473634;
      17663: inst = 32'd136314880;
      17664: inst = 32'd268468224;
      17665: inst = 32'd201347360;
      17666: inst = 32'd203459697;
      17667: inst = 32'd136314880;
      17668: inst = 32'd268468224;
      17669: inst = 32'd201347361;
      17670: inst = 32'd203472375;
      17671: inst = 32'd136314880;
      17672: inst = 32'd268468224;
      17673: inst = 32'd201347362;
      17674: inst = 32'd203472375;
      17675: inst = 32'd136314880;
      17676: inst = 32'd268468224;
      17677: inst = 32'd201347363;
      17678: inst = 32'd203472375;
      17679: inst = 32'd136314880;
      17680: inst = 32'd268468224;
      17681: inst = 32'd201347364;
      17682: inst = 32'd203472375;
      17683: inst = 32'd136314880;
      17684: inst = 32'd268468224;
      17685: inst = 32'd201347365;
      17686: inst = 32'd203472375;
      17687: inst = 32'd136314880;
      17688: inst = 32'd268468224;
      17689: inst = 32'd201347366;
      17690: inst = 32'd203472375;
      17691: inst = 32'd136314880;
      17692: inst = 32'd268468224;
      17693: inst = 32'd201347367;
      17694: inst = 32'd203472375;
      17695: inst = 32'd136314880;
      17696: inst = 32'd268468224;
      17697: inst = 32'd201347368;
      17698: inst = 32'd203472375;
      17699: inst = 32'd136314880;
      17700: inst = 32'd268468224;
      17701: inst = 32'd201347369;
      17702: inst = 32'd203472343;
      17703: inst = 32'd136314880;
      17704: inst = 32'd268468224;
      17705: inst = 32'd201347370;
      17706: inst = 32'd203459729;
      17707: inst = 32'd136314880;
      17708: inst = 32'd268468224;
      17709: inst = 32'd201347371;
      17710: inst = 32'd203470262;
      17711: inst = 32'd136314880;
      17712: inst = 32'd268468224;
      17713: inst = 32'd201347372;
      17714: inst = 32'd203474456;
      17715: inst = 32'd136314880;
      17716: inst = 32'd268468224;
      17717: inst = 32'd201347373;
      17718: inst = 32'd203470295;
      17719: inst = 32'd136314880;
      17720: inst = 32'd268468224;
      17721: inst = 32'd201347374;
      17722: inst = 32'd203472408;
      17723: inst = 32'd136314880;
      17724: inst = 32'd268468224;
      17725: inst = 32'd201347375;
      17726: inst = 32'd203470295;
      17727: inst = 32'd136314880;
      17728: inst = 32'd268468224;
      17729: inst = 32'd201347376;
      17730: inst = 32'd203470327;
      17731: inst = 32'd136314880;
      17732: inst = 32'd268468224;
      17733: inst = 32'd201347377;
      17734: inst = 32'd203472406;
      17735: inst = 32'd136314880;
      17736: inst = 32'd268468224;
      17737: inst = 32'd201347378;
      17738: inst = 32'd203470325;
      17739: inst = 32'd136314880;
      17740: inst = 32'd268468224;
      17741: inst = 32'd201347379;
      17742: inst = 32'd203472375;
      17743: inst = 32'd136314880;
      17744: inst = 32'd268468224;
      17745: inst = 32'd201347380;
      17746: inst = 32'd203459666;
      17747: inst = 32'd136314880;
      17748: inst = 32'd268468224;
      17749: inst = 32'd201347381;
      17750: inst = 32'd203453294;
      17751: inst = 32'd136314880;
      17752: inst = 32'd268468224;
      17753: inst = 32'd201347382;
      17754: inst = 32'd203453260;
      17755: inst = 32'd136314880;
      17756: inst = 32'd268468224;
      17757: inst = 32'd201347383;
      17758: inst = 32'd203482839;
      17759: inst = 32'd136314880;
      17760: inst = 32'd268468224;
      17761: inst = 32'd201347384;
      17762: inst = 32'd203484886;
      17763: inst = 32'd136314880;
      17764: inst = 32'd268468224;
      17765: inst = 32'd201347385;
      17766: inst = 32'd203484853;
      17767: inst = 32'd136314880;
      17768: inst = 32'd268468224;
      17769: inst = 32'd201347386;
      17770: inst = 32'd203486934;
      17771: inst = 32'd136314880;
      17772: inst = 32'd268468224;
      17773: inst = 32'd201347387;
      17774: inst = 32'd203484822;
      17775: inst = 32'd136314880;
      17776: inst = 32'd268468224;
      17777: inst = 32'd201347388;
      17778: inst = 32'd203484854;
      17779: inst = 32'd136314880;
      17780: inst = 32'd268468224;
      17781: inst = 32'd201347389;
      17782: inst = 32'd203484887;
      17783: inst = 32'd136314880;
      17784: inst = 32'd268468224;
      17785: inst = 32'd201347390;
      17786: inst = 32'd203482744;
      17787: inst = 32'd136314880;
      17788: inst = 32'd268468224;
      17789: inst = 32'd201347391;
      17790: inst = 32'd203453132;
      17791: inst = 32'd136314880;
      17792: inst = 32'd268468224;
      17793: inst = 32'd201347392;
      17794: inst = 32'd203447019;
      17795: inst = 32'd136314880;
      17796: inst = 32'd268468224;
      17797: inst = 32'd201347393;
      17798: inst = 32'd203447084;
      17799: inst = 32'd136314880;
      17800: inst = 32'd268468224;
      17801: inst = 32'd201347394;
      17802: inst = 32'd203444907;
      17803: inst = 32'd136314880;
      17804: inst = 32'd268468224;
      17805: inst = 32'd201347395;
      17806: inst = 32'd203442827;
      17807: inst = 32'd136314880;
      17808: inst = 32'd268468224;
      17809: inst = 32'd201347396;
      17810: inst = 32'd203442795;
      17811: inst = 32'd136314880;
      17812: inst = 32'd268468224;
      17813: inst = 32'd201347397;
      17814: inst = 32'd203444907;
      17815: inst = 32'd136314880;
      17816: inst = 32'd268468224;
      17817: inst = 32'd201347398;
      17818: inst = 32'd203451181;
      17819: inst = 32'd136314880;
      17820: inst = 32'd268468224;
      17821: inst = 32'd201347399;
      17822: inst = 32'd203449034;
      17823: inst = 32'd136314880;
      17824: inst = 32'd268468224;
      17825: inst = 32'd201347400;
      17826: inst = 32'd203482841;
      17827: inst = 32'd136314880;
      17828: inst = 32'd268468224;
      17829: inst = 32'd201347401;
      17830: inst = 32'd203480662;
      17831: inst = 32'd136314880;
      17832: inst = 32'd268468224;
      17833: inst = 32'd201347402;
      17834: inst = 32'd203487000;
      17835: inst = 32'd136314880;
      17836: inst = 32'd268468224;
      17837: inst = 32'd201347403;
      17838: inst = 32'd203484887;
      17839: inst = 32'd136314880;
      17840: inst = 32'd268468224;
      17841: inst = 32'd201347404;
      17842: inst = 32'd203482774;
      17843: inst = 32'd136314880;
      17844: inst = 32'd268468224;
      17845: inst = 32'd201347405;
      17846: inst = 32'd203486935;
      17847: inst = 32'd136314880;
      17848: inst = 32'd268468224;
      17849: inst = 32'd201347406;
      17850: inst = 32'd203482775;
      17851: inst = 32'd136314880;
      17852: inst = 32'd268468224;
      17853: inst = 32'd201347407;
      17854: inst = 32'd203484855;
      17855: inst = 32'd136314880;
      17856: inst = 32'd268468224;
      17857: inst = 32'd201347408;
      17858: inst = 32'd203484855;
      17859: inst = 32'd136314880;
      17860: inst = 32'd268468224;
      17861: inst = 32'd201347409;
      17862: inst = 32'd203482775;
      17863: inst = 32'd136314880;
      17864: inst = 32'd268468224;
      17865: inst = 32'd201347410;
      17866: inst = 32'd203486935;
      17867: inst = 32'd136314880;
      17868: inst = 32'd268468224;
      17869: inst = 32'd201347411;
      17870: inst = 32'd203482774;
      17871: inst = 32'd136314880;
      17872: inst = 32'd268468224;
      17873: inst = 32'd201347412;
      17874: inst = 32'd203484887;
      17875: inst = 32'd136314880;
      17876: inst = 32'd268468224;
      17877: inst = 32'd201347413;
      17878: inst = 32'd203487000;
      17879: inst = 32'd136314880;
      17880: inst = 32'd268468224;
      17881: inst = 32'd201347414;
      17882: inst = 32'd203480662;
      17883: inst = 32'd136314880;
      17884: inst = 32'd268468224;
      17885: inst = 32'd201347415;
      17886: inst = 32'd203482841;
      17887: inst = 32'd136314880;
      17888: inst = 32'd268468224;
      17889: inst = 32'd201347416;
      17890: inst = 32'd203449034;
      17891: inst = 32'd136314880;
      17892: inst = 32'd268468224;
      17893: inst = 32'd201347417;
      17894: inst = 32'd203451181;
      17895: inst = 32'd136314880;
      17896: inst = 32'd268468224;
      17897: inst = 32'd201347418;
      17898: inst = 32'd203444907;
      17899: inst = 32'd136314880;
      17900: inst = 32'd268468224;
      17901: inst = 32'd201347419;
      17902: inst = 32'd203442795;
      17903: inst = 32'd136314880;
      17904: inst = 32'd268468224;
      17905: inst = 32'd201347420;
      17906: inst = 32'd203442827;
      17907: inst = 32'd136314880;
      17908: inst = 32'd268468224;
      17909: inst = 32'd201347421;
      17910: inst = 32'd203444907;
      17911: inst = 32'd136314880;
      17912: inst = 32'd268468224;
      17913: inst = 32'd201347422;
      17914: inst = 32'd203447084;
      17915: inst = 32'd136314880;
      17916: inst = 32'd268468224;
      17917: inst = 32'd201347423;
      17918: inst = 32'd203447019;
      17919: inst = 32'd136314880;
      17920: inst = 32'd268468224;
      17921: inst = 32'd201347424;
      17922: inst = 32'd203451146;
      17923: inst = 32'd136314880;
      17924: inst = 32'd268468224;
      17925: inst = 32'd201347425;
      17926: inst = 32'd203480695;
      17927: inst = 32'd136314880;
      17928: inst = 32'd268468224;
      17929: inst = 32'd201347426;
      17930: inst = 32'd203484888;
      17931: inst = 32'd136314880;
      17932: inst = 32'd268468224;
      17933: inst = 32'd201347427;
      17934: inst = 32'd203482808;
      17935: inst = 32'd136314880;
      17936: inst = 32'd268468224;
      17937: inst = 32'd201347428;
      17938: inst = 32'd203482775;
      17939: inst = 32'd136314880;
      17940: inst = 32'd268468224;
      17941: inst = 32'd201347429;
      17942: inst = 32'd203486935;
      17943: inst = 32'd136314880;
      17944: inst = 32'd268468224;
      17945: inst = 32'd201347430;
      17946: inst = 32'd203484821;
      17947: inst = 32'd136314880;
      17948: inst = 32'd268468224;
      17949: inst = 32'd201347431;
      17950: inst = 32'd203484854;
      17951: inst = 32'd136314880;
      17952: inst = 32'd268468224;
      17953: inst = 32'd201347432;
      17954: inst = 32'd203484887;
      17955: inst = 32'd136314880;
      17956: inst = 32'd268468224;
      17957: inst = 32'd201347433;
      17958: inst = 32'd203484854;
      17959: inst = 32'd136314880;
      17960: inst = 32'd268468224;
      17961: inst = 32'd201347434;
      17962: inst = 32'd203486901;
      17963: inst = 32'd136314880;
      17964: inst = 32'd268468224;
      17965: inst = 32'd201347435;
      17966: inst = 32'd203484853;
      17967: inst = 32'd136314880;
      17968: inst = 32'd268468224;
      17969: inst = 32'd201347436;
      17970: inst = 32'd203482840;
      17971: inst = 32'd136314880;
      17972: inst = 32'd268468224;
      17973: inst = 32'd201347437;
      17974: inst = 32'd203484856;
      17975: inst = 32'd136314880;
      17976: inst = 32'd268468224;
      17977: inst = 32'd201347438;
      17978: inst = 32'd203488884;
      17979: inst = 32'd136314880;
      17980: inst = 32'd268468224;
      17981: inst = 32'd201347439;
      17982: inst = 32'd203471619;
      17983: inst = 32'd136314880;
      17984: inst = 32'd268468224;
      17985: inst = 32'd201347440;
      17986: inst = 32'd203480005;
      17987: inst = 32'd136314880;
      17988: inst = 32'd268468224;
      17989: inst = 32'd201347441;
      17990: inst = 32'd203480005;
      17991: inst = 32'd136314880;
      17992: inst = 32'd268468224;
      17993: inst = 32'd201347442;
      17994: inst = 32'd203480005;
      17995: inst = 32'd136314880;
      17996: inst = 32'd268468224;
      17997: inst = 32'd201347443;
      17998: inst = 32'd203480005;
      17999: inst = 32'd136314880;
      18000: inst = 32'd268468224;
      18001: inst = 32'd201347444;
      18002: inst = 32'd203480005;
      18003: inst = 32'd136314880;
      18004: inst = 32'd268468224;
      18005: inst = 32'd201347445;
      18006: inst = 32'd203480005;
      18007: inst = 32'd136314880;
      18008: inst = 32'd268468224;
      18009: inst = 32'd201347446;
      18010: inst = 32'd203480005;
      18011: inst = 32'd136314880;
      18012: inst = 32'd268468224;
      18013: inst = 32'd201347447;
      18014: inst = 32'd203480005;
      18015: inst = 32'd136314880;
      18016: inst = 32'd268468224;
      18017: inst = 32'd201347448;
      18018: inst = 32'd203480005;
      18019: inst = 32'd136314880;
      18020: inst = 32'd268468224;
      18021: inst = 32'd201347449;
      18022: inst = 32'd203480005;
      18023: inst = 32'd136314880;
      18024: inst = 32'd268468224;
      18025: inst = 32'd201347450;
      18026: inst = 32'd203479973;
      18027: inst = 32'd136314880;
      18028: inst = 32'd268468224;
      18029: inst = 32'd201347451;
      18030: inst = 32'd203480005;
      18031: inst = 32'd136314880;
      18032: inst = 32'd268468224;
      18033: inst = 32'd201347452;
      18034: inst = 32'd203479973;
      18035: inst = 32'd136314880;
      18036: inst = 32'd268468224;
      18037: inst = 32'd201347453;
      18038: inst = 32'd203480005;
      18039: inst = 32'd136314880;
      18040: inst = 32'd268468224;
      18041: inst = 32'd201347454;
      18042: inst = 32'd203479973;
      18043: inst = 32'd136314880;
      18044: inst = 32'd268468224;
      18045: inst = 32'd201347455;
      18046: inst = 32'd203473634;
      18047: inst = 32'd136314880;
      18048: inst = 32'd268468224;
      18049: inst = 32'd201347456;
      18050: inst = 32'd203459697;
      18051: inst = 32'd136314880;
      18052: inst = 32'd268468224;
      18053: inst = 32'd201347457;
      18054: inst = 32'd203472375;
      18055: inst = 32'd136314880;
      18056: inst = 32'd268468224;
      18057: inst = 32'd201347458;
      18058: inst = 32'd203472375;
      18059: inst = 32'd136314880;
      18060: inst = 32'd268468224;
      18061: inst = 32'd201347459;
      18062: inst = 32'd203472375;
      18063: inst = 32'd136314880;
      18064: inst = 32'd268468224;
      18065: inst = 32'd201347460;
      18066: inst = 32'd203472375;
      18067: inst = 32'd136314880;
      18068: inst = 32'd268468224;
      18069: inst = 32'd201347461;
      18070: inst = 32'd203472375;
      18071: inst = 32'd136314880;
      18072: inst = 32'd268468224;
      18073: inst = 32'd201347462;
      18074: inst = 32'd203472375;
      18075: inst = 32'd136314880;
      18076: inst = 32'd268468224;
      18077: inst = 32'd201347463;
      18078: inst = 32'd203472375;
      18079: inst = 32'd136314880;
      18080: inst = 32'd268468224;
      18081: inst = 32'd201347464;
      18082: inst = 32'd203472343;
      18083: inst = 32'd136314880;
      18084: inst = 32'd268468224;
      18085: inst = 32'd201347465;
      18086: inst = 32'd203472343;
      18087: inst = 32'd136314880;
      18088: inst = 32'd268468224;
      18089: inst = 32'd201347466;
      18090: inst = 32'd203459729;
      18091: inst = 32'd136314880;
      18092: inst = 32'd268468224;
      18093: inst = 32'd201347467;
      18094: inst = 32'd203472375;
      18095: inst = 32'd136314880;
      18096: inst = 32'd268468224;
      18097: inst = 32'd201347468;
      18098: inst = 32'd203470295;
      18099: inst = 32'd136314880;
      18100: inst = 32'd268468224;
      18101: inst = 32'd201347469;
      18102: inst = 32'd203470295;
      18103: inst = 32'd136314880;
      18104: inst = 32'd268468224;
      18105: inst = 32'd201347470;
      18106: inst = 32'd203472408;
      18107: inst = 32'd136314880;
      18108: inst = 32'd268468224;
      18109: inst = 32'd201347471;
      18110: inst = 32'd203470295;
      18111: inst = 32'd136314880;
      18112: inst = 32'd268468224;
      18113: inst = 32'd201347472;
      18114: inst = 32'd203470326;
      18115: inst = 32'd136314880;
      18116: inst = 32'd268468224;
      18117: inst = 32'd201347473;
      18118: inst = 32'd203472405;
      18119: inst = 32'd136314880;
      18120: inst = 32'd268468224;
      18121: inst = 32'd201347474;
      18122: inst = 32'd203470325;
      18123: inst = 32'd136314880;
      18124: inst = 32'd268468224;
      18125: inst = 32'd201347475;
      18126: inst = 32'd203472374;
      18127: inst = 32'd136314880;
      18128: inst = 32'd268468224;
      18129: inst = 32'd201347476;
      18130: inst = 32'd203459697;
      18131: inst = 32'd136314880;
      18132: inst = 32'd268468224;
      18133: inst = 32'd201347477;
      18134: inst = 32'd203453294;
      18135: inst = 32'd136314880;
      18136: inst = 32'd268468224;
      18137: inst = 32'd201347478;
      18138: inst = 32'd203453260;
      18139: inst = 32'd136314880;
      18140: inst = 32'd268468224;
      18141: inst = 32'd201347479;
      18142: inst = 32'd203484887;
      18143: inst = 32'd136314880;
      18144: inst = 32'd268468224;
      18145: inst = 32'd201347480;
      18146: inst = 32'd203484853;
      18147: inst = 32'd136314880;
      18148: inst = 32'd268468224;
      18149: inst = 32'd201347481;
      18150: inst = 32'd203484821;
      18151: inst = 32'd136314880;
      18152: inst = 32'd268468224;
      18153: inst = 32'd201347482;
      18154: inst = 32'd203486935;
      18155: inst = 32'd136314880;
      18156: inst = 32'd268468224;
      18157: inst = 32'd201347483;
      18158: inst = 32'd203484854;
      18159: inst = 32'd136314880;
      18160: inst = 32'd268468224;
      18161: inst = 32'd201347484;
      18162: inst = 32'd203484855;
      18163: inst = 32'd136314880;
      18164: inst = 32'd268468224;
      18165: inst = 32'd201347485;
      18166: inst = 32'd203482775;
      18167: inst = 32'd136314880;
      18168: inst = 32'd268468224;
      18169: inst = 32'd201347486;
      18170: inst = 32'd203478487;
      18171: inst = 32'd136314880;
      18172: inst = 32'd268468224;
      18173: inst = 32'd201347487;
      18174: inst = 32'd203451052;
      18175: inst = 32'd136314880;
      18176: inst = 32'd268468224;
      18177: inst = 32'd201347488;
      18178: inst = 32'd203447083;
      18179: inst = 32'd136314880;
      18180: inst = 32'd268468224;
      18181: inst = 32'd201347489;
      18182: inst = 32'd203447084;
      18183: inst = 32'd136314880;
      18184: inst = 32'd268468224;
      18185: inst = 32'd201347490;
      18186: inst = 32'd203440746;
      18187: inst = 32'd136314880;
      18188: inst = 32'd268468224;
      18189: inst = 32'd201347491;
      18190: inst = 32'd203442827;
      18191: inst = 32'd136314880;
      18192: inst = 32'd268468224;
      18193: inst = 32'd201347492;
      18194: inst = 32'd203440747;
      18195: inst = 32'd136314880;
      18196: inst = 32'd268468224;
      18197: inst = 32'd201347493;
      18198: inst = 32'd203440746;
      18199: inst = 32'd136314880;
      18200: inst = 32'd268468224;
      18201: inst = 32'd201347494;
      18202: inst = 32'd203449100;
      18203: inst = 32'd136314880;
      18204: inst = 32'd268468224;
      18205: inst = 32'd201347495;
      18206: inst = 32'd203449099;
      18207: inst = 32'd136314880;
      18208: inst = 32'd268468224;
      18209: inst = 32'd201347496;
      18210: inst = 32'd203461743;
      18211: inst = 32'd136314880;
      18212: inst = 32'd268468224;
      18213: inst = 32'd201347497;
      18214: inst = 32'd203463823;
      18215: inst = 32'd136314880;
      18216: inst = 32'd268468224;
      18217: inst = 32'd201347498;
      18218: inst = 32'd203480726;
      18219: inst = 32'd136314880;
      18220: inst = 32'd268468224;
      18221: inst = 32'd201347499;
      18222: inst = 32'd203484887;
      18223: inst = 32'd136314880;
      18224: inst = 32'd268468224;
      18225: inst = 32'd201347500;
      18226: inst = 32'd203482774;
      18227: inst = 32'd136314880;
      18228: inst = 32'd268468224;
      18229: inst = 32'd201347501;
      18230: inst = 32'd203486968;
      18231: inst = 32'd136314880;
      18232: inst = 32'd268468224;
      18233: inst = 32'd201347502;
      18234: inst = 32'd203482743;
      18235: inst = 32'd136314880;
      18236: inst = 32'd268468224;
      18237: inst = 32'd201347503;
      18238: inst = 32'd203484857;
      18239: inst = 32'd136314880;
      18240: inst = 32'd268468224;
      18241: inst = 32'd201347504;
      18242: inst = 32'd203484857;
      18243: inst = 32'd136314880;
      18244: inst = 32'd268468224;
      18245: inst = 32'd201347505;
      18246: inst = 32'd203482743;
      18247: inst = 32'd136314880;
      18248: inst = 32'd268468224;
      18249: inst = 32'd201347506;
      18250: inst = 32'd203486968;
      18251: inst = 32'd136314880;
      18252: inst = 32'd268468224;
      18253: inst = 32'd201347507;
      18254: inst = 32'd203482774;
      18255: inst = 32'd136314880;
      18256: inst = 32'd268468224;
      18257: inst = 32'd201347508;
      18258: inst = 32'd203484887;
      18259: inst = 32'd136314880;
      18260: inst = 32'd268468224;
      18261: inst = 32'd201347509;
      18262: inst = 32'd203480726;
      18263: inst = 32'd136314880;
      18264: inst = 32'd268468224;
      18265: inst = 32'd201347510;
      18266: inst = 32'd203463823;
      18267: inst = 32'd136314880;
      18268: inst = 32'd268468224;
      18269: inst = 32'd201347511;
      18270: inst = 32'd203461743;
      18271: inst = 32'd136314880;
      18272: inst = 32'd268468224;
      18273: inst = 32'd201347512;
      18274: inst = 32'd203449099;
      18275: inst = 32'd136314880;
      18276: inst = 32'd268468224;
      18277: inst = 32'd201347513;
      18278: inst = 32'd203447052;
      18279: inst = 32'd136314880;
      18280: inst = 32'd268468224;
      18281: inst = 32'd201347514;
      18282: inst = 32'd203440746;
      18283: inst = 32'd136314880;
      18284: inst = 32'd268468224;
      18285: inst = 32'd201347515;
      18286: inst = 32'd203440747;
      18287: inst = 32'd136314880;
      18288: inst = 32'd268468224;
      18289: inst = 32'd201347516;
      18290: inst = 32'd203442827;
      18291: inst = 32'd136314880;
      18292: inst = 32'd268468224;
      18293: inst = 32'd201347517;
      18294: inst = 32'd203440746;
      18295: inst = 32'd136314880;
      18296: inst = 32'd268468224;
      18297: inst = 32'd201347518;
      18298: inst = 32'd203447084;
      18299: inst = 32'd136314880;
      18300: inst = 32'd268468224;
      18301: inst = 32'd201347519;
      18302: inst = 32'd203447083;
      18303: inst = 32'd136314880;
      18304: inst = 32'd268468224;
      18305: inst = 32'd201347520;
      18306: inst = 32'd203449065;
      18307: inst = 32'd136314880;
      18308: inst = 32'd268468224;
      18309: inst = 32'd201347521;
      18310: inst = 32'd203476469;
      18311: inst = 32'd136314880;
      18312: inst = 32'd268468224;
      18313: inst = 32'd201347522;
      18314: inst = 32'd203482775;
      18315: inst = 32'd136314880;
      18316: inst = 32'd268468224;
      18317: inst = 32'd201347523;
      18318: inst = 32'd203482840;
      18319: inst = 32'd136314880;
      18320: inst = 32'd268468224;
      18321: inst = 32'd201347524;
      18322: inst = 32'd203482808;
      18323: inst = 32'd136314880;
      18324: inst = 32'd268468224;
      18325: inst = 32'd201347525;
      18326: inst = 32'd203486967;
      18327: inst = 32'd136314880;
      18328: inst = 32'd268468224;
      18329: inst = 32'd201347526;
      18330: inst = 32'd203484821;
      18331: inst = 32'd136314880;
      18332: inst = 32'd268468224;
      18333: inst = 32'd201347527;
      18334: inst = 32'd203484854;
      18335: inst = 32'd136314880;
      18336: inst = 32'd268468224;
      18337: inst = 32'd201347528;
      18338: inst = 32'd203482839;
      18339: inst = 32'd136314880;
      18340: inst = 32'd268468224;
      18341: inst = 32'd201347529;
      18342: inst = 32'd203484854;
      18343: inst = 32'd136314880;
      18344: inst = 32'd268468224;
      18345: inst = 32'd201347530;
      18346: inst = 32'd203486901;
      18347: inst = 32'd136314880;
      18348: inst = 32'd268468224;
      18349: inst = 32'd201347531;
      18350: inst = 32'd203484853;
      18351: inst = 32'd136314880;
      18352: inst = 32'd268468224;
      18353: inst = 32'd201347532;
      18354: inst = 32'd203482840;
      18355: inst = 32'd136314880;
      18356: inst = 32'd268468224;
      18357: inst = 32'd201347533;
      18358: inst = 32'd203484856;
      18359: inst = 32'd136314880;
      18360: inst = 32'd268468224;
      18361: inst = 32'd201347534;
      18362: inst = 32'd203488884;
      18363: inst = 32'd136314880;
      18364: inst = 32'd268468224;
      18365: inst = 32'd201347535;
      18366: inst = 32'd203471619;
      18367: inst = 32'd136314880;
      18368: inst = 32'd268468224;
      18369: inst = 32'd201347536;
      18370: inst = 32'd203480005;
      18371: inst = 32'd136314880;
      18372: inst = 32'd268468224;
      18373: inst = 32'd201347537;
      18374: inst = 32'd203480005;
      18375: inst = 32'd136314880;
      18376: inst = 32'd268468224;
      18377: inst = 32'd201347538;
      18378: inst = 32'd203480005;
      18379: inst = 32'd136314880;
      18380: inst = 32'd268468224;
      18381: inst = 32'd201347539;
      18382: inst = 32'd203480005;
      18383: inst = 32'd136314880;
      18384: inst = 32'd268468224;
      18385: inst = 32'd201347540;
      18386: inst = 32'd203480005;
      18387: inst = 32'd136314880;
      18388: inst = 32'd268468224;
      18389: inst = 32'd201347541;
      18390: inst = 32'd203480005;
      18391: inst = 32'd136314880;
      18392: inst = 32'd268468224;
      18393: inst = 32'd201347542;
      18394: inst = 32'd203480005;
      18395: inst = 32'd136314880;
      18396: inst = 32'd268468224;
      18397: inst = 32'd201347543;
      18398: inst = 32'd203480005;
      18399: inst = 32'd136314880;
      18400: inst = 32'd268468224;
      18401: inst = 32'd201347544;
      18402: inst = 32'd203480005;
      18403: inst = 32'd136314880;
      18404: inst = 32'd268468224;
      18405: inst = 32'd201347545;
      18406: inst = 32'd203480005;
      18407: inst = 32'd136314880;
      18408: inst = 32'd268468224;
      18409: inst = 32'd201347546;
      18410: inst = 32'd203479973;
      18411: inst = 32'd136314880;
      18412: inst = 32'd268468224;
      18413: inst = 32'd201347547;
      18414: inst = 32'd203480005;
      18415: inst = 32'd136314880;
      18416: inst = 32'd268468224;
      18417: inst = 32'd201347548;
      18418: inst = 32'd203479973;
      18419: inst = 32'd136314880;
      18420: inst = 32'd268468224;
      18421: inst = 32'd201347549;
      18422: inst = 32'd203480005;
      18423: inst = 32'd136314880;
      18424: inst = 32'd268468224;
      18425: inst = 32'd201347550;
      18426: inst = 32'd203479973;
      18427: inst = 32'd136314880;
      18428: inst = 32'd268468224;
      18429: inst = 32'd201347551;
      18430: inst = 32'd203473634;
      18431: inst = 32'd136314880;
      18432: inst = 32'd268468224;
      18433: inst = 32'd201347552;
      18434: inst = 32'd203459665;
      18435: inst = 32'd136314880;
      18436: inst = 32'd268468224;
      18437: inst = 32'd201347553;
      18438: inst = 32'd203472375;
      18439: inst = 32'd136314880;
      18440: inst = 32'd268468224;
      18441: inst = 32'd201347554;
      18442: inst = 32'd203472375;
      18443: inst = 32'd136314880;
      18444: inst = 32'd268468224;
      18445: inst = 32'd201347555;
      18446: inst = 32'd203470295;
      18447: inst = 32'd136314880;
      18448: inst = 32'd268468224;
      18449: inst = 32'd201347556;
      18450: inst = 32'd203472408;
      18451: inst = 32'd136314880;
      18452: inst = 32'd268468224;
      18453: inst = 32'd201347557;
      18454: inst = 32'd203472343;
      18455: inst = 32'd136314880;
      18456: inst = 32'd268468224;
      18457: inst = 32'd201347558;
      18458: inst = 32'd203472343;
      18459: inst = 32'd136314880;
      18460: inst = 32'd268468224;
      18461: inst = 32'd201347559;
      18462: inst = 32'd203472375;
      18463: inst = 32'd136314880;
      18464: inst = 32'd268468224;
      18465: inst = 32'd201347560;
      18466: inst = 32'd203472375;
      18467: inst = 32'd136314880;
      18468: inst = 32'd268468224;
      18469: inst = 32'd201347561;
      18470: inst = 32'd203470295;
      18471: inst = 32'd136314880;
      18472: inst = 32'd268468224;
      18473: inst = 32'd201347562;
      18474: inst = 32'd203459697;
      18475: inst = 32'd136314880;
      18476: inst = 32'd268468224;
      18477: inst = 32'd201347563;
      18478: inst = 32'd203472375;
      18479: inst = 32'd136314880;
      18480: inst = 32'd268468224;
      18481: inst = 32'd201347564;
      18482: inst = 32'd203472343;
      18483: inst = 32'd136314880;
      18484: inst = 32'd268468224;
      18485: inst = 32'd201347565;
      18486: inst = 32'd203472375;
      18487: inst = 32'd136314880;
      18488: inst = 32'd268468224;
      18489: inst = 32'd201347566;
      18490: inst = 32'd203472375;
      18491: inst = 32'd136314880;
      18492: inst = 32'd268468224;
      18493: inst = 32'd201347567;
      18494: inst = 32'd203472343;
      18495: inst = 32'd136314880;
      18496: inst = 32'd268468224;
      18497: inst = 32'd201347568;
      18498: inst = 32'd203470293;
      18499: inst = 32'd136314880;
      18500: inst = 32'd268468224;
      18501: inst = 32'd201347569;
      18502: inst = 32'd203472439;
      18503: inst = 32'd136314880;
      18504: inst = 32'd268468224;
      18505: inst = 32'd201347570;
      18506: inst = 32'd203472342;
      18507: inst = 32'd136314880;
      18508: inst = 32'd268468224;
      18509: inst = 32'd201347571;
      18510: inst = 32'd203472343;
      18511: inst = 32'd136314880;
      18512: inst = 32'd268468224;
      18513: inst = 32'd201347572;
      18514: inst = 32'd203461713;
      18515: inst = 32'd136314880;
      18516: inst = 32'd268468224;
      18517: inst = 32'd201347573;
      18518: inst = 32'd203455341;
      18519: inst = 32'd136314880;
      18520: inst = 32'd268468224;
      18521: inst = 32'd201347574;
      18522: inst = 32'd203455308;
      18523: inst = 32'd136314880;
      18524: inst = 32'd268468224;
      18525: inst = 32'd201347575;
      18526: inst = 32'd203484856;
      18527: inst = 32'd136314880;
      18528: inst = 32'd268468224;
      18529: inst = 32'd201347576;
      18530: inst = 32'd203486936;
      18531: inst = 32'd136314880;
      18532: inst = 32'd268468224;
      18533: inst = 32'd201347577;
      18534: inst = 32'd203482774;
      18535: inst = 32'd136314880;
      18536: inst = 32'd268468224;
      18537: inst = 32'd201347578;
      18538: inst = 32'd203484886;
      18539: inst = 32'd136314880;
      18540: inst = 32'd268468224;
      18541: inst = 32'd201347579;
      18542: inst = 32'd203482807;
      18543: inst = 32'd136314880;
      18544: inst = 32'd268468224;
      18545: inst = 32'd201347580;
      18546: inst = 32'd203482840;
      18547: inst = 32'd136314880;
      18548: inst = 32'd268468224;
      18549: inst = 32'd201347581;
      18550: inst = 32'd203478648;
      18551: inst = 32'd136314880;
      18552: inst = 32'd268468224;
      18553: inst = 32'd201347582;
      18554: inst = 32'd203459632;
      18555: inst = 32'd136314880;
      18556: inst = 32'd268468224;
      18557: inst = 32'd201347583;
      18558: inst = 32'd203451180;
      18559: inst = 32'd136314880;
      18560: inst = 32'd268468224;
      18561: inst = 32'd201347584;
      18562: inst = 32'd203449132;
      18563: inst = 32'd136314880;
      18564: inst = 32'd268468224;
      18565: inst = 32'd201347585;
      18566: inst = 32'd203444971;
      18567: inst = 32'd136314880;
      18568: inst = 32'd268468224;
      18569: inst = 32'd201347586;
      18570: inst = 32'd203442793;
      18571: inst = 32'd136314880;
      18572: inst = 32'd268468224;
      18573: inst = 32'd201347587;
      18574: inst = 32'd203442826;
      18575: inst = 32'd136314880;
      18576: inst = 32'd268468224;
      18577: inst = 32'd201347588;
      18578: inst = 32'd203442794;
      18579: inst = 32'd136314880;
      18580: inst = 32'd268468224;
      18581: inst = 32'd201347589;
      18582: inst = 32'd203444906;
      18583: inst = 32'd136314880;
      18584: inst = 32'd268468224;
      18585: inst = 32'd201347590;
      18586: inst = 32'd203449067;
      18587: inst = 32'd136314880;
      18588: inst = 32'd268468224;
      18589: inst = 32'd201347591;
      18590: inst = 32'd203449035;
      18591: inst = 32'd136314880;
      18592: inst = 32'd268468224;
      18593: inst = 32'd201347592;
      18594: inst = 32'd203461745;
      18595: inst = 32'd136314880;
      18596: inst = 32'd268468224;
      18597: inst = 32'd201347593;
      18598: inst = 32'd203461647;
      18599: inst = 32'd136314880;
      18600: inst = 32'd268468224;
      18601: inst = 32'd201347594;
      18602: inst = 32'd203484889;
      18603: inst = 32'd136314880;
      18604: inst = 32'd268468224;
      18605: inst = 32'd201347595;
      18606: inst = 32'd203484791;
      18607: inst = 32'd136314880;
      18608: inst = 32'd268468224;
      18609: inst = 32'd201347596;
      18610: inst = 32'd203486903;
      18611: inst = 32'd136314880;
      18612: inst = 32'd268468224;
      18613: inst = 32'd201347597;
      18614: inst = 32'd203486902;
      18615: inst = 32'd136314880;
      18616: inst = 32'd268468224;
      18617: inst = 32'd201347598;
      18618: inst = 32'd203486870;
      18619: inst = 32'd136314880;
      18620: inst = 32'd268468224;
      18621: inst = 32'd201347599;
      18622: inst = 32'd203486869;
      18623: inst = 32'd136314880;
      18624: inst = 32'd268468224;
      18625: inst = 32'd201347600;
      18626: inst = 32'd203486869;
      18627: inst = 32'd136314880;
      18628: inst = 32'd268468224;
      18629: inst = 32'd201347601;
      18630: inst = 32'd203486870;
      18631: inst = 32'd136314880;
      18632: inst = 32'd268468224;
      18633: inst = 32'd201347602;
      18634: inst = 32'd203486902;
      18635: inst = 32'd136314880;
      18636: inst = 32'd268468224;
      18637: inst = 32'd201347603;
      18638: inst = 32'd203486903;
      18639: inst = 32'd136314880;
      18640: inst = 32'd268468224;
      18641: inst = 32'd201347604;
      18642: inst = 32'd203484823;
      18643: inst = 32'd136314880;
      18644: inst = 32'd268468224;
      18645: inst = 32'd201347605;
      18646: inst = 32'd203484889;
      18647: inst = 32'd136314880;
      18648: inst = 32'd268468224;
      18649: inst = 32'd201347606;
      18650: inst = 32'd203461679;
      18651: inst = 32'd136314880;
      18652: inst = 32'd268468224;
      18653: inst = 32'd201347607;
      18654: inst = 32'd203463793;
      18655: inst = 32'd136314880;
      18656: inst = 32'd268468224;
      18657: inst = 32'd201347608;
      18658: inst = 32'd203449035;
      18659: inst = 32'd136314880;
      18660: inst = 32'd268468224;
      18661: inst = 32'd201347609;
      18662: inst = 32'd203449067;
      18663: inst = 32'd136314880;
      18664: inst = 32'd268468224;
      18665: inst = 32'd201347610;
      18666: inst = 32'd203444906;
      18667: inst = 32'd136314880;
      18668: inst = 32'd268468224;
      18669: inst = 32'd201347611;
      18670: inst = 32'd203442794;
      18671: inst = 32'd136314880;
      18672: inst = 32'd268468224;
      18673: inst = 32'd201347612;
      18674: inst = 32'd203442826;
      18675: inst = 32'd136314880;
      18676: inst = 32'd268468224;
      18677: inst = 32'd201347613;
      18678: inst = 32'd203442793;
      18679: inst = 32'd136314880;
      18680: inst = 32'd268468224;
      18681: inst = 32'd201347614;
      18682: inst = 32'd203444971;
      18683: inst = 32'd136314880;
      18684: inst = 32'd268468224;
      18685: inst = 32'd201347615;
      18686: inst = 32'd203449132;
      18687: inst = 32'd136314880;
      18688: inst = 32'd268468224;
      18689: inst = 32'd201347616;
      18690: inst = 32'd203449131;
      18691: inst = 32'd136314880;
      18692: inst = 32'd268468224;
      18693: inst = 32'd201347617;
      18694: inst = 32'd203459695;
      18695: inst = 32'd136314880;
      18696: inst = 32'd268468224;
      18697: inst = 32'd201347618;
      18698: inst = 32'd203478614;
      18699: inst = 32'd136314880;
      18700: inst = 32'd268468224;
      18701: inst = 32'd201347619;
      18702: inst = 32'd203484919;
      18703: inst = 32'd136314880;
      18704: inst = 32'd268468224;
      18705: inst = 32'd201347620;
      18706: inst = 32'd203484854;
      18707: inst = 32'd136314880;
      18708: inst = 32'd268468224;
      18709: inst = 32'd201347621;
      18710: inst = 32'd203484821;
      18711: inst = 32'd136314880;
      18712: inst = 32'd268468224;
      18713: inst = 32'd201347622;
      18714: inst = 32'd203484853;
      18715: inst = 32'd136314880;
      18716: inst = 32'd268468224;
      18717: inst = 32'd201347623;
      18718: inst = 32'd203486934;
      18719: inst = 32'd136314880;
      18720: inst = 32'd268468224;
      18721: inst = 32'd201347624;
      18722: inst = 32'd203484854;
      18723: inst = 32'd136314880;
      18724: inst = 32'd268468224;
      18725: inst = 32'd201347625;
      18726: inst = 32'd203484886;
      18727: inst = 32'd136314880;
      18728: inst = 32'd268468224;
      18729: inst = 32'd201347626;
      18730: inst = 32'd203484854;
      18731: inst = 32'd136314880;
      18732: inst = 32'd268468224;
      18733: inst = 32'd201347627;
      18734: inst = 32'd203486901;
      18735: inst = 32'd136314880;
      18736: inst = 32'd268468224;
      18737: inst = 32'd201347628;
      18738: inst = 32'd203488916;
      18739: inst = 32'd136314880;
      18740: inst = 32'd268468224;
      18741: inst = 32'd201347629;
      18742: inst = 32'd203488850;
      18743: inst = 32'd136314880;
      18744: inst = 32'd268468224;
      18745: inst = 32'd201347630;
      18746: inst = 32'd203488946;
      18747: inst = 32'd136314880;
      18748: inst = 32'd268468224;
      18749: inst = 32'd201347631;
      18750: inst = 32'd203465508;
      18751: inst = 32'd136314880;
      18752: inst = 32'd268468224;
      18753: inst = 32'd201347632;
      18754: inst = 32'd203482021;
      18755: inst = 32'd136314880;
      18756: inst = 32'd268468224;
      18757: inst = 32'd201347633;
      18758: inst = 32'd203482021;
      18759: inst = 32'd136314880;
      18760: inst = 32'd268468224;
      18761: inst = 32'd201347634;
      18762: inst = 32'd203482021;
      18763: inst = 32'd136314880;
      18764: inst = 32'd268468224;
      18765: inst = 32'd201347635;
      18766: inst = 32'd203482021;
      18767: inst = 32'd136314880;
      18768: inst = 32'd268468224;
      18769: inst = 32'd201347636;
      18770: inst = 32'd203482021;
      18771: inst = 32'd136314880;
      18772: inst = 32'd268468224;
      18773: inst = 32'd201347637;
      18774: inst = 32'd203482021;
      18775: inst = 32'd136314880;
      18776: inst = 32'd268468224;
      18777: inst = 32'd201347638;
      18778: inst = 32'd203482021;
      18779: inst = 32'd136314880;
      18780: inst = 32'd268468224;
      18781: inst = 32'd201347639;
      18782: inst = 32'd203482021;
      18783: inst = 32'd136314880;
      18784: inst = 32'd268468224;
      18785: inst = 32'd201347640;
      18786: inst = 32'd203482021;
      18787: inst = 32'd136314880;
      18788: inst = 32'd268468224;
      18789: inst = 32'd201347641;
      18790: inst = 32'd203482021;
      18791: inst = 32'd136314880;
      18792: inst = 32'd268468224;
      18793: inst = 32'd201347642;
      18794: inst = 32'd203482053;
      18795: inst = 32'd136314880;
      18796: inst = 32'd268468224;
      18797: inst = 32'd201347643;
      18798: inst = 32'd203482021;
      18799: inst = 32'd136314880;
      18800: inst = 32'd268468224;
      18801: inst = 32'd201347644;
      18802: inst = 32'd203482021;
      18803: inst = 32'd136314880;
      18804: inst = 32'd268468224;
      18805: inst = 32'd201347645;
      18806: inst = 32'd203484101;
      18807: inst = 32'd136314880;
      18808: inst = 32'd268468224;
      18809: inst = 32'd201347646;
      18810: inst = 32'd203479940;
      18811: inst = 32'd136314880;
      18812: inst = 32'd268468224;
      18813: inst = 32'd201347647;
      18814: inst = 32'd203475682;
      18815: inst = 32'd136314880;
      18816: inst = 32'd268468224;
      18817: inst = 32'd201347648;
      18818: inst = 32'd203461811;
      18819: inst = 32'd136314880;
      18820: inst = 32'd268468224;
      18821: inst = 32'd201347649;
      18822: inst = 32'd203470295;
      18823: inst = 32'd136314880;
      18824: inst = 32'd268468224;
      18825: inst = 32'd201347650;
      18826: inst = 32'd203470295;
      18827: inst = 32'd136314880;
      18828: inst = 32'd268468224;
      18829: inst = 32'd201347651;
      18830: inst = 32'd203470263;
      18831: inst = 32'd136314880;
      18832: inst = 32'd268468224;
      18833: inst = 32'd201347652;
      18834: inst = 32'd203472376;
      18835: inst = 32'd136314880;
      18836: inst = 32'd268468224;
      18837: inst = 32'd201347653;
      18838: inst = 32'd203472343;
      18839: inst = 32'd136314880;
      18840: inst = 32'd268468224;
      18841: inst = 32'd201347654;
      18842: inst = 32'd203472343;
      18843: inst = 32'd136314880;
      18844: inst = 32'd268468224;
      18845: inst = 32'd201347655;
      18846: inst = 32'd203472343;
      18847: inst = 32'd136314880;
      18848: inst = 32'd268468224;
      18849: inst = 32'd201347656;
      18850: inst = 32'd203472343;
      18851: inst = 32'd136314880;
      18852: inst = 32'd268468224;
      18853: inst = 32'd201347657;
      18854: inst = 32'd203470263;
      18855: inst = 32'd136314880;
      18856: inst = 32'd268468224;
      18857: inst = 32'd201347658;
      18858: inst = 32'd203463891;
      18859: inst = 32'd136314880;
      18860: inst = 32'd268468224;
      18861: inst = 32'd201347659;
      18862: inst = 32'd203472343;
      18863: inst = 32'd136314880;
      18864: inst = 32'd268468224;
      18865: inst = 32'd201347660;
      18866: inst = 32'd203470263;
      18867: inst = 32'd136314880;
      18868: inst = 32'd268468224;
      18869: inst = 32'd201347661;
      18870: inst = 32'd203472343;
      18871: inst = 32'd136314880;
      18872: inst = 32'd268468224;
      18873: inst = 32'd201347662;
      18874: inst = 32'd203472343;
      18875: inst = 32'd136314880;
      18876: inst = 32'd268468224;
      18877: inst = 32'd201347663;
      18878: inst = 32'd203472343;
      18879: inst = 32'd136314880;
      18880: inst = 32'd268468224;
      18881: inst = 32'd201347664;
      18882: inst = 32'd203470326;
      18883: inst = 32'd136314880;
      18884: inst = 32'd268468224;
      18885: inst = 32'd201347665;
      18886: inst = 32'd203472407;
      18887: inst = 32'd136314880;
      18888: inst = 32'd268468224;
      18889: inst = 32'd201347666;
      18890: inst = 32'd203472375;
      18891: inst = 32'd136314880;
      18892: inst = 32'd268468224;
      18893: inst = 32'd201347667;
      18894: inst = 32'd203472375;
      18895: inst = 32'd136314880;
      18896: inst = 32'd268468224;
      18897: inst = 32'd201347668;
      18898: inst = 32'd203461714;
      18899: inst = 32'd136314880;
      18900: inst = 32'd268468224;
      18901: inst = 32'd201347669;
      18902: inst = 32'd203453196;
      18903: inst = 32'd136314880;
      18904: inst = 32'd268468224;
      18905: inst = 32'd201347670;
      18906: inst = 32'd203455276;
      18907: inst = 32'd136314880;
      18908: inst = 32'd268468224;
      18909: inst = 32'd201347671;
      18910: inst = 32'd203484889;
      18911: inst = 32'd136314880;
      18912: inst = 32'd268468224;
      18913: inst = 32'd201347672;
      18914: inst = 32'd203482775;
      18915: inst = 32'd136314880;
      18916: inst = 32'd268468224;
      18917: inst = 32'd201347673;
      18918: inst = 32'd203484887;
      18919: inst = 32'd136314880;
      18920: inst = 32'd268468224;
      18921: inst = 32'd201347674;
      18922: inst = 32'd203484952;
      18923: inst = 32'd136314880;
      18924: inst = 32'd268468224;
      18925: inst = 32'd201347675;
      18926: inst = 32'd203480727;
      18927: inst = 32'd136314880;
      18928: inst = 32'd268468224;
      18929: inst = 32'd201347676;
      18930: inst = 32'd203480727;
      18931: inst = 32'd136314880;
      18932: inst = 32'd268468224;
      18933: inst = 32'd201347677;
      18934: inst = 32'd203463857;
      18935: inst = 32'd136314880;
      18936: inst = 32'd268468224;
      18937: inst = 32'd201347678;
      18938: inst = 32'd203461778;
      18939: inst = 32'd136314880;
      18940: inst = 32'd268468224;
      18941: inst = 32'd201347679;
      18942: inst = 32'd203449068;
      18943: inst = 32'd136314880;
      18944: inst = 32'd268468224;
      18945: inst = 32'd201347680;
      18946: inst = 32'd203447019;
      18947: inst = 32'd136314880;
      18948: inst = 32'd268468224;
      18949: inst = 32'd201347681;
      18950: inst = 32'd203444939;
      18951: inst = 32'd136314880;
      18952: inst = 32'd268468224;
      18953: inst = 32'd201347682;
      18954: inst = 32'd203442794;
      18955: inst = 32'd136314880;
      18956: inst = 32'd268468224;
      18957: inst = 32'd201347683;
      18958: inst = 32'd203442794;
      18959: inst = 32'd136314880;
      18960: inst = 32'd268468224;
      18961: inst = 32'd201347684;
      18962: inst = 32'd203440713;
      18963: inst = 32'd136314880;
      18964: inst = 32'd268468224;
      18965: inst = 32'd201347685;
      18966: inst = 32'd203442793;
      18967: inst = 32'd136314880;
      18968: inst = 32'd268468224;
      18969: inst = 32'd201347686;
      18970: inst = 32'd203449067;
      18971: inst = 32'd136314880;
      18972: inst = 32'd268468224;
      18973: inst = 32'd201347687;
      18974: inst = 32'd203451180;
      18975: inst = 32'd136314880;
      18976: inst = 32'd268468224;
      18977: inst = 32'd201347688;
      18978: inst = 32'd203461745;
      18979: inst = 32'd136314880;
      18980: inst = 32'd268468224;
      18981: inst = 32'd201347689;
      18982: inst = 32'd203461679;
      18983: inst = 32'd136314880;
      18984: inst = 32'd268468224;
      18985: inst = 32'd201347690;
      18986: inst = 32'd203484889;
      18987: inst = 32'd136314880;
      18988: inst = 32'd268468224;
      18989: inst = 32'd201347691;
      18990: inst = 32'd203484856;
      18991: inst = 32'd136314880;
      18992: inst = 32'd268468224;
      18993: inst = 32'd201347692;
      18994: inst = 32'd203484856;
      18995: inst = 32'd136314880;
      18996: inst = 32'd268468224;
      18997: inst = 32'd201347693;
      18998: inst = 32'd203484823;
      18999: inst = 32'd136314880;
      19000: inst = 32'd268468224;
      19001: inst = 32'd201347694;
      19002: inst = 32'd203484854;
      19003: inst = 32'd136314880;
      19004: inst = 32'd268468224;
      19005: inst = 32'd201347695;
      19006: inst = 32'd203486935;
      19007: inst = 32'd136314880;
      19008: inst = 32'd268468224;
      19009: inst = 32'd201347696;
      19010: inst = 32'd203486903;
      19011: inst = 32'd136314880;
      19012: inst = 32'd268468224;
      19013: inst = 32'd201347697;
      19014: inst = 32'd203484822;
      19015: inst = 32'd136314880;
      19016: inst = 32'd268468224;
      19017: inst = 32'd201347698;
      19018: inst = 32'd203484823;
      19019: inst = 32'd136314880;
      19020: inst = 32'd268468224;
      19021: inst = 32'd201347699;
      19022: inst = 32'd203484855;
      19023: inst = 32'd136314880;
      19024: inst = 32'd268468224;
      19025: inst = 32'd201347700;
      19026: inst = 32'd203482776;
      19027: inst = 32'd136314880;
      19028: inst = 32'd268468224;
      19029: inst = 32'd201347701;
      19030: inst = 32'd203484889;
      19031: inst = 32'd136314880;
      19032: inst = 32'd268468224;
      19033: inst = 32'd201347702;
      19034: inst = 32'd203461679;
      19035: inst = 32'd136314880;
      19036: inst = 32'd268468224;
      19037: inst = 32'd201347703;
      19038: inst = 32'd203461713;
      19039: inst = 32'd136314880;
      19040: inst = 32'd268468224;
      19041: inst = 32'd201347704;
      19042: inst = 32'd203451180;
      19043: inst = 32'd136314880;
      19044: inst = 32'd268468224;
      19045: inst = 32'd201347705;
      19046: inst = 32'd203449067;
      19047: inst = 32'd136314880;
      19048: inst = 32'd268468224;
      19049: inst = 32'd201347706;
      19050: inst = 32'd203442793;
      19051: inst = 32'd136314880;
      19052: inst = 32'd268468224;
      19053: inst = 32'd201347707;
      19054: inst = 32'd203440713;
      19055: inst = 32'd136314880;
      19056: inst = 32'd268468224;
      19057: inst = 32'd201347708;
      19058: inst = 32'd203442794;
      19059: inst = 32'd136314880;
      19060: inst = 32'd268468224;
      19061: inst = 32'd201347709;
      19062: inst = 32'd203442794;
      19063: inst = 32'd136314880;
      19064: inst = 32'd268468224;
      19065: inst = 32'd201347710;
      19066: inst = 32'd203444939;
      19067: inst = 32'd136314880;
      19068: inst = 32'd268468224;
      19069: inst = 32'd201347711;
      19070: inst = 32'd203447019;
      19071: inst = 32'd136314880;
      19072: inst = 32'd268468224;
      19073: inst = 32'd201347712;
      19074: inst = 32'd203447019;
      19075: inst = 32'd136314880;
      19076: inst = 32'd268468224;
      19077: inst = 32'd201347713;
      19078: inst = 32'd203463857;
      19079: inst = 32'd136314880;
      19080: inst = 32'd268468224;
      19081: inst = 32'd201347714;
      19082: inst = 32'd203463856;
      19083: inst = 32'd136314880;
      19084: inst = 32'd268468224;
      19085: inst = 32'd201347715;
      19086: inst = 32'd203480695;
      19087: inst = 32'd136314880;
      19088: inst = 32'd268468224;
      19089: inst = 32'd201347716;
      19090: inst = 32'd203482775;
      19091: inst = 32'd136314880;
      19092: inst = 32'd268468224;
      19093: inst = 32'd201347717;
      19094: inst = 32'd203486935;
      19095: inst = 32'd136314880;
      19096: inst = 32'd268468224;
      19097: inst = 32'd201347718;
      19098: inst = 32'd203486967;
      19099: inst = 32'd136314880;
      19100: inst = 32'd268468224;
      19101: inst = 32'd201347719;
      19102: inst = 32'd203482774;
      19103: inst = 32'd136314880;
      19104: inst = 32'd268468224;
      19105: inst = 32'd201347720;
      19106: inst = 32'd203482807;
      19107: inst = 32'd136314880;
      19108: inst = 32'd268468224;
      19109: inst = 32'd201347721;
      19110: inst = 32'd203484887;
      19111: inst = 32'd136314880;
      19112: inst = 32'd268468224;
      19113: inst = 32'd201347722;
      19114: inst = 32'd203484888;
      19115: inst = 32'd136314880;
      19116: inst = 32'd268468224;
      19117: inst = 32'd201347723;
      19118: inst = 32'd203484854;
      19119: inst = 32'd136314880;
      19120: inst = 32'd268468224;
      19121: inst = 32'd201347724;
      19122: inst = 32'd203488950;
      19123: inst = 32'd136314880;
      19124: inst = 32'd268468224;
      19125: inst = 32'd201347725;
      19126: inst = 32'd203488949;
      19127: inst = 32'd136314880;
      19128: inst = 32'd268468224;
      19129: inst = 32'd201347726;
      19130: inst = 32'd203488884;
      19131: inst = 32'd136314880;
      19132: inst = 32'd268468224;
      19133: inst = 32'd201347727;
      19134: inst = 32'd203463429;
      19135: inst = 32'd136314880;
      19136: inst = 32'd268468224;
      19137: inst = 32'd201347728;
      19138: inst = 32'd203479973;
      19139: inst = 32'd136314880;
      19140: inst = 32'd268468224;
      19141: inst = 32'd201347729;
      19142: inst = 32'd203479973;
      19143: inst = 32'd136314880;
      19144: inst = 32'd268468224;
      19145: inst = 32'd201347730;
      19146: inst = 32'd203479973;
      19147: inst = 32'd136314880;
      19148: inst = 32'd268468224;
      19149: inst = 32'd201347731;
      19150: inst = 32'd203479973;
      19151: inst = 32'd136314880;
      19152: inst = 32'd268468224;
      19153: inst = 32'd201347732;
      19154: inst = 32'd203479973;
      19155: inst = 32'd136314880;
      19156: inst = 32'd268468224;
      19157: inst = 32'd201347733;
      19158: inst = 32'd203479973;
      19159: inst = 32'd136314880;
      19160: inst = 32'd268468224;
      19161: inst = 32'd201347734;
      19162: inst = 32'd203479973;
      19163: inst = 32'd136314880;
      19164: inst = 32'd268468224;
      19165: inst = 32'd201347735;
      19166: inst = 32'd203479973;
      19167: inst = 32'd136314880;
      19168: inst = 32'd268468224;
      19169: inst = 32'd201347736;
      19170: inst = 32'd203479973;
      19171: inst = 32'd136314880;
      19172: inst = 32'd268468224;
      19173: inst = 32'd201347737;
      19174: inst = 32'd203479973;
      19175: inst = 32'd136314880;
      19176: inst = 32'd268468224;
      19177: inst = 32'd201347738;
      19178: inst = 32'd203479973;
      19179: inst = 32'd136314880;
      19180: inst = 32'd268468224;
      19181: inst = 32'd201347739;
      19182: inst = 32'd203479973;
      19183: inst = 32'd136314880;
      19184: inst = 32'd268468224;
      19185: inst = 32'd201347740;
      19186: inst = 32'd203479973;
      19187: inst = 32'd136314880;
      19188: inst = 32'd268468224;
      19189: inst = 32'd201347741;
      19190: inst = 32'd203482053;
      19191: inst = 32'd136314880;
      19192: inst = 32'd268468224;
      19193: inst = 32'd201347742;
      19194: inst = 32'd203479941;
      19195: inst = 32'd136314880;
      19196: inst = 32'd268468224;
      19197: inst = 32'd201347743;
      19198: inst = 32'd203475747;
      19199: inst = 32'd136314880;
      19200: inst = 32'd268468224;
      19201: inst = 32'd201347744;
      19202: inst = 32'd203457553;
      19203: inst = 32'd136314880;
      19204: inst = 32'd268468224;
      19205: inst = 32'd201347745;
      19206: inst = 32'd203461779;
      19207: inst = 32'd136314880;
      19208: inst = 32'd268468224;
      19209: inst = 32'd201347746;
      19210: inst = 32'd203459698;
      19211: inst = 32'd136314880;
      19212: inst = 32'd268468224;
      19213: inst = 32'd201347747;
      19214: inst = 32'd203459666;
      19215: inst = 32'd136314880;
      19216: inst = 32'd268468224;
      19217: inst = 32'd201347748;
      19218: inst = 32'd203459698;
      19219: inst = 32'd136314880;
      19220: inst = 32'd268468224;
      19221: inst = 32'd201347749;
      19222: inst = 32'd203459698;
      19223: inst = 32'd136314880;
      19224: inst = 32'd268468224;
      19225: inst = 32'd201347750;
      19226: inst = 32'd203459698;
      19227: inst = 32'd136314880;
      19228: inst = 32'd268468224;
      19229: inst = 32'd201347751;
      19230: inst = 32'd203459666;
      19231: inst = 32'd136314880;
      19232: inst = 32'd268468224;
      19233: inst = 32'd201347752;
      19234: inst = 32'd203459698;
      19235: inst = 32'd136314880;
      19236: inst = 32'd268468224;
      19237: inst = 32'd201347753;
      19238: inst = 32'd203459698;
      19239: inst = 32'd136314880;
      19240: inst = 32'd268468224;
      19241: inst = 32'd201347754;
      19242: inst = 32'd203457553;
      19243: inst = 32'd136314880;
      19244: inst = 32'd268468224;
      19245: inst = 32'd201347755;
      19246: inst = 32'd203459698;
      19247: inst = 32'd136314880;
      19248: inst = 32'd268468224;
      19249: inst = 32'd201347756;
      19250: inst = 32'd203459698;
      19251: inst = 32'd136314880;
      19252: inst = 32'd268468224;
      19253: inst = 32'd201347757;
      19254: inst = 32'd203459698;
      19255: inst = 32'd136314880;
      19256: inst = 32'd268468224;
      19257: inst = 32'd201347758;
      19258: inst = 32'd203459698;
      19259: inst = 32'd136314880;
      19260: inst = 32'd268468224;
      19261: inst = 32'd201347759;
      19262: inst = 32'd203459698;
      19263: inst = 32'd136314880;
      19264: inst = 32'd268468224;
      19265: inst = 32'd201347760;
      19266: inst = 32'd203457681;
      19267: inst = 32'd136314880;
      19268: inst = 32'd268468224;
      19269: inst = 32'd201347761;
      19270: inst = 32'd203457649;
      19271: inst = 32'd136314880;
      19272: inst = 32'd268468224;
      19273: inst = 32'd201347762;
      19274: inst = 32'd203459666;
      19275: inst = 32'd136314880;
      19276: inst = 32'd268468224;
      19277: inst = 32'd201347763;
      19278: inst = 32'd203461812;
      19279: inst = 32'd136314880;
      19280: inst = 32'd268468224;
      19281: inst = 32'd201347764;
      19282: inst = 32'd203459666;
      19283: inst = 32'd136314880;
      19284: inst = 32'd268468224;
      19285: inst = 32'd201347765;
      19286: inst = 32'd203455375;
      19287: inst = 32'd136314880;
      19288: inst = 32'd268468224;
      19289: inst = 32'd201347766;
      19290: inst = 32'd203457455;
      19291: inst = 32'd136314880;
      19292: inst = 32'd268468224;
      19293: inst = 32'd201347767;
      19294: inst = 32'd203480664;
      19295: inst = 32'd136314880;
      19296: inst = 32'd268468224;
      19297: inst = 32'd201347768;
      19298: inst = 32'd203480728;
      19299: inst = 32'd136314880;
      19300: inst = 32'd268468224;
      19301: inst = 32'd201347769;
      19302: inst = 32'd203484921;
      19303: inst = 32'd136314880;
      19304: inst = 32'd268468224;
      19305: inst = 32'd201347770;
      19306: inst = 32'd203480727;
      19307: inst = 32'd136314880;
      19308: inst = 32'd268468224;
      19309: inst = 32'd201347771;
      19310: inst = 32'd203482840;
      19311: inst = 32'd136314880;
      19312: inst = 32'd268468224;
      19313: inst = 32'd201347772;
      19314: inst = 32'd203472276;
      19315: inst = 32'd136314880;
      19316: inst = 32'd268468224;
      19317: inst = 32'd201347773;
      19318: inst = 32'd203459632;
      19319: inst = 32'd136314880;
      19320: inst = 32'd268468224;
      19321: inst = 32'd201347774;
      19322: inst = 32'd203459665;
      19323: inst = 32'd136314880;
      19324: inst = 32'd268468224;
      19325: inst = 32'd201347775;
      19326: inst = 32'd203446988;
      19327: inst = 32'd136314880;
      19328: inst = 32'd268468224;
      19329: inst = 32'd201347776;
      19330: inst = 32'd203449100;
      19331: inst = 32'd136314880;
      19332: inst = 32'd268468224;
      19333: inst = 32'd201347777;
      19334: inst = 32'd203447019;
      19335: inst = 32'd136314880;
      19336: inst = 32'd268468224;
      19337: inst = 32'd201347778;
      19338: inst = 32'd203442794;
      19339: inst = 32'd136314880;
      19340: inst = 32'd268468224;
      19341: inst = 32'd201347779;
      19342: inst = 32'd203442794;
      19343: inst = 32'd136314880;
      19344: inst = 32'd268468224;
      19345: inst = 32'd201347780;
      19346: inst = 32'd203444874;
      19347: inst = 32'd136314880;
      19348: inst = 32'd268468224;
      19349: inst = 32'd201347781;
      19350: inst = 32'd203444906;
      19351: inst = 32'd136314880;
      19352: inst = 32'd268468224;
      19353: inst = 32'd201347782;
      19354: inst = 32'd203447020;
      19355: inst = 32'd136314880;
      19356: inst = 32'd268468224;
      19357: inst = 32'd201347783;
      19358: inst = 32'd203446987;
      19359: inst = 32'd136314880;
      19360: inst = 32'd268468224;
      19361: inst = 32'd201347784;
      19362: inst = 32'd203459665;
      19363: inst = 32'd136314880;
      19364: inst = 32'd268468224;
      19365: inst = 32'd201347785;
      19366: inst = 32'd203457519;
      19367: inst = 32'd136314880;
      19368: inst = 32'd268468224;
      19369: inst = 32'd201347786;
      19370: inst = 32'd203480697;
      19371: inst = 32'd136314880;
      19372: inst = 32'd268468224;
      19373: inst = 32'd201347787;
      19374: inst = 32'd203482841;
      19375: inst = 32'd136314880;
      19376: inst = 32'd268468224;
      19377: inst = 32'd201347788;
      19378: inst = 32'd203484922;
      19379: inst = 32'd136314880;
      19380: inst = 32'd268468224;
      19381: inst = 32'd201347789;
      19382: inst = 32'd203484889;
      19383: inst = 32'd136314880;
      19384: inst = 32'd268468224;
      19385: inst = 32'd201347790;
      19386: inst = 32'd203482776;
      19387: inst = 32'd136314880;
      19388: inst = 32'd268468224;
      19389: inst = 32'd201347791;
      19390: inst = 32'd203482776;
      19391: inst = 32'd136314880;
      19392: inst = 32'd268468224;
      19393: inst = 32'd201347792;
      19394: inst = 32'd203482808;
      19395: inst = 32'd136314880;
      19396: inst = 32'd268468224;
      19397: inst = 32'd201347793;
      19398: inst = 32'd203482808;
      19399: inst = 32'd136314880;
      19400: inst = 32'd268468224;
      19401: inst = 32'd201347794;
      19402: inst = 32'd203484889;
      19403: inst = 32'd136314880;
      19404: inst = 32'd268468224;
      19405: inst = 32'd201347795;
      19406: inst = 32'd203484954;
      19407: inst = 32'd136314880;
      19408: inst = 32'd268468224;
      19409: inst = 32'd201347796;
      19410: inst = 32'd203482842;
      19411: inst = 32'd136314880;
      19412: inst = 32'd268468224;
      19413: inst = 32'd201347797;
      19414: inst = 32'd203480729;
      19415: inst = 32'd136314880;
      19416: inst = 32'd268468224;
      19417: inst = 32'd201347798;
      19418: inst = 32'd203457519;
      19419: inst = 32'd136314880;
      19420: inst = 32'd268468224;
      19421: inst = 32'd201347799;
      19422: inst = 32'd203459665;
      19423: inst = 32'd136314880;
      19424: inst = 32'd268468224;
      19425: inst = 32'd201347800;
      19426: inst = 32'd203446987;
      19427: inst = 32'd136314880;
      19428: inst = 32'd268468224;
      19429: inst = 32'd201347801;
      19430: inst = 32'd203447020;
      19431: inst = 32'd136314880;
      19432: inst = 32'd268468224;
      19433: inst = 32'd201347802;
      19434: inst = 32'd203444906;
      19435: inst = 32'd136314880;
      19436: inst = 32'd268468224;
      19437: inst = 32'd201347803;
      19438: inst = 32'd203444874;
      19439: inst = 32'd136314880;
      19440: inst = 32'd268468224;
      19441: inst = 32'd201347804;
      19442: inst = 32'd203442794;
      19443: inst = 32'd136314880;
      19444: inst = 32'd268468224;
      19445: inst = 32'd201347805;
      19446: inst = 32'd203442794;
      19447: inst = 32'd136314880;
      19448: inst = 32'd268468224;
      19449: inst = 32'd201347806;
      19450: inst = 32'd203447019;
      19451: inst = 32'd136314880;
      19452: inst = 32'd268468224;
      19453: inst = 32'd201347807;
      19454: inst = 32'd203449100;
      19455: inst = 32'd136314880;
      19456: inst = 32'd268468224;
      19457: inst = 32'd201347808;
      19458: inst = 32'd203447020;
      19459: inst = 32'd136314880;
      19460: inst = 32'd268468224;
      19461: inst = 32'd201347809;
      19462: inst = 32'd203459665;
      19463: inst = 32'd136314880;
      19464: inst = 32'd268468224;
      19465: inst = 32'd201347810;
      19466: inst = 32'd203459600;
      19467: inst = 32'd136314880;
      19468: inst = 32'd268468224;
      19469: inst = 32'd201347811;
      19470: inst = 32'd203472245;
      19471: inst = 32'd136314880;
      19472: inst = 32'd268468224;
      19473: inst = 32'd201347812;
      19474: inst = 32'd203484857;
      19475: inst = 32'd136314880;
      19476: inst = 32'd268468224;
      19477: inst = 32'd201347813;
      19478: inst = 32'd203482743;
      19479: inst = 32'd136314880;
      19480: inst = 32'd268468224;
      19481: inst = 32'd201347814;
      19482: inst = 32'd203486969;
      19483: inst = 32'd136314880;
      19484: inst = 32'd268468224;
      19485: inst = 32'd201347815;
      19486: inst = 32'd203482776;
      19487: inst = 32'd136314880;
      19488: inst = 32'd268468224;
      19489: inst = 32'd201347816;
      19490: inst = 32'd203482809;
      19491: inst = 32'd136314880;
      19492: inst = 32'd268468224;
      19493: inst = 32'd201347817;
      19494: inst = 32'd203482810;
      19495: inst = 32'd136314880;
      19496: inst = 32'd268468224;
      19497: inst = 32'd201347818;
      19498: inst = 32'd203482810;
      19499: inst = 32'd136314880;
      19500: inst = 32'd268468224;
      19501: inst = 32'd201347819;
      19502: inst = 32'd203480729;
      19503: inst = 32'd136314880;
      19504: inst = 32'd268468224;
      19505: inst = 32'd201347820;
      19506: inst = 32'd203484857;
      19507: inst = 32'd136314880;
      19508: inst = 32'd268468224;
      19509: inst = 32'd201347821;
      19510: inst = 32'd203484823;
      19511: inst = 32'd136314880;
      19512: inst = 32'd268468224;
      19513: inst = 32'd201347822;
      19514: inst = 32'd203484693;
      19515: inst = 32'd136314880;
      19516: inst = 32'd268468224;
      19517: inst = 32'd201347823;
      19518: inst = 32'd203465675;
      19519: inst = 32'd136314880;
      19520: inst = 32'd268468224;
      19521: inst = 32'd201347824;
      19522: inst = 32'd203469574;
      19523: inst = 32'd136314880;
      19524: inst = 32'd268468224;
      19525: inst = 32'd201347825;
      19526: inst = 32'd203469574;
      19527: inst = 32'd136314880;
      19528: inst = 32'd268468224;
      19529: inst = 32'd201347826;
      19530: inst = 32'd203469574;
      19531: inst = 32'd136314880;
      19532: inst = 32'd268468224;
      19533: inst = 32'd201347827;
      19534: inst = 32'd203469574;
      19535: inst = 32'd136314880;
      19536: inst = 32'd268468224;
      19537: inst = 32'd201347828;
      19538: inst = 32'd203469574;
      19539: inst = 32'd136314880;
      19540: inst = 32'd268468224;
      19541: inst = 32'd201347829;
      19542: inst = 32'd203469574;
      19543: inst = 32'd136314880;
      19544: inst = 32'd268468224;
      19545: inst = 32'd201347830;
      19546: inst = 32'd203469574;
      19547: inst = 32'd136314880;
      19548: inst = 32'd268468224;
      19549: inst = 32'd201347831;
      19550: inst = 32'd203469574;
      19551: inst = 32'd136314880;
      19552: inst = 32'd268468224;
      19553: inst = 32'd201347832;
      19554: inst = 32'd203469606;
      19555: inst = 32'd136314880;
      19556: inst = 32'd268468224;
      19557: inst = 32'd201347833;
      19558: inst = 32'd203469574;
      19559: inst = 32'd136314880;
      19560: inst = 32'd268468224;
      19561: inst = 32'd201347834;
      19562: inst = 32'd203469574;
      19563: inst = 32'd136314880;
      19564: inst = 32'd268468224;
      19565: inst = 32'd201347835;
      19566: inst = 32'd203469606;
      19567: inst = 32'd136314880;
      19568: inst = 32'd268468224;
      19569: inst = 32'd201347836;
      19570: inst = 32'd203469574;
      19571: inst = 32'd136314880;
      19572: inst = 32'd268468224;
      19573: inst = 32'd201347837;
      19574: inst = 32'd203469606;
      19575: inst = 32'd136314880;
      19576: inst = 32'd268468224;
      19577: inst = 32'd201347838;
      19578: inst = 32'd203469606;
      19579: inst = 32'd136314880;
      19580: inst = 32'd268468224;
      19581: inst = 32'd201347839;
      19582: inst = 32'd203467493;
      19583: inst = 32'd136314880;
      19584: inst = 32'd268468224;
      19585: inst = 32'd201347840;
      19586: inst = 32'd203451279;
      19587: inst = 32'd136314880;
      19588: inst = 32'd268468224;
      19589: inst = 32'd201347841;
      19590: inst = 32'd203451247;
      19591: inst = 32'd136314880;
      19592: inst = 32'd268468224;
      19593: inst = 32'd201347842;
      19594: inst = 32'd203451247;
      19595: inst = 32'd136314880;
      19596: inst = 32'd268468224;
      19597: inst = 32'd201347843;
      19598: inst = 32'd203451247;
      19599: inst = 32'd136314880;
      19600: inst = 32'd268468224;
      19601: inst = 32'd201347844;
      19602: inst = 32'd203451215;
      19603: inst = 32'd136314880;
      19604: inst = 32'd268468224;
      19605: inst = 32'd201347845;
      19606: inst = 32'd203451215;
      19607: inst = 32'd136314880;
      19608: inst = 32'd268468224;
      19609: inst = 32'd201347846;
      19610: inst = 32'd203451247;
      19611: inst = 32'd136314880;
      19612: inst = 32'd268468224;
      19613: inst = 32'd201347847;
      19614: inst = 32'd203449134;
      19615: inst = 32'd136314880;
      19616: inst = 32'd268468224;
      19617: inst = 32'd201347848;
      19618: inst = 32'd203451247;
      19619: inst = 32'd136314880;
      19620: inst = 32'd268468224;
      19621: inst = 32'd201347849;
      19622: inst = 32'd203451215;
      19623: inst = 32'd136314880;
      19624: inst = 32'd268468224;
      19625: inst = 32'd201347850;
      19626: inst = 32'd203451247;
      19627: inst = 32'd136314880;
      19628: inst = 32'd268468224;
      19629: inst = 32'd201347851;
      19630: inst = 32'd203451247;
      19631: inst = 32'd136314880;
      19632: inst = 32'd268468224;
      19633: inst = 32'd201347852;
      19634: inst = 32'd203451215;
      19635: inst = 32'd136314880;
      19636: inst = 32'd268468224;
      19637: inst = 32'd201347853;
      19638: inst = 32'd203451247;
      19639: inst = 32'd136314880;
      19640: inst = 32'd268468224;
      19641: inst = 32'd201347854;
      19642: inst = 32'd203451215;
      19643: inst = 32'd136314880;
      19644: inst = 32'd268468224;
      19645: inst = 32'd201347855;
      19646: inst = 32'd203451247;
      19647: inst = 32'd136314880;
      19648: inst = 32'd268468224;
      19649: inst = 32'd201347856;
      19650: inst = 32'd203451311;
      19651: inst = 32'd136314880;
      19652: inst = 32'd268468224;
      19653: inst = 32'd201347857;
      19654: inst = 32'd203451279;
      19655: inst = 32'd136314880;
      19656: inst = 32'd268468224;
      19657: inst = 32'd201347858;
      19658: inst = 32'd203449167;
      19659: inst = 32'd136314880;
      19660: inst = 32'd268468224;
      19661: inst = 32'd201347859;
      19662: inst = 32'd203449134;
      19663: inst = 32'd136314880;
      19664: inst = 32'd268468224;
      19665: inst = 32'd201347860;
      19666: inst = 32'd203453296;
      19667: inst = 32'd136314880;
      19668: inst = 32'd268468224;
      19669: inst = 32'd201347861;
      19670: inst = 32'd203451182;
      19671: inst = 32'd136314880;
      19672: inst = 32'd268468224;
      19673: inst = 32'd201347862;
      19674: inst = 32'd203449036;
      19675: inst = 32'd136314880;
      19676: inst = 32'd268468224;
      19677: inst = 32'd201347863;
      19678: inst = 32'd203455375;
      19679: inst = 32'd136314880;
      19680: inst = 32'd268468224;
      19681: inst = 32'd201347864;
      19682: inst = 32'd203455406;
      19683: inst = 32'd136314880;
      19684: inst = 32'd268468224;
      19685: inst = 32'd201347865;
      19686: inst = 32'd203451147;
      19687: inst = 32'd136314880;
      19688: inst = 32'd268468224;
      19689: inst = 32'd201347866;
      19690: inst = 32'd203453292;
      19691: inst = 32'd136314880;
      19692: inst = 32'd268468224;
      19693: inst = 32'd201347867;
      19694: inst = 32'd203455438;
      19695: inst = 32'd136314880;
      19696: inst = 32'd268468224;
      19697: inst = 32'd201347868;
      19698: inst = 32'd203459664;
      19699: inst = 32'd136314880;
      19700: inst = 32'd268468224;
      19701: inst = 32'd201347869;
      19702: inst = 32'd203459665;
      19703: inst = 32'd136314880;
      19704: inst = 32'd268468224;
      19705: inst = 32'd201347870;
      19706: inst = 32'd203461779;
      19707: inst = 32'd136314880;
      19708: inst = 32'd268468224;
      19709: inst = 32'd201347871;
      19710: inst = 32'd203459666;
      19711: inst = 32'd136314880;
      19712: inst = 32'd268468224;
      19713: inst = 32'd201347872;
      19714: inst = 32'd203459665;
      19715: inst = 32'd136314880;
      19716: inst = 32'd268468224;
      19717: inst = 32'd201347873;
      19718: inst = 32'd203457519;
      19719: inst = 32'd136314880;
      19720: inst = 32'd268468224;
      19721: inst = 32'd201347874;
      19722: inst = 32'd203444874;
      19723: inst = 32'd136314880;
      19724: inst = 32'd268468224;
      19725: inst = 32'd201347875;
      19726: inst = 32'd203440648;
      19727: inst = 32'd136314880;
      19728: inst = 32'd268468224;
      19729: inst = 32'd201347876;
      19730: inst = 32'd203442761;
      19731: inst = 32'd136314880;
      19732: inst = 32'd268468224;
      19733: inst = 32'd201347877;
      19734: inst = 32'd203453326;
      19735: inst = 32'd136314880;
      19736: inst = 32'd268468224;
      19737: inst = 32'd201347878;
      19738: inst = 32'd203459665;
      19739: inst = 32'd136314880;
      19740: inst = 32'd268468224;
      19741: inst = 32'd201347879;
      19742: inst = 32'd203461778;
      19743: inst = 32'd136314880;
      19744: inst = 32'd268468224;
      19745: inst = 32'd201347880;
      19746: inst = 32'd203461778;
      19747: inst = 32'd136314880;
      19748: inst = 32'd268468224;
      19749: inst = 32'd201347881;
      19750: inst = 32'd203446987;
      19751: inst = 32'd136314880;
      19752: inst = 32'd268468224;
      19753: inst = 32'd201347882;
      19754: inst = 32'd203453358;
      19755: inst = 32'd136314880;
      19756: inst = 32'd268468224;
      19757: inst = 32'd201347883;
      19758: inst = 32'd203451180;
      19759: inst = 32'd136314880;
      19760: inst = 32'd268468224;
      19761: inst = 32'd201347884;
      19762: inst = 32'd203451180;
      19763: inst = 32'd136314880;
      19764: inst = 32'd268468224;
      19765: inst = 32'd201347885;
      19766: inst = 32'd203453260;
      19767: inst = 32'd136314880;
      19768: inst = 32'd268468224;
      19769: inst = 32'd201347886;
      19770: inst = 32'd203453261;
      19771: inst = 32'd136314880;
      19772: inst = 32'd268468224;
      19773: inst = 32'd201347887;
      19774: inst = 32'd203453293;
      19775: inst = 32'd136314880;
      19776: inst = 32'd268468224;
      19777: inst = 32'd201347888;
      19778: inst = 32'd203453293;
      19779: inst = 32'd136314880;
      19780: inst = 32'd268468224;
      19781: inst = 32'd201347889;
      19782: inst = 32'd203453261;
      19783: inst = 32'd136314880;
      19784: inst = 32'd268468224;
      19785: inst = 32'd201347890;
      19786: inst = 32'd203453260;
      19787: inst = 32'd136314880;
      19788: inst = 32'd268468224;
      19789: inst = 32'd201347891;
      19790: inst = 32'd203451180;
      19791: inst = 32'd136314880;
      19792: inst = 32'd268468224;
      19793: inst = 32'd201347892;
      19794: inst = 32'd203451180;
      19795: inst = 32'd136314880;
      19796: inst = 32'd268468224;
      19797: inst = 32'd201347893;
      19798: inst = 32'd203453358;
      19799: inst = 32'd136314880;
      19800: inst = 32'd268468224;
      19801: inst = 32'd201347894;
      19802: inst = 32'd203446987;
      19803: inst = 32'd136314880;
      19804: inst = 32'd268468224;
      19805: inst = 32'd201347895;
      19806: inst = 32'd203459697;
      19807: inst = 32'd136314880;
      19808: inst = 32'd268468224;
      19809: inst = 32'd201347896;
      19810: inst = 32'd203461778;
      19811: inst = 32'd136314880;
      19812: inst = 32'd268468224;
      19813: inst = 32'd201347897;
      19814: inst = 32'd203459665;
      19815: inst = 32'd136314880;
      19816: inst = 32'd268468224;
      19817: inst = 32'd201347898;
      19818: inst = 32'd203453326;
      19819: inst = 32'd136314880;
      19820: inst = 32'd268468224;
      19821: inst = 32'd201347899;
      19822: inst = 32'd203442761;
      19823: inst = 32'd136314880;
      19824: inst = 32'd268468224;
      19825: inst = 32'd201347900;
      19826: inst = 32'd203440648;
      19827: inst = 32'd136314880;
      19828: inst = 32'd268468224;
      19829: inst = 32'd201347901;
      19830: inst = 32'd203444874;
      19831: inst = 32'd136314880;
      19832: inst = 32'd268468224;
      19833: inst = 32'd201347902;
      19834: inst = 32'd203457519;
      19835: inst = 32'd136314880;
      19836: inst = 32'd268468224;
      19837: inst = 32'd201347903;
      19838: inst = 32'd203459665;
      19839: inst = 32'd136314880;
      19840: inst = 32'd268468224;
      19841: inst = 32'd201347904;
      19842: inst = 32'd203459666;
      19843: inst = 32'd136314880;
      19844: inst = 32'd268468224;
      19845: inst = 32'd201347905;
      19846: inst = 32'd203461812;
      19847: inst = 32'd136314880;
      19848: inst = 32'd268468224;
      19849: inst = 32'd201347906;
      19850: inst = 32'd203459633;
      19851: inst = 32'd136314880;
      19852: inst = 32'd268468224;
      19853: inst = 32'd201347907;
      19854: inst = 32'd203461681;
      19855: inst = 32'd136314880;
      19856: inst = 32'd268468224;
      19857: inst = 32'd201347908;
      19858: inst = 32'd203457454;
      19859: inst = 32'd136314880;
      19860: inst = 32'd268468224;
      19861: inst = 32'd201347909;
      19862: inst = 32'd203455309;
      19863: inst = 32'd136314880;
      19864: inst = 32'd268468224;
      19865: inst = 32'd201347910;
      19866: inst = 32'd203451148;
      19867: inst = 32'd136314880;
      19868: inst = 32'd268468224;
      19869: inst = 32'd201347911;
      19870: inst = 32'd203455375;
      19871: inst = 32'd136314880;
      19872: inst = 32'd268468224;
      19873: inst = 32'd201347912;
      19874: inst = 32'd203453295;
      19875: inst = 32'd136314880;
      19876: inst = 32'd268468224;
      19877: inst = 32'd201347913;
      19878: inst = 32'd203451214;
      19879: inst = 32'd136314880;
      19880: inst = 32'd268468224;
      19881: inst = 32'd201347914;
      19882: inst = 32'd203453295;
      19883: inst = 32'd136314880;
      19884: inst = 32'd268468224;
      19885: inst = 32'd201347915;
      19886: inst = 32'd203453295;
      19887: inst = 32'd136314880;
      19888: inst = 32'd268468224;
      19889: inst = 32'd201347916;
      19890: inst = 32'd203455375;
      19891: inst = 32'd136314880;
      19892: inst = 32'd268468224;
      19893: inst = 32'd201347917;
      19894: inst = 32'd203455310;
      19895: inst = 32'd136314880;
      19896: inst = 32'd268468224;
      19897: inst = 32'd201347918;
      19898: inst = 32'd203457390;
      19899: inst = 32'd136314880;
      19900: inst = 32'd268468224;
      19901: inst = 32'd201347919;
      19902: inst = 32'd203453131;
      19903: inst = 32'd136314880;
      19904: inst = 32'd268468224;
      19905: inst = 32'd201347920;
      19906: inst = 32'd203457323;
      19907: inst = 32'd136314880;
      19908: inst = 32'd268468224;
      19909: inst = 32'd201347921;
      19910: inst = 32'd203457323;
      19911: inst = 32'd136314880;
      19912: inst = 32'd268468224;
      19913: inst = 32'd201347922;
      19914: inst = 32'd203457323;
      19915: inst = 32'd136314880;
      19916: inst = 32'd268468224;
      19917: inst = 32'd201347923;
      19918: inst = 32'd203457323;
      19919: inst = 32'd136314880;
      19920: inst = 32'd268468224;
      19921: inst = 32'd201347924;
      19922: inst = 32'd203457323;
      19923: inst = 32'd136314880;
      19924: inst = 32'd268468224;
      19925: inst = 32'd201347925;
      19926: inst = 32'd203457323;
      19927: inst = 32'd136314880;
      19928: inst = 32'd268468224;
      19929: inst = 32'd201347926;
      19930: inst = 32'd203457323;
      19931: inst = 32'd136314880;
      19932: inst = 32'd268468224;
      19933: inst = 32'd201347927;
      19934: inst = 32'd203457323;
      19935: inst = 32'd136314880;
      19936: inst = 32'd268468224;
      19937: inst = 32'd201347928;
      19938: inst = 32'd203457323;
      19939: inst = 32'd136314880;
      19940: inst = 32'd268468224;
      19941: inst = 32'd201347929;
      19942: inst = 32'd203455242;
      19943: inst = 32'd136314880;
      19944: inst = 32'd268468224;
      19945: inst = 32'd201347930;
      19946: inst = 32'd203457291;
      19947: inst = 32'd136314880;
      19948: inst = 32'd268468224;
      19949: inst = 32'd201347931;
      19950: inst = 32'd203457323;
      19951: inst = 32'd136314880;
      19952: inst = 32'd268468224;
      19953: inst = 32'd201347932;
      19954: inst = 32'd203457291;
      19955: inst = 32'd136314880;
      19956: inst = 32'd268468224;
      19957: inst = 32'd201347933;
      19958: inst = 32'd203457291;
      19959: inst = 32'd136314880;
      19960: inst = 32'd268468224;
      19961: inst = 32'd201347934;
      19962: inst = 32'd203457323;
      19963: inst = 32'd136314880;
      19964: inst = 32'd268468224;
      19965: inst = 32'd201347935;
      19966: inst = 32'd203457323;
      19967: inst = 32'd136314880;
      19968: inst = 32'd268468224;
      19969: inst = 32'd201347936;
      19970: inst = 32'd203451247;
      19971: inst = 32'd136314880;
      19972: inst = 32'd268468224;
      19973: inst = 32'd201347937;
      19974: inst = 32'd203449135;
      19975: inst = 32'd136314880;
      19976: inst = 32'd268468224;
      19977: inst = 32'd201347938;
      19978: inst = 32'd203451215;
      19979: inst = 32'd136314880;
      19980: inst = 32'd268468224;
      19981: inst = 32'd201347939;
      19982: inst = 32'd203451247;
      19983: inst = 32'd136314880;
      19984: inst = 32'd268468224;
      19985: inst = 32'd201347940;
      19986: inst = 32'd203451215;
      19987: inst = 32'd136314880;
      19988: inst = 32'd268468224;
      19989: inst = 32'd201347941;
      19990: inst = 32'd203451247;
      19991: inst = 32'd136314880;
      19992: inst = 32'd268468224;
      19993: inst = 32'd201347942;
      19994: inst = 32'd203451247;
      19995: inst = 32'd136314880;
      19996: inst = 32'd268468224;
      19997: inst = 32'd201347943;
      19998: inst = 32'd203451247;
      19999: inst = 32'd136314880;
      20000: inst = 32'd268468224;
      20001: inst = 32'd201347944;
      20002: inst = 32'd203451247;
      20003: inst = 32'd136314880;
      20004: inst = 32'd268468224;
      20005: inst = 32'd201347945;
      20006: inst = 32'd203451215;
      20007: inst = 32'd136314880;
      20008: inst = 32'd268468224;
      20009: inst = 32'd201347946;
      20010: inst = 32'd203451280;
      20011: inst = 32'd136314880;
      20012: inst = 32'd268468224;
      20013: inst = 32'd201347947;
      20014: inst = 32'd203449167;
      20015: inst = 32'd136314880;
      20016: inst = 32'd268468224;
      20017: inst = 32'd201347948;
      20018: inst = 32'd203451215;
      20019: inst = 32'd136314880;
      20020: inst = 32'd268468224;
      20021: inst = 32'd201347949;
      20022: inst = 32'd203451247;
      20023: inst = 32'd136314880;
      20024: inst = 32'd268468224;
      20025: inst = 32'd201347950;
      20026: inst = 32'd203451215;
      20027: inst = 32'd136314880;
      20028: inst = 32'd268468224;
      20029: inst = 32'd201347951;
      20030: inst = 32'd203451215;
      20031: inst = 32'd136314880;
      20032: inst = 32'd268468224;
      20033: inst = 32'd201347952;
      20034: inst = 32'd203447086;
      20035: inst = 32'd136314880;
      20036: inst = 32'd268468224;
      20037: inst = 32'd201347953;
      20038: inst = 32'd203451247;
      20039: inst = 32'd136314880;
      20040: inst = 32'd268468224;
      20041: inst = 32'd201347954;
      20042: inst = 32'd203451280;
      20043: inst = 32'd136314880;
      20044: inst = 32'd268468224;
      20045: inst = 32'd201347955;
      20046: inst = 32'd203449136;
      20047: inst = 32'd136314880;
      20048: inst = 32'd268468224;
      20049: inst = 32'd201347956;
      20050: inst = 32'd203451249;
      20051: inst = 32'd136314880;
      20052: inst = 32'd268468224;
      20053: inst = 32'd201347957;
      20054: inst = 32'd203453329;
      20055: inst = 32'd136314880;
      20056: inst = 32'd268468224;
      20057: inst = 32'd201347958;
      20058: inst = 32'd203451215;
      20059: inst = 32'd136314880;
      20060: inst = 32'd268468224;
      20061: inst = 32'd201347959;
      20062: inst = 32'd203453295;
      20063: inst = 32'd136314880;
      20064: inst = 32'd268468224;
      20065: inst = 32'd201347960;
      20066: inst = 32'd203451214;
      20067: inst = 32'd136314880;
      20068: inst = 32'd268468224;
      20069: inst = 32'd201347961;
      20070: inst = 32'd203451213;
      20071: inst = 32'd136314880;
      20072: inst = 32'd268468224;
      20073: inst = 32'd201347962;
      20074: inst = 32'd203453325;
      20075: inst = 32'd136314880;
      20076: inst = 32'd268468224;
      20077: inst = 32'd201347963;
      20078: inst = 32'd203461810;
      20079: inst = 32'd136314880;
      20080: inst = 32'd268468224;
      20081: inst = 32'd201347964;
      20082: inst = 32'd203459632;
      20083: inst = 32'd136314880;
      20084: inst = 32'd268468224;
      20085: inst = 32'd201347965;
      20086: inst = 32'd203457585;
      20087: inst = 32'd136314880;
      20088: inst = 32'd268468224;
      20089: inst = 32'd201347966;
      20090: inst = 32'd203442762;
      20091: inst = 32'd136314880;
      20092: inst = 32'd268468224;
      20093: inst = 32'd201347967;
      20094: inst = 32'd203444843;
      20095: inst = 32'd136314880;
      20096: inst = 32'd268468224;
      20097: inst = 32'd201347968;
      20098: inst = 32'd203446987;
      20099: inst = 32'd136314880;
      20100: inst = 32'd268468224;
      20101: inst = 32'd201347969;
      20102: inst = 32'd203453293;
      20103: inst = 32'd136314880;
      20104: inst = 32'd268468224;
      20105: inst = 32'd201347970;
      20106: inst = 32'd203444842;
      20107: inst = 32'd136314880;
      20108: inst = 32'd268468224;
      20109: inst = 32'd201347971;
      20110: inst = 32'd203444874;
      20111: inst = 32'd136314880;
      20112: inst = 32'd268468224;
      20113: inst = 32'd201347972;
      20114: inst = 32'd203444874;
      20115: inst = 32'd136314880;
      20116: inst = 32'd268468224;
      20117: inst = 32'd201347973;
      20118: inst = 32'd203457552;
      20119: inst = 32'd136314880;
      20120: inst = 32'd268468224;
      20121: inst = 32'd201347974;
      20122: inst = 32'd203459665;
      20123: inst = 32'd136314880;
      20124: inst = 32'd268468224;
      20125: inst = 32'd201347975;
      20126: inst = 32'd203459697;
      20127: inst = 32'd136314880;
      20128: inst = 32'd268468224;
      20129: inst = 32'd201347976;
      20130: inst = 32'd203459697;
      20131: inst = 32'd136314880;
      20132: inst = 32'd268468224;
      20133: inst = 32'd201347977;
      20134: inst = 32'd203444907;
      20135: inst = 32'd136314880;
      20136: inst = 32'd268468224;
      20137: inst = 32'd201347978;
      20138: inst = 32'd203451246;
      20139: inst = 32'd136314880;
      20140: inst = 32'd268468224;
      20141: inst = 32'd201347979;
      20142: inst = 32'd203451246;
      20143: inst = 32'd136314880;
      20144: inst = 32'd268468224;
      20145: inst = 32'd201347980;
      20146: inst = 32'd203451279;
      20147: inst = 32'd136314880;
      20148: inst = 32'd268468224;
      20149: inst = 32'd201347981;
      20150: inst = 32'd203453327;
      20151: inst = 32'd136314880;
      20152: inst = 32'd268468224;
      20153: inst = 32'd201347982;
      20154: inst = 32'd203451247;
      20155: inst = 32'd136314880;
      20156: inst = 32'd268468224;
      20157: inst = 32'd201347983;
      20158: inst = 32'd203449166;
      20159: inst = 32'd136314880;
      20160: inst = 32'd268468224;
      20161: inst = 32'd201347984;
      20162: inst = 32'd203449166;
      20163: inst = 32'd136314880;
      20164: inst = 32'd268468224;
      20165: inst = 32'd201347985;
      20166: inst = 32'd203451247;
      20167: inst = 32'd136314880;
      20168: inst = 32'd268468224;
      20169: inst = 32'd201347986;
      20170: inst = 32'd203451279;
      20171: inst = 32'd136314880;
      20172: inst = 32'd268468224;
      20173: inst = 32'd201347987;
      20174: inst = 32'd203451279;
      20175: inst = 32'd136314880;
      20176: inst = 32'd268468224;
      20177: inst = 32'd201347988;
      20178: inst = 32'd203451246;
      20179: inst = 32'd136314880;
      20180: inst = 32'd268468224;
      20181: inst = 32'd201347989;
      20182: inst = 32'd203451246;
      20183: inst = 32'd136314880;
      20184: inst = 32'd268468224;
      20185: inst = 32'd201347990;
      20186: inst = 32'd203444907;
      20187: inst = 32'd136314880;
      20188: inst = 32'd268468224;
      20189: inst = 32'd201347991;
      20190: inst = 32'd203457617;
      20191: inst = 32'd136314880;
      20192: inst = 32'd268468224;
      20193: inst = 32'd201347992;
      20194: inst = 32'd203459697;
      20195: inst = 32'd136314880;
      20196: inst = 32'd268468224;
      20197: inst = 32'd201347993;
      20198: inst = 32'd203459665;
      20199: inst = 32'd136314880;
      20200: inst = 32'd268468224;
      20201: inst = 32'd201347994;
      20202: inst = 32'd203457552;
      20203: inst = 32'd136314880;
      20204: inst = 32'd268468224;
      20205: inst = 32'd201347995;
      20206: inst = 32'd203444874;
      20207: inst = 32'd136314880;
      20208: inst = 32'd268468224;
      20209: inst = 32'd201347996;
      20210: inst = 32'd203444874;
      20211: inst = 32'd136314880;
      20212: inst = 32'd268468224;
      20213: inst = 32'd201347997;
      20214: inst = 32'd203444842;
      20215: inst = 32'd136314880;
      20216: inst = 32'd268468224;
      20217: inst = 32'd201347998;
      20218: inst = 32'd203453293;
      20219: inst = 32'd136314880;
      20220: inst = 32'd268468224;
      20221: inst = 32'd201347999;
      20222: inst = 32'd203446987;
      20223: inst = 32'd136314880;
      20224: inst = 32'd268468224;
      20225: inst = 32'd201348000;
      20226: inst = 32'd203442796;
      20227: inst = 32'd136314880;
      20228: inst = 32'd268468224;
      20229: inst = 32'd201348001;
      20230: inst = 32'd203442763;
      20231: inst = 32'd136314880;
      20232: inst = 32'd268468224;
      20233: inst = 32'd201348002;
      20234: inst = 32'd203457585;
      20235: inst = 32'd136314880;
      20236: inst = 32'd268468224;
      20237: inst = 32'd201348003;
      20238: inst = 32'd203459633;
      20239: inst = 32'd136314880;
      20240: inst = 32'd268468224;
      20241: inst = 32'd201348004;
      20242: inst = 32'd203463826;
      20243: inst = 32'd136314880;
      20244: inst = 32'd268468224;
      20245: inst = 32'd201348005;
      20246: inst = 32'd203455342;
      20247: inst = 32'd136314880;
      20248: inst = 32'd268468224;
      20249: inst = 32'd201348006;
      20250: inst = 32'd203451182;
      20251: inst = 32'd136314880;
      20252: inst = 32'd268468224;
      20253: inst = 32'd201348007;
      20254: inst = 32'd203451215;
      20255: inst = 32'd136314880;
      20256: inst = 32'd268468224;
      20257: inst = 32'd201348008;
      20258: inst = 32'd203451247;
      20259: inst = 32'd136314880;
      20260: inst = 32'd268468224;
      20261: inst = 32'd201348009;
      20262: inst = 32'd203449136;
      20263: inst = 32'd136314880;
      20264: inst = 32'd268468224;
      20265: inst = 32'd201348010;
      20266: inst = 32'd203449169;
      20267: inst = 32'd136314880;
      20268: inst = 32'd268468224;
      20269: inst = 32'd201348011;
      20270: inst = 32'd203449168;
      20271: inst = 32'd136314880;
      20272: inst = 32'd268468224;
      20273: inst = 32'd201348012;
      20274: inst = 32'd203451216;
      20275: inst = 32'd136314880;
      20276: inst = 32'd268468224;
      20277: inst = 32'd201348013;
      20278: inst = 32'd203449103;
      20279: inst = 32'd136314880;
      20280: inst = 32'd268468224;
      20281: inst = 32'd201348014;
      20282: inst = 32'd203453264;
      20283: inst = 32'd136314880;
      20284: inst = 32'd268468224;
      20285: inst = 32'd201348015;
      20286: inst = 32'd203455344;
      20287: inst = 32'd136314880;
      20288: inst = 32'd268468224;
      20289: inst = 32'd201348016;
      20290: inst = 32'd203449233;
      20291: inst = 32'd136314880;
      20292: inst = 32'd268468224;
      20293: inst = 32'd201348017;
      20294: inst = 32'd203449233;
      20295: inst = 32'd136314880;
      20296: inst = 32'd268468224;
      20297: inst = 32'd201348018;
      20298: inst = 32'd203449233;
      20299: inst = 32'd136314880;
      20300: inst = 32'd268468224;
      20301: inst = 32'd201348019;
      20302: inst = 32'd203449233;
      20303: inst = 32'd136314880;
      20304: inst = 32'd268468224;
      20305: inst = 32'd201348020;
      20306: inst = 32'd203449233;
      20307: inst = 32'd136314880;
      20308: inst = 32'd268468224;
      20309: inst = 32'd201348021;
      20310: inst = 32'd203449233;
      20311: inst = 32'd136314880;
      20312: inst = 32'd268468224;
      20313: inst = 32'd201348022;
      20314: inst = 32'd203449233;
      20315: inst = 32'd136314880;
      20316: inst = 32'd268468224;
      20317: inst = 32'd201348023;
      20318: inst = 32'd203449233;
      20319: inst = 32'd136314880;
      20320: inst = 32'd268468224;
      20321: inst = 32'd201348024;
      20322: inst = 32'd203449233;
      20323: inst = 32'd136314880;
      20324: inst = 32'd268468224;
      20325: inst = 32'd201348025;
      20326: inst = 32'd203449200;
      20327: inst = 32'd136314880;
      20328: inst = 32'd268468224;
      20329: inst = 32'd201348026;
      20330: inst = 32'd203449201;
      20331: inst = 32'd136314880;
      20332: inst = 32'd268468224;
      20333: inst = 32'd201348027;
      20334: inst = 32'd203449233;
      20335: inst = 32'd136314880;
      20336: inst = 32'd268468224;
      20337: inst = 32'd201348028;
      20338: inst = 32'd203449201;
      20339: inst = 32'd136314880;
      20340: inst = 32'd268468224;
      20341: inst = 32'd201348029;
      20342: inst = 32'd203449201;
      20343: inst = 32'd136314880;
      20344: inst = 32'd268468224;
      20345: inst = 32'd201348030;
      20346: inst = 32'd203449233;
      20347: inst = 32'd136314880;
      20348: inst = 32'd268468224;
      20349: inst = 32'd201348031;
      20350: inst = 32'd203449233;
      20351: inst = 32'd136314880;
      20352: inst = 32'd268468224;
      20353: inst = 32'd201348032;
      20354: inst = 32'd203451248;
      20355: inst = 32'd136314880;
      20356: inst = 32'd268468224;
      20357: inst = 32'd201348033;
      20358: inst = 32'd203449135;
      20359: inst = 32'd136314880;
      20360: inst = 32'd268468224;
      20361: inst = 32'd201348034;
      20362: inst = 32'd203451248;
      20363: inst = 32'd136314880;
      20364: inst = 32'd268468224;
      20365: inst = 32'd201348035;
      20366: inst = 32'd203451248;
      20367: inst = 32'd136314880;
      20368: inst = 32'd268468224;
      20369: inst = 32'd201348036;
      20370: inst = 32'd203449167;
      20371: inst = 32'd136314880;
      20372: inst = 32'd268468224;
      20373: inst = 32'd201348037;
      20374: inst = 32'd203451248;
      20375: inst = 32'd136314880;
      20376: inst = 32'd268468224;
      20377: inst = 32'd201348038;
      20378: inst = 32'd203451215;
      20379: inst = 32'd136314880;
      20380: inst = 32'd268468224;
      20381: inst = 32'd201348039;
      20382: inst = 32'd203451248;
      20383: inst = 32'd136314880;
      20384: inst = 32'd268468224;
      20385: inst = 32'd201348040;
      20386: inst = 32'd203451216;
      20387: inst = 32'd136314880;
      20388: inst = 32'd268468224;
      20389: inst = 32'd201348041;
      20390: inst = 32'd203449167;
      20391: inst = 32'd136314880;
      20392: inst = 32'd268468224;
      20393: inst = 32'd201348042;
      20394: inst = 32'd203451248;
      20395: inst = 32'd136314880;
      20396: inst = 32'd268468224;
      20397: inst = 32'd201348043;
      20398: inst = 32'd203449167;
      20399: inst = 32'd136314880;
      20400: inst = 32'd268468224;
      20401: inst = 32'd201348044;
      20402: inst = 32'd203451216;
      20403: inst = 32'd136314880;
      20404: inst = 32'd268468224;
      20405: inst = 32'd201348045;
      20406: inst = 32'd203451248;
      20407: inst = 32'd136314880;
      20408: inst = 32'd268468224;
      20409: inst = 32'd201348046;
      20410: inst = 32'd203451215;
      20411: inst = 32'd136314880;
      20412: inst = 32'd268468224;
      20413: inst = 32'd201348047;
      20414: inst = 32'd203451215;
      20415: inst = 32'd136314880;
      20416: inst = 32'd268468224;
      20417: inst = 32'd201348048;
      20418: inst = 32'd203449199;
      20419: inst = 32'd136314880;
      20420: inst = 32'd268468224;
      20421: inst = 32'd201348049;
      20422: inst = 32'd203449200;
      20423: inst = 32'd136314880;
      20424: inst = 32'd268468224;
      20425: inst = 32'd201348050;
      20426: inst = 32'd203451248;
      20427: inst = 32'd136314880;
      20428: inst = 32'd268468224;
      20429: inst = 32'd201348051;
      20430: inst = 32'd203449168;
      20431: inst = 32'd136314880;
      20432: inst = 32'd268468224;
      20433: inst = 32'd201348052;
      20434: inst = 32'd203449169;
      20435: inst = 32'd136314880;
      20436: inst = 32'd268468224;
      20437: inst = 32'd201348053;
      20438: inst = 32'd203449168;
      20439: inst = 32'd136314880;
      20440: inst = 32'd268468224;
      20441: inst = 32'd201348054;
      20442: inst = 32'd203449136;
      20443: inst = 32'd136314880;
      20444: inst = 32'd268468224;
      20445: inst = 32'd201348055;
      20446: inst = 32'd203449167;
      20447: inst = 32'd136314880;
      20448: inst = 32'd268468224;
      20449: inst = 32'd201348056;
      20450: inst = 32'd203451247;
      20451: inst = 32'd136314880;
      20452: inst = 32'd268468224;
      20453: inst = 32'd201348057;
      20454: inst = 32'd203453359;
      20455: inst = 32'd136314880;
      20456: inst = 32'd268468224;
      20457: inst = 32'd201348058;
      20458: inst = 32'd203459665;
      20459: inst = 32'd136314880;
      20460: inst = 32'd268468224;
      20461: inst = 32'd201348059;
      20462: inst = 32'd203459665;
      20463: inst = 32'd136314880;
      20464: inst = 32'd268468224;
      20465: inst = 32'd201348060;
      20466: inst = 32'd203459698;
      20467: inst = 32'd136314880;
      20468: inst = 32'd268468224;
      20469: inst = 32'd201348061;
      20470: inst = 32'd203446955;
      20471: inst = 32'd136314880;
      20472: inst = 32'd268468224;
      20473: inst = 32'd201348062;
      20474: inst = 32'd203442794;
      20475: inst = 32'd136314880;
      20476: inst = 32'd268468224;
      20477: inst = 32'd201348063;
      20478: inst = 32'd203442795;
      20479: inst = 32'd136314880;
      20480: inst = 32'd268468224;
      20481: inst = 32'd201348064;
      20482: inst = 32'd203453326;
      20483: inst = 32'd136314880;
      20484: inst = 32'd268468224;
      20485: inst = 32'd201348065;
      20486: inst = 32'd203457487;
      20487: inst = 32'd136314880;
      20488: inst = 32'd268468224;
      20489: inst = 32'd201348066;
      20490: inst = 32'd203444874;
      20491: inst = 32'd136314880;
      20492: inst = 32'd268468224;
      20493: inst = 32'd201348067;
      20494: inst = 32'd203444841;
      20495: inst = 32'd136314880;
      20496: inst = 32'd268468224;
      20497: inst = 32'd201348068;
      20498: inst = 32'd203446986;
      20499: inst = 32'd136314880;
      20500: inst = 32'd268468224;
      20501: inst = 32'd201348069;
      20502: inst = 32'd203459665;
      20503: inst = 32'd136314880;
      20504: inst = 32'd268468224;
      20505: inst = 32'd201348070;
      20506: inst = 32'd203459697;
      20507: inst = 32'd136314880;
      20508: inst = 32'd268468224;
      20509: inst = 32'd201348071;
      20510: inst = 32'd203459697;
      20511: inst = 32'd136314880;
      20512: inst = 32'd268468224;
      20513: inst = 32'd201348072;
      20514: inst = 32'd203457585;
      20515: inst = 32'd136314880;
      20516: inst = 32'd268468224;
      20517: inst = 32'd201348073;
      20518: inst = 32'd203444939;
      20519: inst = 32'd136314880;
      20520: inst = 32'd268468224;
      20521: inst = 32'd201348074;
      20522: inst = 32'd203449198;
      20523: inst = 32'd136314880;
      20524: inst = 32'd268468224;
      20525: inst = 32'd201348075;
      20526: inst = 32'd203449199;
      20527: inst = 32'd136314880;
      20528: inst = 32'd268468224;
      20529: inst = 32'd201348076;
      20530: inst = 32'd203449167;
      20531: inst = 32'd136314880;
      20532: inst = 32'd268468224;
      20533: inst = 32'd201348077;
      20534: inst = 32'd203449167;
      20535: inst = 32'd136314880;
      20536: inst = 32'd268468224;
      20537: inst = 32'd201348078;
      20538: inst = 32'd203449168;
      20539: inst = 32'd136314880;
      20540: inst = 32'd268468224;
      20541: inst = 32'd201348079;
      20542: inst = 32'd203449200;
      20543: inst = 32'd136314880;
      20544: inst = 32'd268468224;
      20545: inst = 32'd201348080;
      20546: inst = 32'd203449200;
      20547: inst = 32'd136314880;
      20548: inst = 32'd268468224;
      20549: inst = 32'd201348081;
      20550: inst = 32'd203449200;
      20551: inst = 32'd136314880;
      20552: inst = 32'd268468224;
      20553: inst = 32'd201348082;
      20554: inst = 32'd203449168;
      20555: inst = 32'd136314880;
      20556: inst = 32'd268468224;
      20557: inst = 32'd201348083;
      20558: inst = 32'd203449199;
      20559: inst = 32'd136314880;
      20560: inst = 32'd268468224;
      20561: inst = 32'd201348084;
      20562: inst = 32'd203449199;
      20563: inst = 32'd136314880;
      20564: inst = 32'd268468224;
      20565: inst = 32'd201348085;
      20566: inst = 32'd203449199;
      20567: inst = 32'd136314880;
      20568: inst = 32'd268468224;
      20569: inst = 32'd201348086;
      20570: inst = 32'd203444940;
      20571: inst = 32'd136314880;
      20572: inst = 32'd268468224;
      20573: inst = 32'd201348087;
      20574: inst = 32'd203457617;
      20575: inst = 32'd136314880;
      20576: inst = 32'd268468224;
      20577: inst = 32'd201348088;
      20578: inst = 32'd203459697;
      20579: inst = 32'd136314880;
      20580: inst = 32'd268468224;
      20581: inst = 32'd201348089;
      20582: inst = 32'd203459697;
      20583: inst = 32'd136314880;
      20584: inst = 32'd268468224;
      20585: inst = 32'd201348090;
      20586: inst = 32'd203459665;
      20587: inst = 32'd136314880;
      20588: inst = 32'd268468224;
      20589: inst = 32'd201348091;
      20590: inst = 32'd203446986;
      20591: inst = 32'd136314880;
      20592: inst = 32'd268468224;
      20593: inst = 32'd201348092;
      20594: inst = 32'd203444841;
      20595: inst = 32'd136314880;
      20596: inst = 32'd268468224;
      20597: inst = 32'd201348093;
      20598: inst = 32'd203444874;
      20599: inst = 32'd136314880;
      20600: inst = 32'd268468224;
      20601: inst = 32'd201348094;
      20602: inst = 32'd203457487;
      20603: inst = 32'd136314880;
      20604: inst = 32'd268468224;
      20605: inst = 32'd201348095;
      20606: inst = 32'd203453326;
      20607: inst = 32'd136314880;
      20608: inst = 32'd268468224;
      20609: inst = 32'd201348096;
      20610: inst = 32'd203442795;
      20611: inst = 32'd136314880;
      20612: inst = 32'd268468224;
      20613: inst = 32'd201348097;
      20614: inst = 32'd203442762;
      20615: inst = 32'd136314880;
      20616: inst = 32'd268468224;
      20617: inst = 32'd201348098;
      20618: inst = 32'd203446988;
      20619: inst = 32'd136314880;
      20620: inst = 32'd268468224;
      20621: inst = 32'd201348099;
      20622: inst = 32'd203459665;
      20623: inst = 32'd136314880;
      20624: inst = 32'd268468224;
      20625: inst = 32'd201348100;
      20626: inst = 32'd203459633;
      20627: inst = 32'd136314880;
      20628: inst = 32'd268468224;
      20629: inst = 32'd201348101;
      20630: inst = 32'd203459666;
      20631: inst = 32'd136314880;
      20632: inst = 32'd268468224;
      20633: inst = 32'd201348102;
      20634: inst = 32'd203453327;
      20635: inst = 32'd136314880;
      20636: inst = 32'd268468224;
      20637: inst = 32'd201348103;
      20638: inst = 32'd203451215;
      20639: inst = 32'd136314880;
      20640: inst = 32'd268468224;
      20641: inst = 32'd201348104;
      20642: inst = 32'd203451280;
      20643: inst = 32'd136314880;
      20644: inst = 32'd268468224;
      20645: inst = 32'd201348105;
      20646: inst = 32'd203451281;
      20647: inst = 32'd136314880;
      20648: inst = 32'd268468224;
      20649: inst = 32'd201348106;
      20650: inst = 32'd203449234;
      20651: inst = 32'd136314880;
      20652: inst = 32'd268468224;
      20653: inst = 32'd201348107;
      20654: inst = 32'd203449202;
      20655: inst = 32'd136314880;
      20656: inst = 32'd268468224;
      20657: inst = 32'd201348108;
      20658: inst = 32'd203449202;
      20659: inst = 32'd136314880;
      20660: inst = 32'd268468224;
      20661: inst = 32'd201348109;
      20662: inst = 32'd203449169;
      20663: inst = 32'd136314880;
      20664: inst = 32'd268468224;
      20665: inst = 32'd201348110;
      20666: inst = 32'd203451217;
      20667: inst = 32'd136314880;
      20668: inst = 32'd268468224;
      20669: inst = 32'd201348111;
      20670: inst = 32'd203449104;
      20671: inst = 32'd136314880;
      20672: inst = 32'd268468224;
      20673: inst = 32'd201348112;
      20674: inst = 32'd203447154;
      20675: inst = 32'd136314880;
      20676: inst = 32'd268468224;
      20677: inst = 32'd201348113;
      20678: inst = 32'd203447154;
      20679: inst = 32'd136314880;
      20680: inst = 32'd268468224;
      20681: inst = 32'd201348114;
      20682: inst = 32'd203447154;
      20683: inst = 32'd136314880;
      20684: inst = 32'd268468224;
      20685: inst = 32'd201348115;
      20686: inst = 32'd203447154;
      20687: inst = 32'd136314880;
      20688: inst = 32'd268468224;
      20689: inst = 32'd201348116;
      20690: inst = 32'd203447154;
      20691: inst = 32'd136314880;
      20692: inst = 32'd268468224;
      20693: inst = 32'd201348117;
      20694: inst = 32'd203447154;
      20695: inst = 32'd136314880;
      20696: inst = 32'd268468224;
      20697: inst = 32'd201348118;
      20698: inst = 32'd203447154;
      20699: inst = 32'd136314880;
      20700: inst = 32'd268468224;
      20701: inst = 32'd201348119;
      20702: inst = 32'd203447154;
      20703: inst = 32'd136314880;
      20704: inst = 32'd268468224;
      20705: inst = 32'd201348120;
      20706: inst = 32'd203447186;
      20707: inst = 32'd136314880;
      20708: inst = 32'd268468224;
      20709: inst = 32'd201348121;
      20710: inst = 32'd203445105;
      20711: inst = 32'd136314880;
      20712: inst = 32'd268468224;
      20713: inst = 32'd201348122;
      20714: inst = 32'd203447154;
      20715: inst = 32'd136314880;
      20716: inst = 32'd268468224;
      20717: inst = 32'd201348123;
      20718: inst = 32'd203447186;
      20719: inst = 32'd136314880;
      20720: inst = 32'd268468224;
      20721: inst = 32'd201348124;
      20722: inst = 32'd203445106;
      20723: inst = 32'd136314880;
      20724: inst = 32'd268468224;
      20725: inst = 32'd201348125;
      20726: inst = 32'd203445106;
      20727: inst = 32'd136314880;
      20728: inst = 32'd268468224;
      20729: inst = 32'd201348126;
      20730: inst = 32'd203447186;
      20731: inst = 32'd136314880;
      20732: inst = 32'd268468224;
      20733: inst = 32'd201348127;
      20734: inst = 32'd203445106;
      20735: inst = 32'd136314880;
      20736: inst = 32'd268468224;
      20737: inst = 32'd201348128;
      20738: inst = 32'd203451248;
      20739: inst = 32'd136314880;
      20740: inst = 32'd268468224;
      20741: inst = 32'd201348129;
      20742: inst = 32'd203449168;
      20743: inst = 32'd136314880;
      20744: inst = 32'd268468224;
      20745: inst = 32'd201348130;
      20746: inst = 32'd203451248;
      20747: inst = 32'd136314880;
      20748: inst = 32'd268468224;
      20749: inst = 32'd201348131;
      20750: inst = 32'd203451216;
      20751: inst = 32'd136314880;
      20752: inst = 32'd268468224;
      20753: inst = 32'd201348132;
      20754: inst = 32'd203449167;
      20755: inst = 32'd136314880;
      20756: inst = 32'd268468224;
      20757: inst = 32'd201348133;
      20758: inst = 32'd203451248;
      20759: inst = 32'd136314880;
      20760: inst = 32'd268468224;
      20761: inst = 32'd201348134;
      20762: inst = 32'd203449135;
      20763: inst = 32'd136314880;
      20764: inst = 32'd268468224;
      20765: inst = 32'd201348135;
      20766: inst = 32'd203451216;
      20767: inst = 32'd136314880;
      20768: inst = 32'd268468224;
      20769: inst = 32'd201348136;
      20770: inst = 32'd203451216;
      20771: inst = 32'd136314880;
      20772: inst = 32'd268468224;
      20773: inst = 32'd201348137;
      20774: inst = 32'd203451216;
      20775: inst = 32'd136314880;
      20776: inst = 32'd268468224;
      20777: inst = 32'd201348138;
      20778: inst = 32'd203449167;
      20779: inst = 32'd136314880;
      20780: inst = 32'd268468224;
      20781: inst = 32'd201348139;
      20782: inst = 32'd203451248;
      20783: inst = 32'd136314880;
      20784: inst = 32'd268468224;
      20785: inst = 32'd201348140;
      20786: inst = 32'd203451216;
      20787: inst = 32'd136314880;
      20788: inst = 32'd268468224;
      20789: inst = 32'd201348141;
      20790: inst = 32'd203451216;
      20791: inst = 32'd136314880;
      20792: inst = 32'd268468224;
      20793: inst = 32'd201348142;
      20794: inst = 32'd203451216;
      20795: inst = 32'd136314880;
      20796: inst = 32'd268468224;
      20797: inst = 32'd201348143;
      20798: inst = 32'd203451216;
      20799: inst = 32'd136314880;
      20800: inst = 32'd268468224;
      20801: inst = 32'd201348144;
      20802: inst = 32'd203451248;
      20803: inst = 32'd136314880;
      20804: inst = 32'd268468224;
      20805: inst = 32'd201348145;
      20806: inst = 32'd203449168;
      20807: inst = 32'd136314880;
      20808: inst = 32'd268468224;
      20809: inst = 32'd201348146;
      20810: inst = 32'd203449136;
      20811: inst = 32'd136314880;
      20812: inst = 32'd268468224;
      20813: inst = 32'd201348147;
      20814: inst = 32'd203451249;
      20815: inst = 32'd136314880;
      20816: inst = 32'd268468224;
      20817: inst = 32'd201348148;
      20818: inst = 32'd203451249;
      20819: inst = 32'd136314880;
      20820: inst = 32'd268468224;
      20821: inst = 32'd201348149;
      20822: inst = 32'd203451249;
      20823: inst = 32'd136314880;
      20824: inst = 32'd268468224;
      20825: inst = 32'd201348150;
      20826: inst = 32'd203451281;
      20827: inst = 32'd136314880;
      20828: inst = 32'd268468224;
      20829: inst = 32'd201348151;
      20830: inst = 32'd203451248;
      20831: inst = 32'd136314880;
      20832: inst = 32'd268468224;
      20833: inst = 32'd201348152;
      20834: inst = 32'd203449134;
      20835: inst = 32'd136314880;
      20836: inst = 32'd268468224;
      20837: inst = 32'd201348153;
      20838: inst = 32'd203455537;
      20839: inst = 32'd136314880;
      20840: inst = 32'd268468224;
      20841: inst = 32'd201348154;
      20842: inst = 32'd203457617;
      20843: inst = 32'd136314880;
      20844: inst = 32'd268468224;
      20845: inst = 32'd201348155;
      20846: inst = 32'd203459730;
      20847: inst = 32'd136314880;
      20848: inst = 32'd268468224;
      20849: inst = 32'd201348156;
      20850: inst = 32'd203451213;
      20851: inst = 32'd136314880;
      20852: inst = 32'd268468224;
      20853: inst = 32'd201348157;
      20854: inst = 32'd203442794;
      20855: inst = 32'd136314880;
      20856: inst = 32'd268468224;
      20857: inst = 32'd201348158;
      20858: inst = 32'd203442794;
      20859: inst = 32'd136314880;
      20860: inst = 32'd268468224;
      20861: inst = 32'd201348159;
      20862: inst = 32'd203444843;
      20863: inst = 32'd136314880;
      20864: inst = 32'd268468224;
      20865: inst = 32'd201348160;
      20866: inst = 32'd203457552;
      20867: inst = 32'd136314880;
      20868: inst = 32'd268468224;
      20869: inst = 32'd201348161;
      20870: inst = 32'd203455407;
      20871: inst = 32'd136314880;
      20872: inst = 32'd268468224;
      20873: inst = 32'd201348162;
      20874: inst = 32'd203444842;
      20875: inst = 32'd136314880;
      20876: inst = 32'd268468224;
      20877: inst = 32'd201348163;
      20878: inst = 32'd203442761;
      20879: inst = 32'd136314880;
      20880: inst = 32'd268468224;
      20881: inst = 32'd201348164;
      20882: inst = 32'd203451213;
      20883: inst = 32'd136314880;
      20884: inst = 32'd268468224;
      20885: inst = 32'd201348165;
      20886: inst = 32'd203459665;
      20887: inst = 32'd136314880;
      20888: inst = 32'd268468224;
      20889: inst = 32'd201348166;
      20890: inst = 32'd203459729;
      20891: inst = 32'd136314880;
      20892: inst = 32'd268468224;
      20893: inst = 32'd201348167;
      20894: inst = 32'd203457649;
      20895: inst = 32'd136314880;
      20896: inst = 32'd268468224;
      20897: inst = 32'd201348168;
      20898: inst = 32'd203453424;
      20899: inst = 32'd136314880;
      20900: inst = 32'd268468224;
      20901: inst = 32'd201348169;
      20902: inst = 32'd203442891;
      20903: inst = 32'd136314880;
      20904: inst = 32'd268468224;
      20905: inst = 32'd201348170;
      20906: inst = 32'd203449199;
      20907: inst = 32'd136314880;
      20908: inst = 32'd268468224;
      20909: inst = 32'd201348171;
      20910: inst = 32'd203449232;
      20911: inst = 32'd136314880;
      20912: inst = 32'd268468224;
      20913: inst = 32'd201348172;
      20914: inst = 32'd203449168;
      20915: inst = 32'd136314880;
      20916: inst = 32'd268468224;
      20917: inst = 32'd201348173;
      20918: inst = 32'd203449168;
      20919: inst = 32'd136314880;
      20920: inst = 32'd268468224;
      20921: inst = 32'd201348174;
      20922: inst = 32'd203449201;
      20923: inst = 32'd136314880;
      20924: inst = 32'd268468224;
      20925: inst = 32'd201348175;
      20926: inst = 32'd203451282;
      20927: inst = 32'd136314880;
      20928: inst = 32'd268468224;
      20929: inst = 32'd201348176;
      20930: inst = 32'd203449201;
      20931: inst = 32'd136314880;
      20932: inst = 32'd268468224;
      20933: inst = 32'd201348177;
      20934: inst = 32'd203449201;
      20935: inst = 32'd136314880;
      20936: inst = 32'd268468224;
      20937: inst = 32'd201348178;
      20938: inst = 32'd203447120;
      20939: inst = 32'd136314880;
      20940: inst = 32'd268468224;
      20941: inst = 32'd201348179;
      20942: inst = 32'd203447087;
      20943: inst = 32'd136314880;
      20944: inst = 32'd268468224;
      20945: inst = 32'd201348180;
      20946: inst = 32'd203449199;
      20947: inst = 32'd136314880;
      20948: inst = 32'd268468224;
      20949: inst = 32'd201348181;
      20950: inst = 32'd203449166;
      20951: inst = 32'd136314880;
      20952: inst = 32'd268468224;
      20953: inst = 32'd201348182;
      20954: inst = 32'd203442859;
      20955: inst = 32'd136314880;
      20956: inst = 32'd268468224;
      20957: inst = 32'd201348183;
      20958: inst = 32'd203453391;
      20959: inst = 32'd136314880;
      20960: inst = 32'd268468224;
      20961: inst = 32'd201348184;
      20962: inst = 32'd203457649;
      20963: inst = 32'd136314880;
      20964: inst = 32'd268468224;
      20965: inst = 32'd201348185;
      20966: inst = 32'd203459729;
      20967: inst = 32'd136314880;
      20968: inst = 32'd268468224;
      20969: inst = 32'd201348186;
      20970: inst = 32'd203459665;
      20971: inst = 32'd136314880;
      20972: inst = 32'd268468224;
      20973: inst = 32'd201348187;
      20974: inst = 32'd203451213;
      20975: inst = 32'd136314880;
      20976: inst = 32'd268468224;
      20977: inst = 32'd201348188;
      20978: inst = 32'd203442761;
      20979: inst = 32'd136314880;
      20980: inst = 32'd268468224;
      20981: inst = 32'd201348189;
      20982: inst = 32'd203444842;
      20983: inst = 32'd136314880;
      20984: inst = 32'd268468224;
      20985: inst = 32'd201348190;
      20986: inst = 32'd203455407;
      20987: inst = 32'd136314880;
      20988: inst = 32'd268468224;
      20989: inst = 32'd201348191;
      20990: inst = 32'd203457552;
      20991: inst = 32'd136314880;
      20992: inst = 32'd268468224;
      20993: inst = 32'd201348192;
      20994: inst = 32'd203442826;
      20995: inst = 32'd136314880;
      20996: inst = 32'd268468224;
      20997: inst = 32'd201348193;
      20998: inst = 32'd203442793;
      20999: inst = 32'd136314880;
      21000: inst = 32'd268468224;
      21001: inst = 32'd201348194;
      21002: inst = 32'd203442826;
      21003: inst = 32'd136314880;
      21004: inst = 32'd268468224;
      21005: inst = 32'd201348195;
      21006: inst = 32'd203451213;
      21007: inst = 32'd136314880;
      21008: inst = 32'd268468224;
      21009: inst = 32'd201348196;
      21010: inst = 32'd203461745;
      21011: inst = 32'd136314880;
      21012: inst = 32'd268468224;
      21013: inst = 32'd201348197;
      21014: inst = 32'd203459697;
      21015: inst = 32'd136314880;
      21016: inst = 32'd268468224;
      21017: inst = 32'd201348198;
      21018: inst = 32'd203457552;
      21019: inst = 32'd136314880;
      21020: inst = 32'd268468224;
      21021: inst = 32'd201348199;
      21022: inst = 32'd203449166;
      21023: inst = 32'd136314880;
      21024: inst = 32'd268468224;
      21025: inst = 32'd201348200;
      21026: inst = 32'd203447087;
      21027: inst = 32'd136314880;
      21028: inst = 32'd268468224;
      21029: inst = 32'd201348201;
      21030: inst = 32'd203449201;
      21031: inst = 32'd136314880;
      21032: inst = 32'd268468224;
      21033: inst = 32'd201348202;
      21034: inst = 32'd203447120;
      21035: inst = 32'd136314880;
      21036: inst = 32'd268468224;
      21037: inst = 32'd201348203;
      21038: inst = 32'd203447153;
      21039: inst = 32'd136314880;
      21040: inst = 32'd268468224;
      21041: inst = 32'd201348204;
      21042: inst = 32'd203449202;
      21043: inst = 32'd136314880;
      21044: inst = 32'd268468224;
      21045: inst = 32'd201348205;
      21046: inst = 32'd203449234;
      21047: inst = 32'd136314880;
      21048: inst = 32'd268468224;
      21049: inst = 32'd201348206;
      21050: inst = 32'd203451282;
      21051: inst = 32'd136314880;
      21052: inst = 32'd268468224;
      21053: inst = 32'd201348207;
      21054: inst = 32'd203449169;
      21055: inst = 32'd136314880;
      21056: inst = 32'd268468224;
      21057: inst = 32'd201348208;
      21058: inst = 32'd203451216;
      21059: inst = 32'd136314880;
      21060: inst = 32'd268468224;
      21061: inst = 32'd201348209;
      21062: inst = 32'd203451216;
      21063: inst = 32'd136314880;
      21064: inst = 32'd268468224;
      21065: inst = 32'd201348210;
      21066: inst = 32'd203451216;
      21067: inst = 32'd136314880;
      21068: inst = 32'd268468224;
      21069: inst = 32'd201348211;
      21070: inst = 32'd203451216;
      21071: inst = 32'd136314880;
      21072: inst = 32'd268468224;
      21073: inst = 32'd201348212;
      21074: inst = 32'd203451216;
      21075: inst = 32'd136314880;
      21076: inst = 32'd268468224;
      21077: inst = 32'd201348213;
      21078: inst = 32'd203451216;
      21079: inst = 32'd136314880;
      21080: inst = 32'd268468224;
      21081: inst = 32'd201348214;
      21082: inst = 32'd203451216;
      21083: inst = 32'd136314880;
      21084: inst = 32'd268468224;
      21085: inst = 32'd201348215;
      21086: inst = 32'd203451216;
      21087: inst = 32'd136314880;
      21088: inst = 32'd268468224;
      21089: inst = 32'd201348216;
      21090: inst = 32'd203451248;
      21091: inst = 32'd136314880;
      21092: inst = 32'd268468224;
      21093: inst = 32'd201348217;
      21094: inst = 32'd203451215;
      21095: inst = 32'd136314880;
      21096: inst = 32'd268468224;
      21097: inst = 32'd201348218;
      21098: inst = 32'd203451248;
      21099: inst = 32'd136314880;
      21100: inst = 32'd268468224;
      21101: inst = 32'd201348219;
      21102: inst = 32'd203451248;
      21103: inst = 32'd136314880;
      21104: inst = 32'd268468224;
      21105: inst = 32'd201348220;
      21106: inst = 32'd203449167;
      21107: inst = 32'd136314880;
      21108: inst = 32'd268468224;
      21109: inst = 32'd201348221;
      21110: inst = 32'd203451216;
      21111: inst = 32'd136314880;
      21112: inst = 32'd268468224;
      21113: inst = 32'd201348222;
      21114: inst = 32'd203451248;
      21115: inst = 32'd136314880;
      21116: inst = 32'd268468224;
      21117: inst = 32'd201348223;
      21118: inst = 32'd203451215;
      21119: inst = 32'd136314880;
      21120: inst = 32'd268468224;
      21121: inst = 32'd201348224;
      21122: inst = 32'd203451248;
      21123: inst = 32'd136314880;
      21124: inst = 32'd268468224;
      21125: inst = 32'd201348225;
      21126: inst = 32'd203451216;
      21127: inst = 32'd136314880;
      21128: inst = 32'd268468224;
      21129: inst = 32'd201348226;
      21130: inst = 32'd203451248;
      21131: inst = 32'd136314880;
      21132: inst = 32'd268468224;
      21133: inst = 32'd201348227;
      21134: inst = 32'd203449135;
      21135: inst = 32'd136314880;
      21136: inst = 32'd268468224;
      21137: inst = 32'd201348228;
      21138: inst = 32'd203451216;
      21139: inst = 32'd136314880;
      21140: inst = 32'd268468224;
      21141: inst = 32'd201348229;
      21142: inst = 32'd203451281;
      21143: inst = 32'd136314880;
      21144: inst = 32'd268468224;
      21145: inst = 32'd201348230;
      21146: inst = 32'd203449167;
      21147: inst = 32'd136314880;
      21148: inst = 32'd268468224;
      21149: inst = 32'd201348231;
      21150: inst = 32'd203451248;
      21151: inst = 32'd136314880;
      21152: inst = 32'd268468224;
      21153: inst = 32'd201348232;
      21154: inst = 32'd203451216;
      21155: inst = 32'd136314880;
      21156: inst = 32'd268468224;
      21157: inst = 32'd201348233;
      21158: inst = 32'd203451248;
      21159: inst = 32'd136314880;
      21160: inst = 32'd268468224;
      21161: inst = 32'd201348234;
      21162: inst = 32'd203449135;
      21163: inst = 32'd136314880;
      21164: inst = 32'd268468224;
      21165: inst = 32'd201348235;
      21166: inst = 32'd203451281;
      21167: inst = 32'd136314880;
      21168: inst = 32'd268468224;
      21169: inst = 32'd201348236;
      21170: inst = 32'd203451216;
      21171: inst = 32'd136314880;
      21172: inst = 32'd268468224;
      21173: inst = 32'd201348237;
      21174: inst = 32'd203451216;
      21175: inst = 32'd136314880;
      21176: inst = 32'd268468224;
      21177: inst = 32'd201348238;
      21178: inst = 32'd203451216;
      21179: inst = 32'd136314880;
      21180: inst = 32'd268468224;
      21181: inst = 32'd201348239;
      21182: inst = 32'd203451248;
      21183: inst = 32'd136314880;
      21184: inst = 32'd268468224;
      21185: inst = 32'd201348240;
      21186: inst = 32'd203451215;
      21187: inst = 32'd136314880;
      21188: inst = 32'd268468224;
      21189: inst = 32'd201348241;
      21190: inst = 32'd203451216;
      21191: inst = 32'd136314880;
      21192: inst = 32'd268468224;
      21193: inst = 32'd201348242;
      21194: inst = 32'd203449168;
      21195: inst = 32'd136314880;
      21196: inst = 32'd268468224;
      21197: inst = 32'd201348243;
      21198: inst = 32'd203451281;
      21199: inst = 32'd136314880;
      21200: inst = 32'd268468224;
      21201: inst = 32'd201348244;
      21202: inst = 32'd203449136;
      21203: inst = 32'd136314880;
      21204: inst = 32'd268468224;
      21205: inst = 32'd201348245;
      21206: inst = 32'd203449169;
      21207: inst = 32'd136314880;
      21208: inst = 32'd268468224;
      21209: inst = 32'd201348246;
      21210: inst = 32'd203451248;
      21211: inst = 32'd136314880;
      21212: inst = 32'd268468224;
      21213: inst = 32'd201348247;
      21214: inst = 32'd203449199;
      21215: inst = 32'd136314880;
      21216: inst = 32'd268468224;
      21217: inst = 32'd201348248;
      21218: inst = 32'd203453425;
      21219: inst = 32'd136314880;
      21220: inst = 32'd268468224;
      21221: inst = 32'd201348249;
      21222: inst = 32'd203457650;
      21223: inst = 32'd136314880;
      21224: inst = 32'd268468224;
      21225: inst = 32'd201348250;
      21226: inst = 32'd203457650;
      21227: inst = 32'd136314880;
      21228: inst = 32'd268468224;
      21229: inst = 32'd201348251;
      21230: inst = 32'd203455504;
      21231: inst = 32'd136314880;
      21232: inst = 32'd268468224;
      21233: inst = 32'd201348252;
      21234: inst = 32'd203442761;
      21235: inst = 32'd136314880;
      21236: inst = 32'd268468224;
      21237: inst = 32'd201348253;
      21238: inst = 32'd203442793;
      21239: inst = 32'd136314880;
      21240: inst = 32'd268468224;
      21241: inst = 32'd201348254;
      21242: inst = 32'd203446955;
      21243: inst = 32'd136314880;
      21244: inst = 32'd268468224;
      21245: inst = 32'd201348255;
      21246: inst = 32'd203446955;
      21247: inst = 32'd136314880;
      21248: inst = 32'd268468224;
      21249: inst = 32'd201348256;
      21250: inst = 32'd203444842;
      21251: inst = 32'd136314880;
      21252: inst = 32'd268468224;
      21253: inst = 32'd201348257;
      21254: inst = 32'd203444842;
      21255: inst = 32'd136314880;
      21256: inst = 32'd268468224;
      21257: inst = 32'd201348258;
      21258: inst = 32'd203442761;
      21259: inst = 32'd136314880;
      21260: inst = 32'd268468224;
      21261: inst = 32'd201348259;
      21262: inst = 32'd203444874;
      21263: inst = 32'd136314880;
      21264: inst = 32'd268468224;
      21265: inst = 32'd201348260;
      21266: inst = 32'd203457552;
      21267: inst = 32'd136314880;
      21268: inst = 32'd268468224;
      21269: inst = 32'd201348261;
      21270: inst = 32'd203459665;
      21271: inst = 32'd136314880;
      21272: inst = 32'd268468224;
      21273: inst = 32'd201348262;
      21274: inst = 32'd203461778;
      21275: inst = 32'd136314880;
      21276: inst = 32'd268468224;
      21277: inst = 32'd201348263;
      21278: inst = 32'd203459697;
      21279: inst = 32'd136314880;
      21280: inst = 32'd268468224;
      21281: inst = 32'd201348264;
      21282: inst = 32'd203451278;
      21283: inst = 32'd136314880;
      21284: inst = 32'd268468224;
      21285: inst = 32'd201348265;
      21286: inst = 32'd203442826;
      21287: inst = 32'd136314880;
      21288: inst = 32'd268468224;
      21289: inst = 32'd201348266;
      21290: inst = 32'd203449166;
      21291: inst = 32'd136314880;
      21292: inst = 32'd268468224;
      21293: inst = 32'd201348267;
      21294: inst = 32'd203451280;
      21295: inst = 32'd136314880;
      21296: inst = 32'd268468224;
      21297: inst = 32'd201348268;
      21298: inst = 32'd203449200;
      21299: inst = 32'd136314880;
      21300: inst = 32'd268468224;
      21301: inst = 32'd201348269;
      21302: inst = 32'd203449201;
      21303: inst = 32'd136314880;
      21304: inst = 32'd268468224;
      21305: inst = 32'd201348270;
      21306: inst = 32'd203449201;
      21307: inst = 32'd136314880;
      21308: inst = 32'd268468224;
      21309: inst = 32'd201348271;
      21310: inst = 32'd203447089;
      21311: inst = 32'd136314880;
      21312: inst = 32'd268468224;
      21313: inst = 32'd201348272;
      21314: inst = 32'd203447089;
      21315: inst = 32'd136314880;
      21316: inst = 32'd268468224;
      21317: inst = 32'd201348273;
      21318: inst = 32'd203449201;
      21319: inst = 32'd136314880;
      21320: inst = 32'd268468224;
      21321: inst = 32'd201348274;
      21322: inst = 32'd203449201;
      21323: inst = 32'd136314880;
      21324: inst = 32'd268468224;
      21325: inst = 32'd201348275;
      21326: inst = 32'd203449200;
      21327: inst = 32'd136314880;
      21328: inst = 32'd268468224;
      21329: inst = 32'd201348276;
      21330: inst = 32'd203451312;
      21331: inst = 32'd136314880;
      21332: inst = 32'd268468224;
      21333: inst = 32'd201348277;
      21334: inst = 32'd203449198;
      21335: inst = 32'd136314880;
      21336: inst = 32'd268468224;
      21337: inst = 32'd201348278;
      21338: inst = 32'd203442827;
      21339: inst = 32'd136314880;
      21340: inst = 32'd268468224;
      21341: inst = 32'd201348279;
      21342: inst = 32'd203451278;
      21343: inst = 32'd136314880;
      21344: inst = 32'd268468224;
      21345: inst = 32'd201348280;
      21346: inst = 32'd203459697;
      21347: inst = 32'd136314880;
      21348: inst = 32'd268468224;
      21349: inst = 32'd201348281;
      21350: inst = 32'd203461778;
      21351: inst = 32'd136314880;
      21352: inst = 32'd268468224;
      21353: inst = 32'd201348282;
      21354: inst = 32'd203459665;
      21355: inst = 32'd136314880;
      21356: inst = 32'd268468224;
      21357: inst = 32'd201348283;
      21358: inst = 32'd203457552;
      21359: inst = 32'd136314880;
      21360: inst = 32'd268468224;
      21361: inst = 32'd201348284;
      21362: inst = 32'd203444874;
      21363: inst = 32'd136314880;
      21364: inst = 32'd268468224;
      21365: inst = 32'd201348285;
      21366: inst = 32'd203442761;
      21367: inst = 32'd136314880;
      21368: inst = 32'd268468224;
      21369: inst = 32'd201348286;
      21370: inst = 32'd203444842;
      21371: inst = 32'd136314880;
      21372: inst = 32'd268468224;
      21373: inst = 32'd201348287;
      21374: inst = 32'd203444842;
      21375: inst = 32'd136314880;
      21376: inst = 32'd268468224;
      21377: inst = 32'd201348288;
      21378: inst = 32'd203444938;
      21379: inst = 32'd136314880;
      21380: inst = 32'd268468224;
      21381: inst = 32'd201348289;
      21382: inst = 32'd203442858;
      21383: inst = 32'd136314880;
      21384: inst = 32'd268468224;
      21385: inst = 32'd201348290;
      21386: inst = 32'd203442825;
      21387: inst = 32'd136314880;
      21388: inst = 32'd268468224;
      21389: inst = 32'd201348291;
      21390: inst = 32'd203442760;
      21391: inst = 32'd136314880;
      21392: inst = 32'd268468224;
      21393: inst = 32'd201348292;
      21394: inst = 32'd203455503;
      21395: inst = 32'd136314880;
      21396: inst = 32'd268468224;
      21397: inst = 32'd201348293;
      21398: inst = 32'd203459729;
      21399: inst = 32'd136314880;
      21400: inst = 32'd268468224;
      21401: inst = 32'd201348294;
      21402: inst = 32'd203457617;
      21403: inst = 32'd136314880;
      21404: inst = 32'd268468224;
      21405: inst = 32'd201348295;
      21406: inst = 32'd203455504;
      21407: inst = 32'd136314880;
      21408: inst = 32'd268468224;
      21409: inst = 32'd201348296;
      21410: inst = 32'd203451279;
      21411: inst = 32'd136314880;
      21412: inst = 32'd268468224;
      21413: inst = 32'd201348297;
      21414: inst = 32'd203451280;
      21415: inst = 32'd136314880;
      21416: inst = 32'd268468224;
      21417: inst = 32'd201348298;
      21418: inst = 32'd203447120;
      21419: inst = 32'd136314880;
      21420: inst = 32'd268468224;
      21421: inst = 32'd201348299;
      21422: inst = 32'd203449233;
      21423: inst = 32'd136314880;
      21424: inst = 32'd268468224;
      21425: inst = 32'd201348300;
      21426: inst = 32'd203449201;
      21427: inst = 32'd136314880;
      21428: inst = 32'd268468224;
      21429: inst = 32'd201348301;
      21430: inst = 32'd203447088;
      21431: inst = 32'd136314880;
      21432: inst = 32'd268468224;
      21433: inst = 32'd201348302;
      21434: inst = 32'd203451281;
      21435: inst = 32'd136314880;
      21436: inst = 32'd268468224;
      21437: inst = 32'd201348303;
      21438: inst = 32'd203451249;
      21439: inst = 32'd136314880;
      21440: inst = 32'd268468224;
      21441: inst = 32'd201348304;
      21442: inst = 32'd203453262;
      21443: inst = 32'd136314880;
      21444: inst = 32'd268468224;
      21445: inst = 32'd201348305;
      21446: inst = 32'd203453262;
      21447: inst = 32'd136314880;
      21448: inst = 32'd268468224;
      21449: inst = 32'd201348306;
      21450: inst = 32'd203453262;
      21451: inst = 32'd136314880;
      21452: inst = 32'd268468224;
      21453: inst = 32'd201348307;
      21454: inst = 32'd203453262;
      21455: inst = 32'd136314880;
      21456: inst = 32'd268468224;
      21457: inst = 32'd201348308;
      21458: inst = 32'd203453262;
      21459: inst = 32'd136314880;
      21460: inst = 32'd268468224;
      21461: inst = 32'd201348309;
      21462: inst = 32'd203453262;
      21463: inst = 32'd136314880;
      21464: inst = 32'd268468224;
      21465: inst = 32'd201348310;
      21466: inst = 32'd203453262;
      21467: inst = 32'd136314880;
      21468: inst = 32'd268468224;
      21469: inst = 32'd201348311;
      21470: inst = 32'd203453262;
      21471: inst = 32'd136314880;
      21472: inst = 32'd268468224;
      21473: inst = 32'd201348312;
      21474: inst = 32'd203453262;
      21475: inst = 32'd136314880;
      21476: inst = 32'd268468224;
      21477: inst = 32'd201348313;
      21478: inst = 32'd203453262;
      21479: inst = 32'd136314880;
      21480: inst = 32'd268468224;
      21481: inst = 32'd201348314;
      21482: inst = 32'd203453262;
      21483: inst = 32'd136314880;
      21484: inst = 32'd268468224;
      21485: inst = 32'd201348315;
      21486: inst = 32'd203453262;
      21487: inst = 32'd136314880;
      21488: inst = 32'd268468224;
      21489: inst = 32'd201348316;
      21490: inst = 32'd203453230;
      21491: inst = 32'd136314880;
      21492: inst = 32'd268468224;
      21493: inst = 32'd201348317;
      21494: inst = 32'd203453262;
      21495: inst = 32'd136314880;
      21496: inst = 32'd268468224;
      21497: inst = 32'd201348318;
      21498: inst = 32'd203453295;
      21499: inst = 32'd136314880;
      21500: inst = 32'd268468224;
      21501: inst = 32'd201348319;
      21502: inst = 32'd203453262;
      21503: inst = 32'd136314880;
      21504: inst = 32'd268468224;
      21505: inst = 32'd201348320;
      21506: inst = 32'd203449200;
      21507: inst = 32'd136314880;
      21508: inst = 32'd268468224;
      21509: inst = 32'd201348321;
      21510: inst = 32'd203449200;
      21511: inst = 32'd136314880;
      21512: inst = 32'd268468224;
      21513: inst = 32'd201348322;
      21514: inst = 32'd203449200;
      21515: inst = 32'd136314880;
      21516: inst = 32'd268468224;
      21517: inst = 32'd201348323;
      21518: inst = 32'd203449200;
      21519: inst = 32'd136314880;
      21520: inst = 32'd268468224;
      21521: inst = 32'd201348324;
      21522: inst = 32'd203449200;
      21523: inst = 32'd136314880;
      21524: inst = 32'd268468224;
      21525: inst = 32'd201348325;
      21526: inst = 32'd203449200;
      21527: inst = 32'd136314880;
      21528: inst = 32'd268468224;
      21529: inst = 32'd201348326;
      21530: inst = 32'd203449200;
      21531: inst = 32'd136314880;
      21532: inst = 32'd268468224;
      21533: inst = 32'd201348327;
      21534: inst = 32'd203449200;
      21535: inst = 32'd136314880;
      21536: inst = 32'd268468224;
      21537: inst = 32'd201348328;
      21538: inst = 32'd203449200;
      21539: inst = 32'd136314880;
      21540: inst = 32'd268468224;
      21541: inst = 32'd201348329;
      21542: inst = 32'd203449200;
      21543: inst = 32'd136314880;
      21544: inst = 32'd268468224;
      21545: inst = 32'd201348330;
      21546: inst = 32'd203449200;
      21547: inst = 32'd136314880;
      21548: inst = 32'd268468224;
      21549: inst = 32'd201348331;
      21550: inst = 32'd203449200;
      21551: inst = 32'd136314880;
      21552: inst = 32'd268468224;
      21553: inst = 32'd201348332;
      21554: inst = 32'd203449200;
      21555: inst = 32'd136314880;
      21556: inst = 32'd268468224;
      21557: inst = 32'd201348333;
      21558: inst = 32'd203449200;
      21559: inst = 32'd136314880;
      21560: inst = 32'd268468224;
      21561: inst = 32'd201348334;
      21562: inst = 32'd203449200;
      21563: inst = 32'd136314880;
      21564: inst = 32'd268468224;
      21565: inst = 32'd201348335;
      21566: inst = 32'd203449200;
      21567: inst = 32'd136314880;
      21568: inst = 32'd268468224;
      21569: inst = 32'd201348336;
      21570: inst = 32'd203451215;
      21571: inst = 32'd136314880;
      21572: inst = 32'd268468224;
      21573: inst = 32'd201348337;
      21574: inst = 32'd203451216;
      21575: inst = 32'd136314880;
      21576: inst = 32'd268468224;
      21577: inst = 32'd201348338;
      21578: inst = 32'd203451248;
      21579: inst = 32'd136314880;
      21580: inst = 32'd268468224;
      21581: inst = 32'd201348339;
      21582: inst = 32'd203451216;
      21583: inst = 32'd136314880;
      21584: inst = 32'd268468224;
      21585: inst = 32'd201348340;
      21586: inst = 32'd203451216;
      21587: inst = 32'd136314880;
      21588: inst = 32'd268468224;
      21589: inst = 32'd201348341;
      21590: inst = 32'd203449168;
      21591: inst = 32'd136314880;
      21592: inst = 32'd268468224;
      21593: inst = 32'd201348342;
      21594: inst = 32'd203451280;
      21595: inst = 32'd136314880;
      21596: inst = 32'd268468224;
      21597: inst = 32'd201348343;
      21598: inst = 32'd203451312;
      21599: inst = 32'd136314880;
      21600: inst = 32'd268468224;
      21601: inst = 32'd201348344;
      21602: inst = 32'd203457651;
      21603: inst = 32'd136314880;
      21604: inst = 32'd268468224;
      21605: inst = 32'd201348345;
      21606: inst = 32'd203459698;
      21607: inst = 32'd136314880;
      21608: inst = 32'd268468224;
      21609: inst = 32'd201348346;
      21610: inst = 32'd203459697;
      21611: inst = 32'd136314880;
      21612: inst = 32'd268468224;
      21613: inst = 32'd201348347;
      21614: inst = 32'd203444939;
      21615: inst = 32'd136314880;
      21616: inst = 32'd268468224;
      21617: inst = 32'd201348348;
      21618: inst = 32'd203444874;
      21619: inst = 32'd136314880;
      21620: inst = 32'd268468224;
      21621: inst = 32'd201348349;
      21622: inst = 32'd203442793;
      21623: inst = 32'd136314880;
      21624: inst = 32'd268468224;
      21625: inst = 32'd201348350;
      21626: inst = 32'd203444841;
      21627: inst = 32'd136314880;
      21628: inst = 32'd268468224;
      21629: inst = 32'd201348351;
      21630: inst = 32'd203455374;
      21631: inst = 32'd136314880;
      21632: inst = 32'd268468224;
      21633: inst = 32'd201348352;
      21634: inst = 32'd203459666;
      21635: inst = 32'd136314880;
      21636: inst = 32'd268468224;
      21637: inst = 32'd201348353;
      21638: inst = 32'd203455472;
      21639: inst = 32'd136314880;
      21640: inst = 32'd268468224;
      21641: inst = 32'd201348354;
      21642: inst = 32'd203442761;
      21643: inst = 32'd136314880;
      21644: inst = 32'd268468224;
      21645: inst = 32'd201348355;
      21646: inst = 32'd203446987;
      21647: inst = 32'd136314880;
      21648: inst = 32'd268468224;
      21649: inst = 32'd201348356;
      21650: inst = 32'd203459697;
      21651: inst = 32'd136314880;
      21652: inst = 32'd268468224;
      21653: inst = 32'd201348357;
      21654: inst = 32'd203459697;
      21655: inst = 32'd136314880;
      21656: inst = 32'd268468224;
      21657: inst = 32'd201348358;
      21658: inst = 32'd203459729;
      21659: inst = 32'd136314880;
      21660: inst = 32'd268468224;
      21661: inst = 32'd201348359;
      21662: inst = 32'd203459665;
      21663: inst = 32'd136314880;
      21664: inst = 32'd268468224;
      21665: inst = 32'd201348360;
      21666: inst = 32'd203449132;
      21667: inst = 32'd136314880;
      21668: inst = 32'd268468224;
      21669: inst = 32'd201348361;
      21670: inst = 32'd203444907;
      21671: inst = 32'd136314880;
      21672: inst = 32'd268468224;
      21673: inst = 32'd201348362;
      21674: inst = 32'd203451247;
      21675: inst = 32'd136314880;
      21676: inst = 32'd268468224;
      21677: inst = 32'd201348363;
      21678: inst = 32'd203451247;
      21679: inst = 32'd136314880;
      21680: inst = 32'd268468224;
      21681: inst = 32'd201348364;
      21682: inst = 32'd203451248;
      21683: inst = 32'd136314880;
      21684: inst = 32'd268468224;
      21685: inst = 32'd201348365;
      21686: inst = 32'd203449168;
      21687: inst = 32'd136314880;
      21688: inst = 32'd268468224;
      21689: inst = 32'd201348366;
      21690: inst = 32'd203449169;
      21691: inst = 32'd136314880;
      21692: inst = 32'd268468224;
      21693: inst = 32'd201348367;
      21694: inst = 32'd203451217;
      21695: inst = 32'd136314880;
      21696: inst = 32'd268468224;
      21697: inst = 32'd201348368;
      21698: inst = 32'd203451217;
      21699: inst = 32'd136314880;
      21700: inst = 32'd268468224;
      21701: inst = 32'd201348369;
      21702: inst = 32'd203449169;
      21703: inst = 32'd136314880;
      21704: inst = 32'd268468224;
      21705: inst = 32'd201348370;
      21706: inst = 32'd203449168;
      21707: inst = 32'd136314880;
      21708: inst = 32'd268468224;
      21709: inst = 32'd201348371;
      21710: inst = 32'd203451248;
      21711: inst = 32'd136314880;
      21712: inst = 32'd268468224;
      21713: inst = 32'd201348372;
      21714: inst = 32'd203451247;
      21715: inst = 32'd136314880;
      21716: inst = 32'd268468224;
      21717: inst = 32'd201348373;
      21718: inst = 32'd203451247;
      21719: inst = 32'd136314880;
      21720: inst = 32'd268468224;
      21721: inst = 32'd201348374;
      21722: inst = 32'd203444907;
      21723: inst = 32'd136314880;
      21724: inst = 32'd268468224;
      21725: inst = 32'd201348375;
      21726: inst = 32'd203449132;
      21727: inst = 32'd136314880;
      21728: inst = 32'd268468224;
      21729: inst = 32'd201348376;
      21730: inst = 32'd203459697;
      21731: inst = 32'd136314880;
      21732: inst = 32'd268468224;
      21733: inst = 32'd201348377;
      21734: inst = 32'd203459697;
      21735: inst = 32'd136314880;
      21736: inst = 32'd268468224;
      21737: inst = 32'd201348378;
      21738: inst = 32'd203459665;
      21739: inst = 32'd136314880;
      21740: inst = 32'd268468224;
      21741: inst = 32'd201348379;
      21742: inst = 32'd203459697;
      21743: inst = 32'd136314880;
      21744: inst = 32'd268468224;
      21745: inst = 32'd201348380;
      21746: inst = 32'd203447019;
      21747: inst = 32'd136314880;
      21748: inst = 32'd268468224;
      21749: inst = 32'd201348381;
      21750: inst = 32'd203442729;
      21751: inst = 32'd136314880;
      21752: inst = 32'd268468224;
      21753: inst = 32'd201348382;
      21754: inst = 32'd203455440;
      21755: inst = 32'd136314880;
      21756: inst = 32'd268468224;
      21757: inst = 32'd201348383;
      21758: inst = 32'd203459666;
      21759: inst = 32'd136314880;
      21760: inst = 32'd268468224;
      21761: inst = 32'd201348384;
      21762: inst = 32'd203451309;
      21763: inst = 32'd136314880;
      21764: inst = 32'd268468224;
      21765: inst = 32'd201348385;
      21766: inst = 32'd203442825;
      21767: inst = 32'd136314880;
      21768: inst = 32'd268468224;
      21769: inst = 32'd201348386;
      21770: inst = 32'd203442825;
      21771: inst = 32'd136314880;
      21772: inst = 32'd268468224;
      21773: inst = 32'd201348387;
      21774: inst = 32'd203444873;
      21775: inst = 32'd136314880;
      21776: inst = 32'd268468224;
      21777: inst = 32'd201348388;
      21778: inst = 32'd203444938;
      21779: inst = 32'd136314880;
      21780: inst = 32'd268468224;
      21781: inst = 32'd201348389;
      21782: inst = 32'd203459664;
      21783: inst = 32'd136314880;
      21784: inst = 32'd268468224;
      21785: inst = 32'd201348390;
      21786: inst = 32'd203459697;
      21787: inst = 32'd136314880;
      21788: inst = 32'd268468224;
      21789: inst = 32'd201348391;
      21790: inst = 32'd203459697;
      21791: inst = 32'd136314880;
      21792: inst = 32'd268468224;
      21793: inst = 32'd201348392;
      21794: inst = 32'd203453359;
      21795: inst = 32'd136314880;
      21796: inst = 32'd268468224;
      21797: inst = 32'd201348393;
      21798: inst = 32'd203451279;
      21799: inst = 32'd136314880;
      21800: inst = 32'd268468224;
      21801: inst = 32'd201348394;
      21802: inst = 32'd203449199;
      21803: inst = 32'd136314880;
      21804: inst = 32'd268468224;
      21805: inst = 32'd201348395;
      21806: inst = 32'd203449199;
      21807: inst = 32'd136314880;
      21808: inst = 32'd268468224;
      21809: inst = 32'd201348396;
      21810: inst = 32'd203449200;
      21811: inst = 32'd136314880;
      21812: inst = 32'd268468224;
      21813: inst = 32'd201348397;
      21814: inst = 32'd203451248;
      21815: inst = 32'd136314880;
      21816: inst = 32'd268468224;
      21817: inst = 32'd201348398;
      21818: inst = 32'd203451248;
      21819: inst = 32'd136314880;
      21820: inst = 32'd268468224;
      21821: inst = 32'd201348399;
      21822: inst = 32'd203451216;
      21823: inst = 32'd136314880;
      21824: inst = 32'd268468224;
      21825: inst = 32'd201348400;
      21826: inst = 32'd203453263;
      21827: inst = 32'd136314880;
      21828: inst = 32'd268468224;
      21829: inst = 32'd201348401;
      21830: inst = 32'd203453263;
      21831: inst = 32'd136314880;
      21832: inst = 32'd268468224;
      21833: inst = 32'd201348402;
      21834: inst = 32'd203453263;
      21835: inst = 32'd136314880;
      21836: inst = 32'd268468224;
      21837: inst = 32'd201348403;
      21838: inst = 32'd203453263;
      21839: inst = 32'd136314880;
      21840: inst = 32'd268468224;
      21841: inst = 32'd201348404;
      21842: inst = 32'd203453263;
      21843: inst = 32'd136314880;
      21844: inst = 32'd268468224;
      21845: inst = 32'd201348405;
      21846: inst = 32'd203453263;
      21847: inst = 32'd136314880;
      21848: inst = 32'd268468224;
      21849: inst = 32'd201348406;
      21850: inst = 32'd203453263;
      21851: inst = 32'd136314880;
      21852: inst = 32'd268468224;
      21853: inst = 32'd201348407;
      21854: inst = 32'd203453263;
      21855: inst = 32'd136314880;
      21856: inst = 32'd268468224;
      21857: inst = 32'd201348408;
      21858: inst = 32'd203453263;
      21859: inst = 32'd136314880;
      21860: inst = 32'd268468224;
      21861: inst = 32'd201348409;
      21862: inst = 32'd203453263;
      21863: inst = 32'd136314880;
      21864: inst = 32'd268468224;
      21865: inst = 32'd201348410;
      21866: inst = 32'd203453263;
      21867: inst = 32'd136314880;
      21868: inst = 32'd268468224;
      21869: inst = 32'd201348411;
      21870: inst = 32'd203453263;
      21871: inst = 32'd136314880;
      21872: inst = 32'd268468224;
      21873: inst = 32'd201348412;
      21874: inst = 32'd203453263;
      21875: inst = 32'd136314880;
      21876: inst = 32'd268468224;
      21877: inst = 32'd201348413;
      21878: inst = 32'd203453263;
      21879: inst = 32'd136314880;
      21880: inst = 32'd268468224;
      21881: inst = 32'd201348414;
      21882: inst = 32'd203453263;
      21883: inst = 32'd136314880;
      21884: inst = 32'd268468224;
      21885: inst = 32'd201348415;
      21886: inst = 32'd203453263;
      21887: inst = 32'd136314880;
      21888: inst = 32'd268468224;
      21889: inst = 32'd201348416;
      21890: inst = 32'd203449200;
      21891: inst = 32'd136314880;
      21892: inst = 32'd268468224;
      21893: inst = 32'd201348417;
      21894: inst = 32'd203449200;
      21895: inst = 32'd136314880;
      21896: inst = 32'd268468224;
      21897: inst = 32'd201348418;
      21898: inst = 32'd203449200;
      21899: inst = 32'd136314880;
      21900: inst = 32'd268468224;
      21901: inst = 32'd201348419;
      21902: inst = 32'd203449200;
      21903: inst = 32'd136314880;
      21904: inst = 32'd268468224;
      21905: inst = 32'd201348420;
      21906: inst = 32'd203449200;
      21907: inst = 32'd136314880;
      21908: inst = 32'd268468224;
      21909: inst = 32'd201348421;
      21910: inst = 32'd203449200;
      21911: inst = 32'd136314880;
      21912: inst = 32'd268468224;
      21913: inst = 32'd201348422;
      21914: inst = 32'd203449200;
      21915: inst = 32'd136314880;
      21916: inst = 32'd268468224;
      21917: inst = 32'd201348423;
      21918: inst = 32'd203449200;
      21919: inst = 32'd136314880;
      21920: inst = 32'd268468224;
      21921: inst = 32'd201348424;
      21922: inst = 32'd203449200;
      21923: inst = 32'd136314880;
      21924: inst = 32'd268468224;
      21925: inst = 32'd201348425;
      21926: inst = 32'd203449200;
      21927: inst = 32'd136314880;
      21928: inst = 32'd268468224;
      21929: inst = 32'd201348426;
      21930: inst = 32'd203449200;
      21931: inst = 32'd136314880;
      21932: inst = 32'd268468224;
      21933: inst = 32'd201348427;
      21934: inst = 32'd203449200;
      21935: inst = 32'd136314880;
      21936: inst = 32'd268468224;
      21937: inst = 32'd201348428;
      21938: inst = 32'd203449200;
      21939: inst = 32'd136314880;
      21940: inst = 32'd268468224;
      21941: inst = 32'd201348429;
      21942: inst = 32'd203449200;
      21943: inst = 32'd136314880;
      21944: inst = 32'd268468224;
      21945: inst = 32'd201348430;
      21946: inst = 32'd203449200;
      21947: inst = 32'd136314880;
      21948: inst = 32'd268468224;
      21949: inst = 32'd201348431;
      21950: inst = 32'd203449200;
      21951: inst = 32'd136314880;
      21952: inst = 32'd268468224;
      21953: inst = 32'd201348432;
      21954: inst = 32'd203451215;
      21955: inst = 32'd136314880;
      21956: inst = 32'd268468224;
      21957: inst = 32'd201348433;
      21958: inst = 32'd203451183;
      21959: inst = 32'd136314880;
      21960: inst = 32'd268468224;
      21961: inst = 32'd201348434;
      21962: inst = 32'd203451215;
      21963: inst = 32'd136314880;
      21964: inst = 32'd268468224;
      21965: inst = 32'd201348435;
      21966: inst = 32'd203453296;
      21967: inst = 32'd136314880;
      21968: inst = 32'd268468224;
      21969: inst = 32'd201348436;
      21970: inst = 32'd203451247;
      21971: inst = 32'd136314880;
      21972: inst = 32'd268468224;
      21973: inst = 32'd201348437;
      21974: inst = 32'd203449167;
      21975: inst = 32'd136314880;
      21976: inst = 32'd268468224;
      21977: inst = 32'd201348438;
      21978: inst = 32'd203453360;
      21979: inst = 32'd136314880;
      21980: inst = 32'd268468224;
      21981: inst = 32'd201348439;
      21982: inst = 32'd203457586;
      21983: inst = 32'd136314880;
      21984: inst = 32'd268468224;
      21985: inst = 32'd201348440;
      21986: inst = 32'd203459730;
      21987: inst = 32'd136314880;
      21988: inst = 32'd268468224;
      21989: inst = 32'd201348441;
      21990: inst = 32'd203459698;
      21991: inst = 32'd136314880;
      21992: inst = 32'd268468224;
      21993: inst = 32'd201348442;
      21994: inst = 32'd203451213;
      21995: inst = 32'd136314880;
      21996: inst = 32'd268468224;
      21997: inst = 32'd201348443;
      21998: inst = 32'd203442793;
      21999: inst = 32'd136314880;
      22000: inst = 32'd268468224;
      22001: inst = 32'd201348444;
      22002: inst = 32'd203442760;
      22003: inst = 32'd136314880;
      22004: inst = 32'd268468224;
      22005: inst = 32'd201348445;
      22006: inst = 32'd203444873;
      22007: inst = 32'd136314880;
      22008: inst = 32'd268468224;
      22009: inst = 32'd201348446;
      22010: inst = 32'd203444841;
      22011: inst = 32'd136314880;
      22012: inst = 32'd268468224;
      22013: inst = 32'd201348447;
      22014: inst = 32'd203459664;
      22015: inst = 32'd136314880;
      22016: inst = 32'd268468224;
      22017: inst = 32'd201348448;
      22018: inst = 32'd203459666;
      22019: inst = 32'd136314880;
      22020: inst = 32'd268468224;
      22021: inst = 32'd201348449;
      22022: inst = 32'd203455472;
      22023: inst = 32'd136314880;
      22024: inst = 32'd268468224;
      22025: inst = 32'd201348450;
      22026: inst = 32'd203442761;
      22027: inst = 32'd136314880;
      22028: inst = 32'd268468224;
      22029: inst = 32'd201348451;
      22030: inst = 32'd203451213;
      22031: inst = 32'd136314880;
      22032: inst = 32'd268468224;
      22033: inst = 32'd201348452;
      22034: inst = 32'd203459665;
      22035: inst = 32'd136314880;
      22036: inst = 32'd268468224;
      22037: inst = 32'd201348453;
      22038: inst = 32'd203461778;
      22039: inst = 32'd136314880;
      22040: inst = 32'd268468224;
      22041: inst = 32'd201348454;
      22042: inst = 32'd203459697;
      22043: inst = 32'd136314880;
      22044: inst = 32'd268468224;
      22045: inst = 32'd201348455;
      22046: inst = 32'd203459697;
      22047: inst = 32'd136314880;
      22048: inst = 32'd268468224;
      22049: inst = 32'd201348456;
      22050: inst = 32'd203447020;
      22051: inst = 32'd136314880;
      22052: inst = 32'd268468224;
      22053: inst = 32'd201348457;
      22054: inst = 32'd203444874;
      22055: inst = 32'd136314880;
      22056: inst = 32'd268468224;
      22057: inst = 32'd201348458;
      22058: inst = 32'd203451214;
      22059: inst = 32'd136314880;
      22060: inst = 32'd268468224;
      22061: inst = 32'd201348459;
      22062: inst = 32'd203451215;
      22063: inst = 32'd136314880;
      22064: inst = 32'd268468224;
      22065: inst = 32'd201348460;
      22066: inst = 32'd203451248;
      22067: inst = 32'd136314880;
      22068: inst = 32'd268468224;
      22069: inst = 32'd201348461;
      22070: inst = 32'd203451216;
      22071: inst = 32'd136314880;
      22072: inst = 32'd268468224;
      22073: inst = 32'd201348462;
      22074: inst = 32'd203451216;
      22075: inst = 32'd136314880;
      22076: inst = 32'd268468224;
      22077: inst = 32'd201348463;
      22078: inst = 32'd203451217;
      22079: inst = 32'd136314880;
      22080: inst = 32'd268468224;
      22081: inst = 32'd201348464;
      22082: inst = 32'd203451217;
      22083: inst = 32'd136314880;
      22084: inst = 32'd268468224;
      22085: inst = 32'd201348465;
      22086: inst = 32'd203451216;
      22087: inst = 32'd136314880;
      22088: inst = 32'd268468224;
      22089: inst = 32'd201348466;
      22090: inst = 32'd203451216;
      22091: inst = 32'd136314880;
      22092: inst = 32'd268468224;
      22093: inst = 32'd201348467;
      22094: inst = 32'd203451248;
      22095: inst = 32'd136314880;
      22096: inst = 32'd268468224;
      22097: inst = 32'd201348468;
      22098: inst = 32'd203451215;
      22099: inst = 32'd136314880;
      22100: inst = 32'd268468224;
      22101: inst = 32'd201348469;
      22102: inst = 32'd203451214;
      22103: inst = 32'd136314880;
      22104: inst = 32'd268468224;
      22105: inst = 32'd201348470;
      22106: inst = 32'd203444874;
      22107: inst = 32'd136314880;
      22108: inst = 32'd268468224;
      22109: inst = 32'd201348471;
      22110: inst = 32'd203447020;
      22111: inst = 32'd136314880;
      22112: inst = 32'd268468224;
      22113: inst = 32'd201348472;
      22114: inst = 32'd203459697;
      22115: inst = 32'd136314880;
      22116: inst = 32'd268468224;
      22117: inst = 32'd201348473;
      22118: inst = 32'd203459697;
      22119: inst = 32'd136314880;
      22120: inst = 32'd268468224;
      22121: inst = 32'd201348474;
      22122: inst = 32'd203461778;
      22123: inst = 32'd136314880;
      22124: inst = 32'd268468224;
      22125: inst = 32'd201348475;
      22126: inst = 32'd203459665;
      22127: inst = 32'd136314880;
      22128: inst = 32'd268468224;
      22129: inst = 32'd201348476;
      22130: inst = 32'd203451245;
      22131: inst = 32'd136314880;
      22132: inst = 32'd268468224;
      22133: inst = 32'd201348477;
      22134: inst = 32'd203440713;
      22135: inst = 32'd136314880;
      22136: inst = 32'd268468224;
      22137: inst = 32'd201348478;
      22138: inst = 32'd203455472;
      22139: inst = 32'd136314880;
      22140: inst = 32'd268468224;
      22141: inst = 32'd201348479;
      22142: inst = 32'd203459698;
      22143: inst = 32'd136314880;
      22144: inst = 32'd268468224;
      22145: inst = 32'd201348480;
      22146: inst = 32'd203457649;
      22147: inst = 32'd136314880;
      22148: inst = 32'd268468224;
      22149: inst = 32'd201348481;
      22150: inst = 32'd203442825;
      22151: inst = 32'd136314880;
      22152: inst = 32'd268468224;
      22153: inst = 32'd201348482;
      22154: inst = 32'd203442825;
      22155: inst = 32'd136314880;
      22156: inst = 32'd268468224;
      22157: inst = 32'd201348483;
      22158: inst = 32'd203442760;
      22159: inst = 32'd136314880;
      22160: inst = 32'd268468224;
      22161: inst = 32'd201348484;
      22162: inst = 32'd203442793;
      22163: inst = 32'd136314880;
      22164: inst = 32'd268468224;
      22165: inst = 32'd201348485;
      22166: inst = 32'd203451212;
      22167: inst = 32'd136314880;
      22168: inst = 32'd268468224;
      22169: inst = 32'd201348486;
      22170: inst = 32'd203459697;
      22171: inst = 32'd136314880;
      22172: inst = 32'd268468224;
      22173: inst = 32'd201348487;
      22174: inst = 32'd203459698;
      22175: inst = 32'd136314880;
      22176: inst = 32'd268468224;
      22177: inst = 32'd201348488;
      22178: inst = 32'd203457585;
      22179: inst = 32'd136314880;
      22180: inst = 32'd268468224;
      22181: inst = 32'd201348489;
      22182: inst = 32'd203453359;
      22183: inst = 32'd136314880;
      22184: inst = 32'd268468224;
      22185: inst = 32'd201348490;
      22186: inst = 32'd203451214;
      22187: inst = 32'd136314880;
      22188: inst = 32'd268468224;
      22189: inst = 32'd201348491;
      22190: inst = 32'd203451247;
      22191: inst = 32'd136314880;
      22192: inst = 32'd268468224;
      22193: inst = 32'd201348492;
      22194: inst = 32'd203451248;
      22195: inst = 32'd136314880;
      22196: inst = 32'd268468224;
      22197: inst = 32'd201348493;
      22198: inst = 32'd203451215;
      22199: inst = 32'd136314880;
      22200: inst = 32'd268468224;
      22201: inst = 32'd201348494;
      22202: inst = 32'd203451183;
      22203: inst = 32'd136314880;
      22204: inst = 32'd268468224;
      22205: inst = 32'd201348495;
      22206: inst = 32'd203451216;
      22207: inst = 32'd136314880;
      22208: inst = 32'd268468224;
      22209: inst = 32'd201348496;
      22210: inst = 32'd203449168;
      22211: inst = 32'd136314880;
      22212: inst = 32'd268468224;
      22213: inst = 32'd201348497;
      22214: inst = 32'd203449168;
      22215: inst = 32'd136314880;
      22216: inst = 32'd268468224;
      22217: inst = 32'd201348498;
      22218: inst = 32'd203449168;
      22219: inst = 32'd136314880;
      22220: inst = 32'd268468224;
      22221: inst = 32'd201348499;
      22222: inst = 32'd203449168;
      22223: inst = 32'd136314880;
      22224: inst = 32'd268468224;
      22225: inst = 32'd201348500;
      22226: inst = 32'd203449168;
      22227: inst = 32'd136314880;
      22228: inst = 32'd268468224;
      22229: inst = 32'd201348501;
      22230: inst = 32'd203449168;
      22231: inst = 32'd136314880;
      22232: inst = 32'd268468224;
      22233: inst = 32'd201348502;
      22234: inst = 32'd203449168;
      22235: inst = 32'd136314880;
      22236: inst = 32'd268468224;
      22237: inst = 32'd201348503;
      22238: inst = 32'd203449168;
      22239: inst = 32'd136314880;
      22240: inst = 32'd268468224;
      22241: inst = 32'd201348504;
      22242: inst = 32'd203449168;
      22243: inst = 32'd136314880;
      22244: inst = 32'd268468224;
      22245: inst = 32'd201348505;
      22246: inst = 32'd203449168;
      22247: inst = 32'd136314880;
      22248: inst = 32'd268468224;
      22249: inst = 32'd201348506;
      22250: inst = 32'd203449168;
      22251: inst = 32'd136314880;
      22252: inst = 32'd268468224;
      22253: inst = 32'd201348507;
      22254: inst = 32'd203449168;
      22255: inst = 32'd136314880;
      22256: inst = 32'd268468224;
      22257: inst = 32'd201348508;
      22258: inst = 32'd203449168;
      22259: inst = 32'd136314880;
      22260: inst = 32'd268468224;
      22261: inst = 32'd201348509;
      22262: inst = 32'd203449168;
      22263: inst = 32'd136314880;
      22264: inst = 32'd268468224;
      22265: inst = 32'd201348510;
      22266: inst = 32'd203449168;
      22267: inst = 32'd136314880;
      22268: inst = 32'd268468224;
      22269: inst = 32'd201348511;
      22270: inst = 32'd203449168;
      22271: inst = 32'd136314880;
      22272: inst = 32'd268468224;
      22273: inst = 32'd201348512;
      22274: inst = 32'd203451247;
      22275: inst = 32'd136314880;
      22276: inst = 32'd268468224;
      22277: inst = 32'd201348513;
      22278: inst = 32'd203451247;
      22279: inst = 32'd136314880;
      22280: inst = 32'd268468224;
      22281: inst = 32'd201348514;
      22282: inst = 32'd203451247;
      22283: inst = 32'd136314880;
      22284: inst = 32'd268468224;
      22285: inst = 32'd201348515;
      22286: inst = 32'd203451247;
      22287: inst = 32'd136314880;
      22288: inst = 32'd268468224;
      22289: inst = 32'd201348516;
      22290: inst = 32'd203451247;
      22291: inst = 32'd136314880;
      22292: inst = 32'd268468224;
      22293: inst = 32'd201348517;
      22294: inst = 32'd203451247;
      22295: inst = 32'd136314880;
      22296: inst = 32'd268468224;
      22297: inst = 32'd201348518;
      22298: inst = 32'd203451247;
      22299: inst = 32'd136314880;
      22300: inst = 32'd268468224;
      22301: inst = 32'd201348519;
      22302: inst = 32'd203451247;
      22303: inst = 32'd136314880;
      22304: inst = 32'd268468224;
      22305: inst = 32'd201348520;
      22306: inst = 32'd203451247;
      22307: inst = 32'd136314880;
      22308: inst = 32'd268468224;
      22309: inst = 32'd201348521;
      22310: inst = 32'd203451247;
      22311: inst = 32'd136314880;
      22312: inst = 32'd268468224;
      22313: inst = 32'd201348522;
      22314: inst = 32'd203451247;
      22315: inst = 32'd136314880;
      22316: inst = 32'd268468224;
      22317: inst = 32'd201348523;
      22318: inst = 32'd203451247;
      22319: inst = 32'd136314880;
      22320: inst = 32'd268468224;
      22321: inst = 32'd201348524;
      22322: inst = 32'd203451247;
      22323: inst = 32'd136314880;
      22324: inst = 32'd268468224;
      22325: inst = 32'd201348525;
      22326: inst = 32'd203451247;
      22327: inst = 32'd136314880;
      22328: inst = 32'd268468224;
      22329: inst = 32'd201348526;
      22330: inst = 32'd203451247;
      22331: inst = 32'd136314880;
      22332: inst = 32'd268468224;
      22333: inst = 32'd201348527;
      22334: inst = 32'd203451247;
      22335: inst = 32'd136314880;
      22336: inst = 32'd268468224;
      22337: inst = 32'd201348528;
      22338: inst = 32'd203453263;
      22339: inst = 32'd136314880;
      22340: inst = 32'd268468224;
      22341: inst = 32'd201348529;
      22342: inst = 32'd203451215;
      22343: inst = 32'd136314880;
      22344: inst = 32'd268468224;
      22345: inst = 32'd201348530;
      22346: inst = 32'd203451215;
      22347: inst = 32'd136314880;
      22348: inst = 32'd268468224;
      22349: inst = 32'd201348531;
      22350: inst = 32'd203451247;
      22351: inst = 32'd136314880;
      22352: inst = 32'd268468224;
      22353: inst = 32'd201348532;
      22354: inst = 32'd203451247;
      22355: inst = 32'd136314880;
      22356: inst = 32'd268468224;
      22357: inst = 32'd201348533;
      22358: inst = 32'd203451279;
      22359: inst = 32'd136314880;
      22360: inst = 32'd268468224;
      22361: inst = 32'd201348534;
      22362: inst = 32'd203455504;
      22363: inst = 32'd136314880;
      22364: inst = 32'd268468224;
      22365: inst = 32'd201348535;
      22366: inst = 32'd203459730;
      22367: inst = 32'd136314880;
      22368: inst = 32'd268468224;
      22369: inst = 32'd201348536;
      22370: inst = 32'd203457617;
      22371: inst = 32'd136314880;
      22372: inst = 32'd268468224;
      22373: inst = 32'd201348537;
      22374: inst = 32'd203453358;
      22375: inst = 32'd136314880;
      22376: inst = 32'd268468224;
      22377: inst = 32'd201348538;
      22378: inst = 32'd203444873;
      22379: inst = 32'd136314880;
      22380: inst = 32'd268468224;
      22381: inst = 32'd201348539;
      22382: inst = 32'd203442793;
      22383: inst = 32'd136314880;
      22384: inst = 32'd268468224;
      22385: inst = 32'd201348540;
      22386: inst = 32'd203442793;
      22387: inst = 32'd136314880;
      22388: inst = 32'd268468224;
      22389: inst = 32'd201348541;
      22390: inst = 32'd203444873;
      22391: inst = 32'd136314880;
      22392: inst = 32'd268468224;
      22393: inst = 32'd201348542;
      22394: inst = 32'd203449066;
      22395: inst = 32'd136314880;
      22396: inst = 32'd268468224;
      22397: inst = 32'd201348543;
      22398: inst = 32'd203461712;
      22399: inst = 32'd136314880;
      22400: inst = 32'd268468224;
      22401: inst = 32'd201348544;
      22402: inst = 32'd203459698;
      22403: inst = 32'd136314880;
      22404: inst = 32'd268468224;
      22405: inst = 32'd201348545;
      22406: inst = 32'd203455440;
      22407: inst = 32'd136314880;
      22408: inst = 32'd268468224;
      22409: inst = 32'd201348546;
      22410: inst = 32'd203442794;
      22411: inst = 32'd136314880;
      22412: inst = 32'd268468224;
      22413: inst = 32'd201348547;
      22414: inst = 32'd203455504;
      22415: inst = 32'd136314880;
      22416: inst = 32'd268468224;
      22417: inst = 32'd201348548;
      22418: inst = 32'd203459665;
      22419: inst = 32'd136314880;
      22420: inst = 32'd268468224;
      22421: inst = 32'd201348549;
      22422: inst = 32'd203461778;
      22423: inst = 32'd136314880;
      22424: inst = 32'd268468224;
      22425: inst = 32'd201348550;
      22426: inst = 32'd203459665;
      22427: inst = 32'd136314880;
      22428: inst = 32'd268468224;
      22429: inst = 32'd201348551;
      22430: inst = 32'd203459697;
      22431: inst = 32'd136314880;
      22432: inst = 32'd268468224;
      22433: inst = 32'd201348552;
      22434: inst = 32'd203446955;
      22435: inst = 32'd136314880;
      22436: inst = 32'd268468224;
      22437: inst = 32'd201348553;
      22438: inst = 32'd203444842;
      22439: inst = 32'd136314880;
      22440: inst = 32'd268468224;
      22441: inst = 32'd201348554;
      22442: inst = 32'd203451214;
      22443: inst = 32'd136314880;
      22444: inst = 32'd268468224;
      22445: inst = 32'd201348555;
      22446: inst = 32'd203451214;
      22447: inst = 32'd136314880;
      22448: inst = 32'd268468224;
      22449: inst = 32'd201348556;
      22450: inst = 32'd203451215;
      22451: inst = 32'd136314880;
      22452: inst = 32'd268468224;
      22453: inst = 32'd201348557;
      22454: inst = 32'd203451215;
      22455: inst = 32'd136314880;
      22456: inst = 32'd268468224;
      22457: inst = 32'd201348558;
      22458: inst = 32'd203451216;
      22459: inst = 32'd136314880;
      22460: inst = 32'd268468224;
      22461: inst = 32'd201348559;
      22462: inst = 32'd203451248;
      22463: inst = 32'd136314880;
      22464: inst = 32'd268468224;
      22465: inst = 32'd201348560;
      22466: inst = 32'd203451248;
      22467: inst = 32'd136314880;
      22468: inst = 32'd268468224;
      22469: inst = 32'd201348561;
      22470: inst = 32'd203451216;
      22471: inst = 32'd136314880;
      22472: inst = 32'd268468224;
      22473: inst = 32'd201348562;
      22474: inst = 32'd203451215;
      22475: inst = 32'd136314880;
      22476: inst = 32'd268468224;
      22477: inst = 32'd201348563;
      22478: inst = 32'd203451215;
      22479: inst = 32'd136314880;
      22480: inst = 32'd268468224;
      22481: inst = 32'd201348564;
      22482: inst = 32'd203451214;
      22483: inst = 32'd136314880;
      22484: inst = 32'd268468224;
      22485: inst = 32'd201348565;
      22486: inst = 32'd203451214;
      22487: inst = 32'd136314880;
      22488: inst = 32'd268468224;
      22489: inst = 32'd201348566;
      22490: inst = 32'd203444842;
      22491: inst = 32'd136314880;
      22492: inst = 32'd268468224;
      22493: inst = 32'd201348567;
      22494: inst = 32'd203446955;
      22495: inst = 32'd136314880;
      22496: inst = 32'd268468224;
      22497: inst = 32'd201348568;
      22498: inst = 32'd203459697;
      22499: inst = 32'd136314880;
      22500: inst = 32'd268468224;
      22501: inst = 32'd201348569;
      22502: inst = 32'd203459697;
      22503: inst = 32'd136314880;
      22504: inst = 32'd268468224;
      22505: inst = 32'd201348570;
      22506: inst = 32'd203461778;
      22507: inst = 32'd136314880;
      22508: inst = 32'd268468224;
      22509: inst = 32'd201348571;
      22510: inst = 32'd203457585;
      22511: inst = 32'd136314880;
      22512: inst = 32'd268468224;
      22513: inst = 32'd201348572;
      22514: inst = 32'd203455472;
      22515: inst = 32'd136314880;
      22516: inst = 32'd268468224;
      22517: inst = 32'd201348573;
      22518: inst = 32'd203442794;
      22519: inst = 32'd136314880;
      22520: inst = 32'd268468224;
      22521: inst = 32'd201348574;
      22522: inst = 32'd203455440;
      22523: inst = 32'd136314880;
      22524: inst = 32'd268468224;
      22525: inst = 32'd201348575;
      22526: inst = 32'd203459698;
      22527: inst = 32'd136314880;
      22528: inst = 32'd268468224;
      22529: inst = 32'd201348576;
      22530: inst = 32'd203459697;
      22531: inst = 32'd136314880;
      22532: inst = 32'd268468224;
      22533: inst = 32'd201348577;
      22534: inst = 32'd203447020;
      22535: inst = 32'd136314880;
      22536: inst = 32'd268468224;
      22537: inst = 32'd201348578;
      22538: inst = 32'd203444874;
      22539: inst = 32'd136314880;
      22540: inst = 32'd268468224;
      22541: inst = 32'd201348579;
      22542: inst = 32'd203442793;
      22543: inst = 32'd136314880;
      22544: inst = 32'd268468224;
      22545: inst = 32'd201348580;
      22546: inst = 32'd203442794;
      22547: inst = 32'd136314880;
      22548: inst = 32'd268468224;
      22549: inst = 32'd201348581;
      22550: inst = 32'd203444874;
      22551: inst = 32'd136314880;
      22552: inst = 32'd268468224;
      22553: inst = 32'd201348582;
      22554: inst = 32'd203453358;
      22555: inst = 32'd136314880;
      22556: inst = 32'd268468224;
      22557: inst = 32'd201348583;
      22558: inst = 32'd203459633;
      22559: inst = 32'd136314880;
      22560: inst = 32'd268468224;
      22561: inst = 32'd201348584;
      22562: inst = 32'd203461746;
      22563: inst = 32'd136314880;
      22564: inst = 32'd268468224;
      22565: inst = 32'd201348585;
      22566: inst = 32'd203457520;
      22567: inst = 32'd136314880;
      22568: inst = 32'd268468224;
      22569: inst = 32'd201348586;
      22570: inst = 32'd203453295;
      22571: inst = 32'd136314880;
      22572: inst = 32'd268468224;
      22573: inst = 32'd201348587;
      22574: inst = 32'd203451215;
      22575: inst = 32'd136314880;
      22576: inst = 32'd268468224;
      22577: inst = 32'd201348588;
      22578: inst = 32'd203451215;
      22579: inst = 32'd136314880;
      22580: inst = 32'd268468224;
      22581: inst = 32'd201348589;
      22582: inst = 32'd203451215;
      22583: inst = 32'd136314880;
      22584: inst = 32'd268468224;
      22585: inst = 32'd201348590;
      22586: inst = 32'd203451183;
      22587: inst = 32'd136314880;
      22588: inst = 32'd268468224;
      22589: inst = 32'd201348591;
      22590: inst = 32'd203451216;
      22591: inst = 32'd136314880;
      22592: inst = 32'd268468224;
      22593: inst = 32'd201348592;
      22594: inst = 32'd203449200;
      22595: inst = 32'd136314880;
      22596: inst = 32'd268468224;
      22597: inst = 32'd201348593;
      22598: inst = 32'd203449200;
      22599: inst = 32'd136314880;
      22600: inst = 32'd268468224;
      22601: inst = 32'd201348594;
      22602: inst = 32'd203449200;
      22603: inst = 32'd136314880;
      22604: inst = 32'd268468224;
      22605: inst = 32'd201348595;
      22606: inst = 32'd203449200;
      22607: inst = 32'd136314880;
      22608: inst = 32'd268468224;
      22609: inst = 32'd201348596;
      22610: inst = 32'd203449200;
      22611: inst = 32'd136314880;
      22612: inst = 32'd268468224;
      22613: inst = 32'd201348597;
      22614: inst = 32'd203449200;
      22615: inst = 32'd136314880;
      22616: inst = 32'd268468224;
      22617: inst = 32'd201348598;
      22618: inst = 32'd203449200;
      22619: inst = 32'd136314880;
      22620: inst = 32'd268468224;
      22621: inst = 32'd201348599;
      22622: inst = 32'd203449200;
      22623: inst = 32'd136314880;
      22624: inst = 32'd268468224;
      22625: inst = 32'd201348600;
      22626: inst = 32'd203449200;
      22627: inst = 32'd136314880;
      22628: inst = 32'd268468224;
      22629: inst = 32'd201348601;
      22630: inst = 32'd203449200;
      22631: inst = 32'd136314880;
      22632: inst = 32'd268468224;
      22633: inst = 32'd201348602;
      22634: inst = 32'd203449200;
      22635: inst = 32'd136314880;
      22636: inst = 32'd268468224;
      22637: inst = 32'd201348603;
      22638: inst = 32'd203449200;
      22639: inst = 32'd136314880;
      22640: inst = 32'd268468224;
      22641: inst = 32'd201348604;
      22642: inst = 32'd203449200;
      22643: inst = 32'd136314880;
      22644: inst = 32'd268468224;
      22645: inst = 32'd201348605;
      22646: inst = 32'd203449200;
      22647: inst = 32'd136314880;
      22648: inst = 32'd268468224;
      22649: inst = 32'd201348606;
      22650: inst = 32'd203449200;
      22651: inst = 32'd136314880;
      22652: inst = 32'd268468224;
      22653: inst = 32'd201348607;
      22654: inst = 32'd203449200;
      22655: inst = 32'd136314880;
      22656: inst = 32'd268468224;
      22657: inst = 32'd201348608;
      22658: inst = 32'd203451247;
      22659: inst = 32'd136314880;
      22660: inst = 32'd268468224;
      22661: inst = 32'd201348609;
      22662: inst = 32'd203451247;
      22663: inst = 32'd136314880;
      22664: inst = 32'd268468224;
      22665: inst = 32'd201348610;
      22666: inst = 32'd203451247;
      22667: inst = 32'd136314880;
      22668: inst = 32'd268468224;
      22669: inst = 32'd201348611;
      22670: inst = 32'd203451247;
      22671: inst = 32'd136314880;
      22672: inst = 32'd268468224;
      22673: inst = 32'd201348612;
      22674: inst = 32'd203451247;
      22675: inst = 32'd136314880;
      22676: inst = 32'd268468224;
      22677: inst = 32'd201348613;
      22678: inst = 32'd203451247;
      22679: inst = 32'd136314880;
      22680: inst = 32'd268468224;
      22681: inst = 32'd201348614;
      22682: inst = 32'd203451247;
      22683: inst = 32'd136314880;
      22684: inst = 32'd268468224;
      22685: inst = 32'd201348615;
      22686: inst = 32'd203451247;
      22687: inst = 32'd136314880;
      22688: inst = 32'd268468224;
      22689: inst = 32'd201348616;
      22690: inst = 32'd203451247;
      22691: inst = 32'd136314880;
      22692: inst = 32'd268468224;
      22693: inst = 32'd201348617;
      22694: inst = 32'd203451247;
      22695: inst = 32'd136314880;
      22696: inst = 32'd268468224;
      22697: inst = 32'd201348618;
      22698: inst = 32'd203451247;
      22699: inst = 32'd136314880;
      22700: inst = 32'd268468224;
      22701: inst = 32'd201348619;
      22702: inst = 32'd203451247;
      22703: inst = 32'd136314880;
      22704: inst = 32'd268468224;
      22705: inst = 32'd201348620;
      22706: inst = 32'd203451247;
      22707: inst = 32'd136314880;
      22708: inst = 32'd268468224;
      22709: inst = 32'd201348621;
      22710: inst = 32'd203451247;
      22711: inst = 32'd136314880;
      22712: inst = 32'd268468224;
      22713: inst = 32'd201348622;
      22714: inst = 32'd203451247;
      22715: inst = 32'd136314880;
      22716: inst = 32'd268468224;
      22717: inst = 32'd201348623;
      22718: inst = 32'd203451247;
      22719: inst = 32'd136314880;
      22720: inst = 32'd268468224;
      22721: inst = 32'd201348624;
      22722: inst = 32'd203451215;
      22723: inst = 32'd136314880;
      22724: inst = 32'd268468224;
      22725: inst = 32'd201348625;
      22726: inst = 32'd203453296;
      22727: inst = 32'd136314880;
      22728: inst = 32'd268468224;
      22729: inst = 32'd201348626;
      22730: inst = 32'd203451215;
      22731: inst = 32'd136314880;
      22732: inst = 32'd268468224;
      22733: inst = 32'd201348627;
      22734: inst = 32'd203451182;
      22735: inst = 32'd136314880;
      22736: inst = 32'd268468224;
      22737: inst = 32'd201348628;
      22738: inst = 32'd203451246;
      22739: inst = 32'd136314880;
      22740: inst = 32'd268468224;
      22741: inst = 32'd201348629;
      22742: inst = 32'd203455504;
      22743: inst = 32'd136314880;
      22744: inst = 32'd268468224;
      22745: inst = 32'd201348630;
      22746: inst = 32'd203459698;
      22747: inst = 32'd136314880;
      22748: inst = 32'd268468224;
      22749: inst = 32'd201348631;
      22750: inst = 32'd203459697;
      22751: inst = 32'd136314880;
      22752: inst = 32'd268468224;
      22753: inst = 32'd201348632;
      22754: inst = 32'd203459697;
      22755: inst = 32'd136314880;
      22756: inst = 32'd268468224;
      22757: inst = 32'd201348633;
      22758: inst = 32'd203447019;
      22759: inst = 32'd136314880;
      22760: inst = 32'd268468224;
      22761: inst = 32'd201348634;
      22762: inst = 32'd203442761;
      22763: inst = 32'd136314880;
      22764: inst = 32'd268468224;
      22765: inst = 32'd201348635;
      22766: inst = 32'd203442793;
      22767: inst = 32'd136314880;
      22768: inst = 32'd268468224;
      22769: inst = 32'd201348636;
      22770: inst = 32'd203442760;
      22771: inst = 32'd136314880;
      22772: inst = 32'd268468224;
      22773: inst = 32'd201348637;
      22774: inst = 32'd203442760;
      22775: inst = 32'd136314880;
      22776: inst = 32'd268468224;
      22777: inst = 32'd201348638;
      22778: inst = 32'd203457551;
      22779: inst = 32'd136314880;
      22780: inst = 32'd268468224;
      22781: inst = 32'd201348639;
      22782: inst = 32'd203461777;
      22783: inst = 32'd136314880;
      22784: inst = 32'd268468224;
      22785: inst = 32'd201348640;
      22786: inst = 32'd203459730;
      22787: inst = 32'd136314880;
      22788: inst = 32'd268468224;
      22789: inst = 32'd201348641;
      22790: inst = 32'd203453359;
      22791: inst = 32'd136314880;
      22792: inst = 32'd268468224;
      22793: inst = 32'd201348642;
      22794: inst = 32'd203444939;
      22795: inst = 32'd136314880;
      22796: inst = 32'd268468224;
      22797: inst = 32'd201348643;
      22798: inst = 32'd203459698;
      22799: inst = 32'd136314880;
      22800: inst = 32'd268468224;
      22801: inst = 32'd201348644;
      22802: inst = 32'd203459665;
      22803: inst = 32'd136314880;
      22804: inst = 32'd268468224;
      22805: inst = 32'd201348645;
      22806: inst = 32'd203461778;
      22807: inst = 32'd136314880;
      22808: inst = 32'd268468224;
      22809: inst = 32'd201348646;
      22810: inst = 32'd203459665;
      22811: inst = 32'd136314880;
      22812: inst = 32'd268468224;
      22813: inst = 32'd201348647;
      22814: inst = 32'd203459665;
      22815: inst = 32'd136314880;
      22816: inst = 32'd268468224;
      22817: inst = 32'd201348648;
      22818: inst = 32'd203444875;
      22819: inst = 32'd136314880;
      22820: inst = 32'd268468224;
      22821: inst = 32'd201348649;
      22822: inst = 32'd203444842;
      22823: inst = 32'd136314880;
      22824: inst = 32'd268468224;
      22825: inst = 32'd201348650;
      22826: inst = 32'd203451214;
      22827: inst = 32'd136314880;
      22828: inst = 32'd268468224;
      22829: inst = 32'd201348651;
      22830: inst = 32'd203451215;
      22831: inst = 32'd136314880;
      22832: inst = 32'd268468224;
      22833: inst = 32'd201348652;
      22834: inst = 32'd203451215;
      22835: inst = 32'd136314880;
      22836: inst = 32'd268468224;
      22837: inst = 32'd201348653;
      22838: inst = 32'd203451215;
      22839: inst = 32'd136314880;
      22840: inst = 32'd268468224;
      22841: inst = 32'd201348654;
      22842: inst = 32'd203451215;
      22843: inst = 32'd136314880;
      22844: inst = 32'd268468224;
      22845: inst = 32'd201348655;
      22846: inst = 32'd203451248;
      22847: inst = 32'd136314880;
      22848: inst = 32'd268468224;
      22849: inst = 32'd201348656;
      22850: inst = 32'd203451248;
      22851: inst = 32'd136314880;
      22852: inst = 32'd268468224;
      22853: inst = 32'd201348657;
      22854: inst = 32'd203451215;
      22855: inst = 32'd136314880;
      22856: inst = 32'd268468224;
      22857: inst = 32'd201348658;
      22858: inst = 32'd203451215;
      22859: inst = 32'd136314880;
      22860: inst = 32'd268468224;
      22861: inst = 32'd201348659;
      22862: inst = 32'd203451215;
      22863: inst = 32'd136314880;
      22864: inst = 32'd268468224;
      22865: inst = 32'd201348660;
      22866: inst = 32'd203451215;
      22867: inst = 32'd136314880;
      22868: inst = 32'd268468224;
      22869: inst = 32'd201348661;
      22870: inst = 32'd203451214;
      22871: inst = 32'd136314880;
      22872: inst = 32'd268468224;
      22873: inst = 32'd201348662;
      22874: inst = 32'd203444842;
      22875: inst = 32'd136314880;
      22876: inst = 32'd268468224;
      22877: inst = 32'd201348663;
      22878: inst = 32'd203444875;
      22879: inst = 32'd136314880;
      22880: inst = 32'd268468224;
      22881: inst = 32'd201348664;
      22882: inst = 32'd203459633;
      22883: inst = 32'd136314880;
      22884: inst = 32'd268468224;
      22885: inst = 32'd201348665;
      22886: inst = 32'd203459697;
      22887: inst = 32'd136314880;
      22888: inst = 32'd268468224;
      22889: inst = 32'd201348666;
      22890: inst = 32'd203461778;
      22891: inst = 32'd136314880;
      22892: inst = 32'd268468224;
      22893: inst = 32'd201348667;
      22894: inst = 32'd203459665;
      22895: inst = 32'd136314880;
      22896: inst = 32'd268468224;
      22897: inst = 32'd201348668;
      22898: inst = 32'd203459665;
      22899: inst = 32'd136314880;
      22900: inst = 32'd268468224;
      22901: inst = 32'd201348669;
      22902: inst = 32'd203446987;
      22903: inst = 32'd136314880;
      22904: inst = 32'd268468224;
      22905: inst = 32'd201348670;
      22906: inst = 32'd203453391;
      22907: inst = 32'd136314880;
      22908: inst = 32'd268468224;
      22909: inst = 32'd201348671;
      22910: inst = 32'd203459698;
      22911: inst = 32'd136314880;
      22912: inst = 32'd268468224;
      22913: inst = 32'd201348672;
      22914: inst = 32'd203459730;
      22915: inst = 32'd136314880;
      22916: inst = 32'd268468224;
      22917: inst = 32'd201348673;
      22918: inst = 32'd203455504;
      22919: inst = 32'd136314880;
      22920: inst = 32'd268468224;
      22921: inst = 32'd201348674;
      22922: inst = 32'd203442761;
      22923: inst = 32'd136314880;
      22924: inst = 32'd268468224;
      22925: inst = 32'd201348675;
      22926: inst = 32'd203440681;
      22927: inst = 32'd136314880;
      22928: inst = 32'd268468224;
      22929: inst = 32'd201348676;
      22930: inst = 32'd203442794;
      22931: inst = 32'd136314880;
      22932: inst = 32'd268468224;
      22933: inst = 32'd201348677;
      22934: inst = 32'd203442762;
      22935: inst = 32'd136314880;
      22936: inst = 32'd268468224;
      22937: inst = 32'd201348678;
      22938: inst = 32'd203446988;
      22939: inst = 32'd136314880;
      22940: inst = 32'd268468224;
      22941: inst = 32'd201348679;
      22942: inst = 32'd203459666;
      22943: inst = 32'd136314880;
      22944: inst = 32'd268468224;
      22945: inst = 32'd201348680;
      22946: inst = 32'd203461746;
      22947: inst = 32'd136314880;
      22948: inst = 32'd268468224;
      22949: inst = 32'd201348681;
      22950: inst = 32'd203459634;
      22951: inst = 32'd136314880;
      22952: inst = 32'd268468224;
      22953: inst = 32'd201348682;
      22954: inst = 32'd203457488;
      22955: inst = 32'd136314880;
      22956: inst = 32'd268468224;
      22957: inst = 32'd201348683;
      22958: inst = 32'd203453263;
      22959: inst = 32'd136314880;
      22960: inst = 32'd268468224;
      22961: inst = 32'd201348684;
      22962: inst = 32'd203451182;
      22963: inst = 32'd136314880;
      22964: inst = 32'd268468224;
      22965: inst = 32'd201348685;
      22966: inst = 32'd203453264;
      22967: inst = 32'd136314880;
      22968: inst = 32'd268468224;
      22969: inst = 32'd201348686;
      22970: inst = 32'd203453296;
      22971: inst = 32'd136314880;
      22972: inst = 32'd268468224;
      22973: inst = 32'd201348687;
      22974: inst = 32'd203451215;
      22975: inst = 32'd136314880;
      22976: inst = 32'd268468224;
      22977: inst = 32'd201348688;
      22978: inst = 32'd203449168;
      22979: inst = 32'd136314880;
      22980: inst = 32'd268468224;
      22981: inst = 32'd201348689;
      22982: inst = 32'd203449168;
      22983: inst = 32'd136314880;
      22984: inst = 32'd268468224;
      22985: inst = 32'd201348690;
      22986: inst = 32'd203449168;
      22987: inst = 32'd136314880;
      22988: inst = 32'd268468224;
      22989: inst = 32'd201348691;
      22990: inst = 32'd203449168;
      22991: inst = 32'd136314880;
      22992: inst = 32'd268468224;
      22993: inst = 32'd201348692;
      22994: inst = 32'd203449168;
      22995: inst = 32'd136314880;
      22996: inst = 32'd268468224;
      22997: inst = 32'd201348693;
      22998: inst = 32'd203449168;
      22999: inst = 32'd136314880;
      23000: inst = 32'd268468224;
      23001: inst = 32'd201348694;
      23002: inst = 32'd203449168;
      23003: inst = 32'd136314880;
      23004: inst = 32'd268468224;
      23005: inst = 32'd201348695;
      23006: inst = 32'd203449168;
      23007: inst = 32'd136314880;
      23008: inst = 32'd268468224;
      23009: inst = 32'd201348696;
      23010: inst = 32'd203449168;
      23011: inst = 32'd136314880;
      23012: inst = 32'd268468224;
      23013: inst = 32'd201348697;
      23014: inst = 32'd203449168;
      23015: inst = 32'd136314880;
      23016: inst = 32'd268468224;
      23017: inst = 32'd201348698;
      23018: inst = 32'd203449168;
      23019: inst = 32'd136314880;
      23020: inst = 32'd268468224;
      23021: inst = 32'd201348699;
      23022: inst = 32'd203449168;
      23023: inst = 32'd136314880;
      23024: inst = 32'd268468224;
      23025: inst = 32'd201348700;
      23026: inst = 32'd203449168;
      23027: inst = 32'd136314880;
      23028: inst = 32'd268468224;
      23029: inst = 32'd201348701;
      23030: inst = 32'd203449168;
      23031: inst = 32'd136314880;
      23032: inst = 32'd268468224;
      23033: inst = 32'd201348702;
      23034: inst = 32'd203449168;
      23035: inst = 32'd136314880;
      23036: inst = 32'd268468224;
      23037: inst = 32'd201348703;
      23038: inst = 32'd203449168;
      23039: inst = 32'd136314880;
      23040: inst = 32'd268468224;
      23041: inst = 32'd201348704;
      23042: inst = 32'd203451247;
      23043: inst = 32'd136314880;
      23044: inst = 32'd268468224;
      23045: inst = 32'd201348705;
      23046: inst = 32'd203451247;
      23047: inst = 32'd136314880;
      23048: inst = 32'd268468224;
      23049: inst = 32'd201348706;
      23050: inst = 32'd203451247;
      23051: inst = 32'd136314880;
      23052: inst = 32'd268468224;
      23053: inst = 32'd201348707;
      23054: inst = 32'd203451247;
      23055: inst = 32'd136314880;
      23056: inst = 32'd268468224;
      23057: inst = 32'd201348708;
      23058: inst = 32'd203451247;
      23059: inst = 32'd136314880;
      23060: inst = 32'd268468224;
      23061: inst = 32'd201348709;
      23062: inst = 32'd203451247;
      23063: inst = 32'd136314880;
      23064: inst = 32'd268468224;
      23065: inst = 32'd201348710;
      23066: inst = 32'd203451247;
      23067: inst = 32'd136314880;
      23068: inst = 32'd268468224;
      23069: inst = 32'd201348711;
      23070: inst = 32'd203451247;
      23071: inst = 32'd136314880;
      23072: inst = 32'd268468224;
      23073: inst = 32'd201348712;
      23074: inst = 32'd203451247;
      23075: inst = 32'd136314880;
      23076: inst = 32'd268468224;
      23077: inst = 32'd201348713;
      23078: inst = 32'd203451247;
      23079: inst = 32'd136314880;
      23080: inst = 32'd268468224;
      23081: inst = 32'd201348714;
      23082: inst = 32'd203451247;
      23083: inst = 32'd136314880;
      23084: inst = 32'd268468224;
      23085: inst = 32'd201348715;
      23086: inst = 32'd203451247;
      23087: inst = 32'd136314880;
      23088: inst = 32'd268468224;
      23089: inst = 32'd201348716;
      23090: inst = 32'd203451247;
      23091: inst = 32'd136314880;
      23092: inst = 32'd268468224;
      23093: inst = 32'd201348717;
      23094: inst = 32'd203451247;
      23095: inst = 32'd136314880;
      23096: inst = 32'd268468224;
      23097: inst = 32'd201348718;
      23098: inst = 32'd203451247;
      23099: inst = 32'd136314880;
      23100: inst = 32'd268468224;
      23101: inst = 32'd201348719;
      23102: inst = 32'd203451247;
      23103: inst = 32'd136314880;
      23104: inst = 32'd268468224;
      23105: inst = 32'd201348720;
      23106: inst = 32'd203451248;
      23107: inst = 32'd136314880;
      23108: inst = 32'd268468224;
      23109: inst = 32'd201348721;
      23110: inst = 32'd203451248;
      23111: inst = 32'd136314880;
      23112: inst = 32'd268468224;
      23113: inst = 32'd201348722;
      23114: inst = 32'd203451215;
      23115: inst = 32'd136314880;
      23116: inst = 32'd268468224;
      23117: inst = 32'd201348723;
      23118: inst = 32'd203451214;
      23119: inst = 32'd136314880;
      23120: inst = 32'd268468224;
      23121: inst = 32'd201348724;
      23122: inst = 32'd203455440;
      23123: inst = 32'd136314880;
      23124: inst = 32'd268468224;
      23125: inst = 32'd201348725;
      23126: inst = 32'd203459666;
      23127: inst = 32'd136314880;
      23128: inst = 32'd268468224;
      23129: inst = 32'd201348726;
      23130: inst = 32'd203461778;
      23131: inst = 32'd136314880;
      23132: inst = 32'd268468224;
      23133: inst = 32'd201348727;
      23134: inst = 32'd203459665;
      23135: inst = 32'd136314880;
      23136: inst = 32'd268468224;
      23137: inst = 32'd201348728;
      23138: inst = 32'd203449100;
      23139: inst = 32'd136314880;
      23140: inst = 32'd268468224;
      23141: inst = 32'd201348729;
      23142: inst = 32'd203440680;
      23143: inst = 32'd136314880;
      23144: inst = 32'd268468224;
      23145: inst = 32'd201348730;
      23146: inst = 32'd203440680;
      23147: inst = 32'd136314880;
      23148: inst = 32'd268468224;
      23149: inst = 32'd201348731;
      23150: inst = 32'd203444874;
      23151: inst = 32'd136314880;
      23152: inst = 32'd268468224;
      23153: inst = 32'd201348732;
      23154: inst = 32'd203444841;
      23155: inst = 32'd136314880;
      23156: inst = 32'd268468224;
      23157: inst = 32'd201348733;
      23158: inst = 32'd203444906;
      23159: inst = 32'd136314880;
      23160: inst = 32'd268468224;
      23161: inst = 32'd201348734;
      23162: inst = 32'd203459664;
      23163: inst = 32'd136314880;
      23164: inst = 32'd268468224;
      23165: inst = 32'd201348735;
      23166: inst = 32'd203459665;
      23167: inst = 32'd136314880;
      23168: inst = 32'd268468224;
      23169: inst = 32'd201348736;
      23170: inst = 32'd203459730;
      23171: inst = 32'd136314880;
      23172: inst = 32'd268468224;
      23173: inst = 32'd201348737;
      23174: inst = 32'd203453358;
      23175: inst = 32'd136314880;
      23176: inst = 32'd268468224;
      23177: inst = 32'd201348738;
      23178: inst = 32'd203451213;
      23179: inst = 32'd136314880;
      23180: inst = 32'd268468224;
      23181: inst = 32'd201348739;
      23182: inst = 32'd203459730;
      23183: inst = 32'd136314880;
      23184: inst = 32'd268468224;
      23185: inst = 32'd201348740;
      23186: inst = 32'd203459698;
      23187: inst = 32'd136314880;
      23188: inst = 32'd268468224;
      23189: inst = 32'd201348741;
      23190: inst = 32'd203459697;
      23191: inst = 32'd136314880;
      23192: inst = 32'd268468224;
      23193: inst = 32'd201348742;
      23194: inst = 32'd203459665;
      23195: inst = 32'd136314880;
      23196: inst = 32'd268468224;
      23197: inst = 32'd201348743;
      23198: inst = 32'd203457520;
      23199: inst = 32'd136314880;
      23200: inst = 32'd268468224;
      23201: inst = 32'd201348744;
      23202: inst = 32'd203444875;
      23203: inst = 32'd136314880;
      23204: inst = 32'd268468224;
      23205: inst = 32'd201348745;
      23206: inst = 32'd203444842;
      23207: inst = 32'd136314880;
      23208: inst = 32'd268468224;
      23209: inst = 32'd201348746;
      23210: inst = 32'd203451247;
      23211: inst = 32'd136314880;
      23212: inst = 32'd268468224;
      23213: inst = 32'd201348747;
      23214: inst = 32'd203451247;
      23215: inst = 32'd136314880;
      23216: inst = 32'd268468224;
      23217: inst = 32'd201348748;
      23218: inst = 32'd203451215;
      23219: inst = 32'd136314880;
      23220: inst = 32'd268468224;
      23221: inst = 32'd201348749;
      23222: inst = 32'd203451215;
      23223: inst = 32'd136314880;
      23224: inst = 32'd268468224;
      23225: inst = 32'd201348750;
      23226: inst = 32'd203451215;
      23227: inst = 32'd136314880;
      23228: inst = 32'd268468224;
      23229: inst = 32'd201348751;
      23230: inst = 32'd203451248;
      23231: inst = 32'd136314880;
      23232: inst = 32'd268468224;
      23233: inst = 32'd201348752;
      23234: inst = 32'd203451248;
      23235: inst = 32'd136314880;
      23236: inst = 32'd268468224;
      23237: inst = 32'd201348753;
      23238: inst = 32'd203451215;
      23239: inst = 32'd136314880;
      23240: inst = 32'd268468224;
      23241: inst = 32'd201348754;
      23242: inst = 32'd203451215;
      23243: inst = 32'd136314880;
      23244: inst = 32'd268468224;
      23245: inst = 32'd201348755;
      23246: inst = 32'd203451215;
      23247: inst = 32'd136314880;
      23248: inst = 32'd268468224;
      23249: inst = 32'd201348756;
      23250: inst = 32'd203451247;
      23251: inst = 32'd136314880;
      23252: inst = 32'd268468224;
      23253: inst = 32'd201348757;
      23254: inst = 32'd203451247;
      23255: inst = 32'd136314880;
      23256: inst = 32'd268468224;
      23257: inst = 32'd201348758;
      23258: inst = 32'd203444842;
      23259: inst = 32'd136314880;
      23260: inst = 32'd268468224;
      23261: inst = 32'd201348759;
      23262: inst = 32'd203444875;
      23263: inst = 32'd136314880;
      23264: inst = 32'd268468224;
      23265: inst = 32'd201348760;
      23266: inst = 32'd203455472;
      23267: inst = 32'd136314880;
      23268: inst = 32'd268468224;
      23269: inst = 32'd201348761;
      23270: inst = 32'd203459698;
      23271: inst = 32'd136314880;
      23272: inst = 32'd268468224;
      23273: inst = 32'd201348762;
      23274: inst = 32'd203459697;
      23275: inst = 32'd136314880;
      23276: inst = 32'd268468224;
      23277: inst = 32'd201348763;
      23278: inst = 32'd203459697;
      23279: inst = 32'd136314880;
      23280: inst = 32'd268468224;
      23281: inst = 32'd201348764;
      23282: inst = 32'd203459698;
      23283: inst = 32'd136314880;
      23284: inst = 32'd268468224;
      23285: inst = 32'd201348765;
      23286: inst = 32'd203451245;
      23287: inst = 32'd136314880;
      23288: inst = 32'd268468224;
      23289: inst = 32'd201348766;
      23290: inst = 32'd203453359;
      23291: inst = 32'd136314880;
      23292: inst = 32'd268468224;
      23293: inst = 32'd201348767;
      23294: inst = 32'd203459730;
      23295: inst = 32'd136314880;
      23296: inst = 32'd268468224;
      23297: inst = 32'd201348768;
      23298: inst = 32'd203459666;
      23299: inst = 32'd136314880;
      23300: inst = 32'd268468224;
      23301: inst = 32'd201348769;
      23302: inst = 32'd203459666;
      23303: inst = 32'd136314880;
      23304: inst = 32'd268468224;
      23305: inst = 32'd201348770;
      23306: inst = 32'd203444907;
      23307: inst = 32'd136314880;
      23308: inst = 32'd268468224;
      23309: inst = 32'd201348771;
      23310: inst = 32'd203442794;
      23311: inst = 32'd136314880;
      23312: inst = 32'd268468224;
      23313: inst = 32'd201348772;
      23314: inst = 32'd203444875;
      23315: inst = 32'd136314880;
      23316: inst = 32'd268468224;
      23317: inst = 32'd201348773;
      23318: inst = 32'd203440681;
      23319: inst = 32'd136314880;
      23320: inst = 32'd268468224;
      23321: inst = 32'd201348774;
      23322: inst = 32'd203440681;
      23323: inst = 32'd136314880;
      23324: inst = 32'd268468224;
      23325: inst = 32'd201348775;
      23326: inst = 32'd203449101;
      23327: inst = 32'd136314880;
      23328: inst = 32'd268468224;
      23329: inst = 32'd201348776;
      23330: inst = 32'd203459666;
      23331: inst = 32'd136314880;
      23332: inst = 32'd268468224;
      23333: inst = 32'd201348777;
      23334: inst = 32'd203461746;
      23335: inst = 32'd136314880;
      23336: inst = 32'd268468224;
      23337: inst = 32'd201348778;
      23338: inst = 32'd203459634;
      23339: inst = 32'd136314880;
      23340: inst = 32'd268468224;
      23341: inst = 32'd201348779;
      23342: inst = 32'd203455408;
      23343: inst = 32'd136314880;
      23344: inst = 32'd268468224;
      23345: inst = 32'd201348780;
      23346: inst = 32'd203451215;
      23347: inst = 32'd136314880;
      23348: inst = 32'd268468224;
      23349: inst = 32'd201348781;
      23350: inst = 32'd203451215;
      23351: inst = 32'd136314880;
      23352: inst = 32'd268468224;
      23353: inst = 32'd201348782;
      23354: inst = 32'd203451248;
      23355: inst = 32'd136314880;
      23356: inst = 32'd268468224;
      23357: inst = 32'd201348783;
      23358: inst = 32'd203451216;
      23359: inst = 32'd136314880;
      23360: inst = 32'd268468224;
      23361: inst = 32'd201348784;
      23362: inst = 32'd203449168;
      23363: inst = 32'd136314880;
      23364: inst = 32'd268468224;
      23365: inst = 32'd201348785;
      23366: inst = 32'd203449168;
      23367: inst = 32'd136314880;
      23368: inst = 32'd268468224;
      23369: inst = 32'd201348786;
      23370: inst = 32'd203449168;
      23371: inst = 32'd136314880;
      23372: inst = 32'd268468224;
      23373: inst = 32'd201348787;
      23374: inst = 32'd203449168;
      23375: inst = 32'd136314880;
      23376: inst = 32'd268468224;
      23377: inst = 32'd201348788;
      23378: inst = 32'd203449168;
      23379: inst = 32'd136314880;
      23380: inst = 32'd268468224;
      23381: inst = 32'd201348789;
      23382: inst = 32'd203449168;
      23383: inst = 32'd136314880;
      23384: inst = 32'd268468224;
      23385: inst = 32'd201348790;
      23386: inst = 32'd203449168;
      23387: inst = 32'd136314880;
      23388: inst = 32'd268468224;
      23389: inst = 32'd201348791;
      23390: inst = 32'd203449168;
      23391: inst = 32'd136314880;
      23392: inst = 32'd268468224;
      23393: inst = 32'd201348792;
      23394: inst = 32'd203449168;
      23395: inst = 32'd136314880;
      23396: inst = 32'd268468224;
      23397: inst = 32'd201348793;
      23398: inst = 32'd203449168;
      23399: inst = 32'd136314880;
      23400: inst = 32'd268468224;
      23401: inst = 32'd201348794;
      23402: inst = 32'd203449168;
      23403: inst = 32'd136314880;
      23404: inst = 32'd268468224;
      23405: inst = 32'd201348795;
      23406: inst = 32'd203449168;
      23407: inst = 32'd136314880;
      23408: inst = 32'd268468224;
      23409: inst = 32'd201348796;
      23410: inst = 32'd203449168;
      23411: inst = 32'd136314880;
      23412: inst = 32'd268468224;
      23413: inst = 32'd201348797;
      23414: inst = 32'd203449168;
      23415: inst = 32'd136314880;
      23416: inst = 32'd268468224;
      23417: inst = 32'd201348798;
      23418: inst = 32'd203449168;
      23419: inst = 32'd136314880;
      23420: inst = 32'd268468224;
      23421: inst = 32'd201348799;
      23422: inst = 32'd203449168;
      23423: inst = 32'd136314880;
      23424: inst = 32'd268468224;
      23425: inst = 32'd201348800;
      23426: inst = 32'd203451216;
      23427: inst = 32'd136314880;
      23428: inst = 32'd268468224;
      23429: inst = 32'd201348801;
      23430: inst = 32'd203451216;
      23431: inst = 32'd136314880;
      23432: inst = 32'd268468224;
      23433: inst = 32'd201348802;
      23434: inst = 32'd203451216;
      23435: inst = 32'd136314880;
      23436: inst = 32'd268468224;
      23437: inst = 32'd201348803;
      23438: inst = 32'd203451216;
      23439: inst = 32'd136314880;
      23440: inst = 32'd268468224;
      23441: inst = 32'd201348804;
      23442: inst = 32'd203451216;
      23443: inst = 32'd136314880;
      23444: inst = 32'd268468224;
      23445: inst = 32'd201348805;
      23446: inst = 32'd203451216;
      23447: inst = 32'd136314880;
      23448: inst = 32'd268468224;
      23449: inst = 32'd201348806;
      23450: inst = 32'd203451216;
      23451: inst = 32'd136314880;
      23452: inst = 32'd268468224;
      23453: inst = 32'd201348807;
      23454: inst = 32'd203451216;
      23455: inst = 32'd136314880;
      23456: inst = 32'd268468224;
      23457: inst = 32'd201348808;
      23458: inst = 32'd203451216;
      23459: inst = 32'd136314880;
      23460: inst = 32'd268468224;
      23461: inst = 32'd201348809;
      23462: inst = 32'd203451216;
      23463: inst = 32'd136314880;
      23464: inst = 32'd268468224;
      23465: inst = 32'd201348810;
      23466: inst = 32'd203451216;
      23467: inst = 32'd136314880;
      23468: inst = 32'd268468224;
      23469: inst = 32'd201348811;
      23470: inst = 32'd203451216;
      23471: inst = 32'd136314880;
      23472: inst = 32'd268468224;
      23473: inst = 32'd201348812;
      23474: inst = 32'd203451216;
      23475: inst = 32'd136314880;
      23476: inst = 32'd268468224;
      23477: inst = 32'd201348813;
      23478: inst = 32'd203451216;
      23479: inst = 32'd136314880;
      23480: inst = 32'd268468224;
      23481: inst = 32'd201348814;
      23482: inst = 32'd203451216;
      23483: inst = 32'd136314880;
      23484: inst = 32'd268468224;
      23485: inst = 32'd201348815;
      23486: inst = 32'd203451216;
      23487: inst = 32'd136314880;
      23488: inst = 32'd268468224;
      23489: inst = 32'd201348816;
      23490: inst = 32'd203451249;
      23491: inst = 32'd136314880;
      23492: inst = 32'd268468224;
      23493: inst = 32'd201348817;
      23494: inst = 32'd203449135;
      23495: inst = 32'd136314880;
      23496: inst = 32'd268468224;
      23497: inst = 32'd201348818;
      23498: inst = 32'd203449135;
      23499: inst = 32'd136314880;
      23500: inst = 32'd268468224;
      23501: inst = 32'd201348819;
      23502: inst = 32'd203455408;
      23503: inst = 32'd136314880;
      23504: inst = 32'd268468224;
      23505: inst = 32'd201348820;
      23506: inst = 32'd203459666;
      23507: inst = 32'd136314880;
      23508: inst = 32'd268468224;
      23509: inst = 32'd201348821;
      23510: inst = 32'd203459698;
      23511: inst = 32'd136314880;
      23512: inst = 32'd268468224;
      23513: inst = 32'd201348822;
      23514: inst = 32'd203459697;
      23515: inst = 32'd136314880;
      23516: inst = 32'd268468224;
      23517: inst = 32'd201348823;
      23518: inst = 32'd203459697;
      23519: inst = 32'd136314880;
      23520: inst = 32'd268468224;
      23521: inst = 32'd201348824;
      23522: inst = 32'd203459697;
      23523: inst = 32'd136314880;
      23524: inst = 32'd268468224;
      23525: inst = 32'd201348825;
      23526: inst = 32'd203463859;
      23527: inst = 32'd136314880;
      23528: inst = 32'd268468224;
      23529: inst = 32'd201348826;
      23530: inst = 32'd203459665;
      23531: inst = 32'd136314880;
      23532: inst = 32'd268468224;
      23533: inst = 32'd201348827;
      23534: inst = 32'd203461811;
      23535: inst = 32'd136314880;
      23536: inst = 32'd268468224;
      23537: inst = 32'd201348828;
      23538: inst = 32'd203459698;
      23539: inst = 32'd136314880;
      23540: inst = 32'd268468224;
      23541: inst = 32'd201348829;
      23542: inst = 32'd203457617;
      23543: inst = 32'd136314880;
      23544: inst = 32'd268468224;
      23545: inst = 32'd201348830;
      23546: inst = 32'd203459665;
      23547: inst = 32'd136314880;
      23548: inst = 32'd268468224;
      23549: inst = 32'd201348831;
      23550: inst = 32'd203459698;
      23551: inst = 32'd136314880;
      23552: inst = 32'd268468224;
      23553: inst = 32'd201348832;
      23554: inst = 32'd203459729;
      23555: inst = 32'd136314880;
      23556: inst = 32'd268468224;
      23557: inst = 32'd201348833;
      23558: inst = 32'd203455439;
      23559: inst = 32'd136314880;
      23560: inst = 32'd268468224;
      23561: inst = 32'd201348834;
      23562: inst = 32'd203455471;
      23563: inst = 32'd136314880;
      23564: inst = 32'd268468224;
      23565: inst = 32'd201348835;
      23566: inst = 32'd203459698;
      23567: inst = 32'd136314880;
      23568: inst = 32'd268468224;
      23569: inst = 32'd201348836;
      23570: inst = 32'd203461778;
      23571: inst = 32'd136314880;
      23572: inst = 32'd268468224;
      23573: inst = 32'd201348837;
      23574: inst = 32'd203459665;
      23575: inst = 32'd136314880;
      23576: inst = 32'd268468224;
      23577: inst = 32'd201348838;
      23578: inst = 32'd203459666;
      23579: inst = 32'd136314880;
      23580: inst = 32'd268468224;
      23581: inst = 32'd201348839;
      23582: inst = 32'd203453327;
      23583: inst = 32'd136314880;
      23584: inst = 32'd268468224;
      23585: inst = 32'd201348840;
      23586: inst = 32'd203444875;
      23587: inst = 32'd136314880;
      23588: inst = 32'd268468224;
      23589: inst = 32'd201348841;
      23590: inst = 32'd203444875;
      23591: inst = 32'd136314880;
      23592: inst = 32'd268468224;
      23593: inst = 32'd201348842;
      23594: inst = 32'd203451247;
      23595: inst = 32'd136314880;
      23596: inst = 32'd268468224;
      23597: inst = 32'd201348843;
      23598: inst = 32'd203451247;
      23599: inst = 32'd136314880;
      23600: inst = 32'd268468224;
      23601: inst = 32'd201348844;
      23602: inst = 32'd203451247;
      23603: inst = 32'd136314880;
      23604: inst = 32'd268468224;
      23605: inst = 32'd201348845;
      23606: inst = 32'd203449199;
      23607: inst = 32'd136314880;
      23608: inst = 32'd268468224;
      23609: inst = 32'd201348846;
      23610: inst = 32'd203449200;
      23611: inst = 32'd136314880;
      23612: inst = 32'd268468224;
      23613: inst = 32'd201348847;
      23614: inst = 32'd203449200;
      23615: inst = 32'd136314880;
      23616: inst = 32'd268468224;
      23617: inst = 32'd201348848;
      23618: inst = 32'd203449200;
      23619: inst = 32'd136314880;
      23620: inst = 32'd268468224;
      23621: inst = 32'd201348849;
      23622: inst = 32'd203449200;
      23623: inst = 32'd136314880;
      23624: inst = 32'd268468224;
      23625: inst = 32'd201348850;
      23626: inst = 32'd203449199;
      23627: inst = 32'd136314880;
      23628: inst = 32'd268468224;
      23629: inst = 32'd201348851;
      23630: inst = 32'd203451247;
      23631: inst = 32'd136314880;
      23632: inst = 32'd268468224;
      23633: inst = 32'd201348852;
      23634: inst = 32'd203451247;
      23635: inst = 32'd136314880;
      23636: inst = 32'd268468224;
      23637: inst = 32'd201348853;
      23638: inst = 32'd203451247;
      23639: inst = 32'd136314880;
      23640: inst = 32'd268468224;
      23641: inst = 32'd201348854;
      23642: inst = 32'd203444875;
      23643: inst = 32'd136314880;
      23644: inst = 32'd268468224;
      23645: inst = 32'd201348855;
      23646: inst = 32'd203444875;
      23647: inst = 32'd136314880;
      23648: inst = 32'd268468224;
      23649: inst = 32'd201348856;
      23650: inst = 32'd203453294;
      23651: inst = 32'd136314880;
      23652: inst = 32'd268468224;
      23653: inst = 32'd201348857;
      23654: inst = 32'd203459666;
      23655: inst = 32'd136314880;
      23656: inst = 32'd268468224;
      23657: inst = 32'd201348858;
      23658: inst = 32'd203459665;
      23659: inst = 32'd136314880;
      23660: inst = 32'd268468224;
      23661: inst = 32'd201348859;
      23662: inst = 32'd203459698;
      23663: inst = 32'd136314880;
      23664: inst = 32'd268468224;
      23665: inst = 32'd201348860;
      23666: inst = 32'd203459697;
      23667: inst = 32'd136314880;
      23668: inst = 32'd268468224;
      23669: inst = 32'd201348861;
      23670: inst = 32'd203455471;
      23671: inst = 32'd136314880;
      23672: inst = 32'd268468224;
      23673: inst = 32'd201348862;
      23674: inst = 32'd203455439;
      23675: inst = 32'd136314880;
      23676: inst = 32'd268468224;
      23677: inst = 32'd201348863;
      23678: inst = 32'd203459697;
      23679: inst = 32'd136314880;
      23680: inst = 32'd268468224;
      23681: inst = 32'd201348864;
      23682: inst = 32'd203459698;
      23683: inst = 32'd136314880;
      23684: inst = 32'd268468224;
      23685: inst = 32'd201348865;
      23686: inst = 32'd203459665;
      23687: inst = 32'd136314880;
      23688: inst = 32'd268468224;
      23689: inst = 32'd201348866;
      23690: inst = 32'd203459665;
      23691: inst = 32'd136314880;
      23692: inst = 32'd268468224;
      23693: inst = 32'd201348867;
      23694: inst = 32'd203459698;
      23695: inst = 32'd136314880;
      23696: inst = 32'd268468224;
      23697: inst = 32'd201348868;
      23698: inst = 32'd203461811;
      23699: inst = 32'd136314880;
      23700: inst = 32'd268468224;
      23701: inst = 32'd201348869;
      23702: inst = 32'd203459665;
      23703: inst = 32'd136314880;
      23704: inst = 32'd268468224;
      23705: inst = 32'd201348870;
      23706: inst = 32'd203461811;
      23707: inst = 32'd136314880;
      23708: inst = 32'd268468224;
      23709: inst = 32'd201348871;
      23710: inst = 32'd203459698;
      23711: inst = 32'd136314880;
      23712: inst = 32'd268468224;
      23713: inst = 32'd201348872;
      23714: inst = 32'd203459698;
      23715: inst = 32'd136314880;
      23716: inst = 32'd268468224;
      23717: inst = 32'd201348873;
      23718: inst = 32'd203461746;
      23719: inst = 32'd136314880;
      23720: inst = 32'd268468224;
      23721: inst = 32'd201348874;
      23722: inst = 32'd203459698;
      23723: inst = 32'd136314880;
      23724: inst = 32'd268468224;
      23725: inst = 32'd201348875;
      23726: inst = 32'd203459634;
      23727: inst = 32'd136314880;
      23728: inst = 32'd268468224;
      23729: inst = 32'd201348876;
      23730: inst = 32'd203455408;
      23731: inst = 32'd136314880;
      23732: inst = 32'd268468224;
      23733: inst = 32'd201348877;
      23734: inst = 32'd203449167;
      23735: inst = 32'd136314880;
      23736: inst = 32'd268468224;
      23737: inst = 32'd201348878;
      23738: inst = 32'd203449167;
      23739: inst = 32'd136314880;
      23740: inst = 32'd268468224;
      23741: inst = 32'd201348879;
      23742: inst = 32'd203451248;
      23743: inst = 32'd136314880;
      23744: inst = 32'd268468224;
      23745: inst = 32'd201348880;
      23746: inst = 32'd203449200;
      23747: inst = 32'd136314880;
      23748: inst = 32'd268468224;
      23749: inst = 32'd201348881;
      23750: inst = 32'd203449200;
      23751: inst = 32'd136314880;
      23752: inst = 32'd268468224;
      23753: inst = 32'd201348882;
      23754: inst = 32'd203449200;
      23755: inst = 32'd136314880;
      23756: inst = 32'd268468224;
      23757: inst = 32'd201348883;
      23758: inst = 32'd203449200;
      23759: inst = 32'd136314880;
      23760: inst = 32'd268468224;
      23761: inst = 32'd201348884;
      23762: inst = 32'd203449200;
      23763: inst = 32'd136314880;
      23764: inst = 32'd268468224;
      23765: inst = 32'd201348885;
      23766: inst = 32'd203449200;
      23767: inst = 32'd136314880;
      23768: inst = 32'd268468224;
      23769: inst = 32'd201348886;
      23770: inst = 32'd203449200;
      23771: inst = 32'd136314880;
      23772: inst = 32'd268468224;
      23773: inst = 32'd201348887;
      23774: inst = 32'd203449200;
      23775: inst = 32'd136314880;
      23776: inst = 32'd268468224;
      23777: inst = 32'd201348888;
      23778: inst = 32'd203449200;
      23779: inst = 32'd136314880;
      23780: inst = 32'd268468224;
      23781: inst = 32'd201348889;
      23782: inst = 32'd203449200;
      23783: inst = 32'd136314880;
      23784: inst = 32'd268468224;
      23785: inst = 32'd201348890;
      23786: inst = 32'd203449200;
      23787: inst = 32'd136314880;
      23788: inst = 32'd268468224;
      23789: inst = 32'd201348891;
      23790: inst = 32'd203449200;
      23791: inst = 32'd136314880;
      23792: inst = 32'd268468224;
      23793: inst = 32'd201348892;
      23794: inst = 32'd203449200;
      23795: inst = 32'd136314880;
      23796: inst = 32'd268468224;
      23797: inst = 32'd201348893;
      23798: inst = 32'd203449200;
      23799: inst = 32'd136314880;
      23800: inst = 32'd268468224;
      23801: inst = 32'd201348894;
      23802: inst = 32'd203449200;
      23803: inst = 32'd136314880;
      23804: inst = 32'd268468224;
      23805: inst = 32'd201348895;
      23806: inst = 32'd203449200;
      23807: inst = 32'd136314880;
      23808: inst = 32'd268468224;
      23809: inst = 32'd201348896;
      23810: inst = 32'd203451216;
      23811: inst = 32'd136314880;
      23812: inst = 32'd268468224;
      23813: inst = 32'd201348897;
      23814: inst = 32'd203451216;
      23815: inst = 32'd136314880;
      23816: inst = 32'd268468224;
      23817: inst = 32'd201348898;
      23818: inst = 32'd203451216;
      23819: inst = 32'd136314880;
      23820: inst = 32'd268468224;
      23821: inst = 32'd201348899;
      23822: inst = 32'd203451216;
      23823: inst = 32'd136314880;
      23824: inst = 32'd268468224;
      23825: inst = 32'd201348900;
      23826: inst = 32'd203451216;
      23827: inst = 32'd136314880;
      23828: inst = 32'd268468224;
      23829: inst = 32'd201348901;
      23830: inst = 32'd203451216;
      23831: inst = 32'd136314880;
      23832: inst = 32'd268468224;
      23833: inst = 32'd201348902;
      23834: inst = 32'd203451216;
      23835: inst = 32'd136314880;
      23836: inst = 32'd268468224;
      23837: inst = 32'd201348903;
      23838: inst = 32'd203451216;
      23839: inst = 32'd136314880;
      23840: inst = 32'd268468224;
      23841: inst = 32'd201348904;
      23842: inst = 32'd203451216;
      23843: inst = 32'd136314880;
      23844: inst = 32'd268468224;
      23845: inst = 32'd201348905;
      23846: inst = 32'd203451216;
      23847: inst = 32'd136314880;
      23848: inst = 32'd268468224;
      23849: inst = 32'd201348906;
      23850: inst = 32'd203451216;
      23851: inst = 32'd136314880;
      23852: inst = 32'd268468224;
      23853: inst = 32'd201348907;
      23854: inst = 32'd203451216;
      23855: inst = 32'd136314880;
      23856: inst = 32'd268468224;
      23857: inst = 32'd201348908;
      23858: inst = 32'd203451216;
      23859: inst = 32'd136314880;
      23860: inst = 32'd268468224;
      23861: inst = 32'd201348909;
      23862: inst = 32'd203451216;
      23863: inst = 32'd136314880;
      23864: inst = 32'd268468224;
      23865: inst = 32'd201348910;
      23866: inst = 32'd203451216;
      23867: inst = 32'd136314880;
      23868: inst = 32'd268468224;
      23869: inst = 32'd201348911;
      23870: inst = 32'd203451216;
      23871: inst = 32'd136314880;
      23872: inst = 32'd268468224;
      23873: inst = 32'd201348912;
      23874: inst = 32'd203451217;
      23875: inst = 32'd136314880;
      23876: inst = 32'd268468224;
      23877: inst = 32'd201348913;
      23878: inst = 32'd203449168;
      23879: inst = 32'd136314880;
      23880: inst = 32'd268468224;
      23881: inst = 32'd201348914;
      23882: inst = 32'd203451280;
      23883: inst = 32'd136314880;
      23884: inst = 32'd268468224;
      23885: inst = 32'd201348915;
      23886: inst = 32'd203457586;
      23887: inst = 32'd136314880;
      23888: inst = 32'd268468224;
      23889: inst = 32'd201348916;
      23890: inst = 32'd203459698;
      23891: inst = 32'd136314880;
      23892: inst = 32'd268468224;
      23893: inst = 32'd201348917;
      23894: inst = 32'd203459698;
      23895: inst = 32'd136314880;
      23896: inst = 32'd268468224;
      23897: inst = 32'd201348918;
      23898: inst = 32'd203459665;
      23899: inst = 32'd136314880;
      23900: inst = 32'd268468224;
      23901: inst = 32'd201348919;
      23902: inst = 32'd203461745;
      23903: inst = 32'd136314880;
      23904: inst = 32'd268468224;
      23905: inst = 32'd201348920;
      23906: inst = 32'd203457584;
      23907: inst = 32'd136314880;
      23908: inst = 32'd268468224;
      23909: inst = 32'd201348921;
      23910: inst = 32'd203461778;
      23911: inst = 32'd136314880;
      23912: inst = 32'd268468224;
      23913: inst = 32'd201348922;
      23914: inst = 32'd203457585;
      23915: inst = 32'd136314880;
      23916: inst = 32'd268468224;
      23917: inst = 32'd201348923;
      23918: inst = 32'd203459665;
      23919: inst = 32'd136314880;
      23920: inst = 32'd268468224;
      23921: inst = 32'd201348924;
      23922: inst = 32'd203459698;
      23923: inst = 32'd136314880;
      23924: inst = 32'd268468224;
      23925: inst = 32'd201348925;
      23926: inst = 32'd203459698;
      23927: inst = 32'd136314880;
      23928: inst = 32'd268468224;
      23929: inst = 32'd201348926;
      23930: inst = 32'd203457618;
      23931: inst = 32'd136314880;
      23932: inst = 32'd268468224;
      23933: inst = 32'd201348927;
      23934: inst = 32'd203461843;
      23935: inst = 32'd136314880;
      23936: inst = 32'd268468224;
      23937: inst = 32'd201348928;
      23938: inst = 32'd203459697;
      23939: inst = 32'd136314880;
      23940: inst = 32'd268468224;
      23941: inst = 32'd201348929;
      23942: inst = 32'd203457583;
      23943: inst = 32'd136314880;
      23944: inst = 32'd268468224;
      23945: inst = 32'd201348930;
      23946: inst = 32'd203459664;
      23947: inst = 32'd136314880;
      23948: inst = 32'd268468224;
      23949: inst = 32'd201348931;
      23950: inst = 32'd203459697;
      23951: inst = 32'd136314880;
      23952: inst = 32'd268468224;
      23953: inst = 32'd201348932;
      23954: inst = 32'd203459697;
      23955: inst = 32'd136314880;
      23956: inst = 32'd268468224;
      23957: inst = 32'd201348933;
      23958: inst = 32'd203459698;
      23959: inst = 32'd136314880;
      23960: inst = 32'd268468224;
      23961: inst = 32'd201348934;
      23962: inst = 32'd203459666;
      23963: inst = 32'd136314880;
      23964: inst = 32'd268468224;
      23965: inst = 32'd201348935;
      23966: inst = 32'd203449101;
      23967: inst = 32'd136314880;
      23968: inst = 32'd268468224;
      23969: inst = 32'd201348936;
      23970: inst = 32'd203444876;
      23971: inst = 32'd136314880;
      23972: inst = 32'd268468224;
      23973: inst = 32'd201348937;
      23974: inst = 32'd203442827;
      23975: inst = 32'd136314880;
      23976: inst = 32'd268468224;
      23977: inst = 32'd201348938;
      23978: inst = 32'd203451247;
      23979: inst = 32'd136314880;
      23980: inst = 32'd268468224;
      23981: inst = 32'd201348939;
      23982: inst = 32'd203449199;
      23983: inst = 32'd136314880;
      23984: inst = 32'd268468224;
      23985: inst = 32'd201348940;
      23986: inst = 32'd203449199;
      23987: inst = 32'd136314880;
      23988: inst = 32'd268468224;
      23989: inst = 32'd201348941;
      23990: inst = 32'd203449200;
      23991: inst = 32'd136314880;
      23992: inst = 32'd268468224;
      23993: inst = 32'd201348942;
      23994: inst = 32'd203449200;
      23995: inst = 32'd136314880;
      23996: inst = 32'd268468224;
      23997: inst = 32'd201348943;
      23998: inst = 32'd203449200;
      23999: inst = 32'd136314880;
      24000: inst = 32'd268468224;
      24001: inst = 32'd201348944;
      24002: inst = 32'd203449200;
      24003: inst = 32'd136314880;
      24004: inst = 32'd268468224;
      24005: inst = 32'd201348945;
      24006: inst = 32'd203449200;
      24007: inst = 32'd136314880;
      24008: inst = 32'd268468224;
      24009: inst = 32'd201348946;
      24010: inst = 32'd203449200;
      24011: inst = 32'd136314880;
      24012: inst = 32'd268468224;
      24013: inst = 32'd201348947;
      24014: inst = 32'd203449199;
      24015: inst = 32'd136314880;
      24016: inst = 32'd268468224;
      24017: inst = 32'd201348948;
      24018: inst = 32'd203449199;
      24019: inst = 32'd136314880;
      24020: inst = 32'd268468224;
      24021: inst = 32'd201348949;
      24022: inst = 32'd203451247;
      24023: inst = 32'd136314880;
      24024: inst = 32'd268468224;
      24025: inst = 32'd201348950;
      24026: inst = 32'd203442827;
      24027: inst = 32'd136314880;
      24028: inst = 32'd268468224;
      24029: inst = 32'd201348951;
      24030: inst = 32'd203444876;
      24031: inst = 32'd136314880;
      24032: inst = 32'd268468224;
      24033: inst = 32'd201348952;
      24034: inst = 32'd203449133;
      24035: inst = 32'd136314880;
      24036: inst = 32'd268468224;
      24037: inst = 32'd201348953;
      24038: inst = 32'd203459666;
      24039: inst = 32'd136314880;
      24040: inst = 32'd268468224;
      24041: inst = 32'd201348954;
      24042: inst = 32'd203459698;
      24043: inst = 32'd136314880;
      24044: inst = 32'd268468224;
      24045: inst = 32'd201348955;
      24046: inst = 32'd203459698;
      24047: inst = 32'd136314880;
      24048: inst = 32'd268468224;
      24049: inst = 32'd201348956;
      24050: inst = 32'd203459697;
      24051: inst = 32'd136314880;
      24052: inst = 32'd268468224;
      24053: inst = 32'd201348957;
      24054: inst = 32'd203459664;
      24055: inst = 32'd136314880;
      24056: inst = 32'd268468224;
      24057: inst = 32'd201348958;
      24058: inst = 32'd203457551;
      24059: inst = 32'd136314880;
      24060: inst = 32'd268468224;
      24061: inst = 32'd201348959;
      24062: inst = 32'd203459697;
      24063: inst = 32'd136314880;
      24064: inst = 32'd268468224;
      24065: inst = 32'd201348960;
      24066: inst = 32'd203463858;
      24067: inst = 32'd136314880;
      24068: inst = 32'd268468224;
      24069: inst = 32'd201348961;
      24070: inst = 32'd203459664;
      24071: inst = 32'd136314880;
      24072: inst = 32'd268468224;
      24073: inst = 32'd201348962;
      24074: inst = 32'd203459697;
      24075: inst = 32'd136314880;
      24076: inst = 32'd268468224;
      24077: inst = 32'd201348963;
      24078: inst = 32'd203459697;
      24079: inst = 32'd136314880;
      24080: inst = 32'd268468224;
      24081: inst = 32'd201348964;
      24082: inst = 32'd203457617;
      24083: inst = 32'd136314880;
      24084: inst = 32'd268468224;
      24085: inst = 32'd201348965;
      24086: inst = 32'd203457584;
      24087: inst = 32'd136314880;
      24088: inst = 32'd268468224;
      24089: inst = 32'd201348966;
      24090: inst = 32'd203461810;
      24091: inst = 32'd136314880;
      24092: inst = 32'd268468224;
      24093: inst = 32'd201348967;
      24094: inst = 32'd203457584;
      24095: inst = 32'd136314880;
      24096: inst = 32'd268468224;
      24097: inst = 32'd201348968;
      24098: inst = 32'd203459697;
      24099: inst = 32'd136314880;
      24100: inst = 32'd268468224;
      24101: inst = 32'd201348969;
      24102: inst = 32'd203459697;
      24103: inst = 32'd136314880;
      24104: inst = 32'd268468224;
      24105: inst = 32'd201348970;
      24106: inst = 32'd203459698;
      24107: inst = 32'd136314880;
      24108: inst = 32'd268468224;
      24109: inst = 32'd201348971;
      24110: inst = 32'd203459730;
      24111: inst = 32'd136314880;
      24112: inst = 32'd268468224;
      24113: inst = 32'd201348972;
      24114: inst = 32'd203457585;
      24115: inst = 32'd136314880;
      24116: inst = 32'd268468224;
      24117: inst = 32'd201348973;
      24118: inst = 32'd203451280;
      24119: inst = 32'd136314880;
      24120: inst = 32'd268468224;
      24121: inst = 32'd201348974;
      24122: inst = 32'd203449199;
      24123: inst = 32'd136314880;
      24124: inst = 32'd268468224;
      24125: inst = 32'd201348975;
      24126: inst = 32'd203449232;
      24127: inst = 32'd136314880;
      24128: inst = 32'd268468224;
      24129: inst = 32'd201348976;
      24130: inst = 32'd203451216;
      24131: inst = 32'd136314880;
      24132: inst = 32'd268468224;
      24133: inst = 32'd201348977;
      24134: inst = 32'd203451216;
      24135: inst = 32'd136314880;
      24136: inst = 32'd268468224;
      24137: inst = 32'd201348978;
      24138: inst = 32'd203451216;
      24139: inst = 32'd136314880;
      24140: inst = 32'd268468224;
      24141: inst = 32'd201348979;
      24142: inst = 32'd203451216;
      24143: inst = 32'd136314880;
      24144: inst = 32'd268468224;
      24145: inst = 32'd201348980;
      24146: inst = 32'd203451216;
      24147: inst = 32'd136314880;
      24148: inst = 32'd268468224;
      24149: inst = 32'd201348981;
      24150: inst = 32'd203451216;
      24151: inst = 32'd136314880;
      24152: inst = 32'd268468224;
      24153: inst = 32'd201348982;
      24154: inst = 32'd203451216;
      24155: inst = 32'd136314880;
      24156: inst = 32'd268468224;
      24157: inst = 32'd201348983;
      24158: inst = 32'd203451216;
      24159: inst = 32'd136314880;
      24160: inst = 32'd268468224;
      24161: inst = 32'd201348984;
      24162: inst = 32'd203451216;
      24163: inst = 32'd136314880;
      24164: inst = 32'd268468224;
      24165: inst = 32'd201348985;
      24166: inst = 32'd203451216;
      24167: inst = 32'd136314880;
      24168: inst = 32'd268468224;
      24169: inst = 32'd201348986;
      24170: inst = 32'd203451216;
      24171: inst = 32'd136314880;
      24172: inst = 32'd268468224;
      24173: inst = 32'd201348987;
      24174: inst = 32'd203451216;
      24175: inst = 32'd136314880;
      24176: inst = 32'd268468224;
      24177: inst = 32'd201348988;
      24178: inst = 32'd203451216;
      24179: inst = 32'd136314880;
      24180: inst = 32'd268468224;
      24181: inst = 32'd201348989;
      24182: inst = 32'd203451216;
      24183: inst = 32'd136314880;
      24184: inst = 32'd268468224;
      24185: inst = 32'd201348990;
      24186: inst = 32'd203451216;
      24187: inst = 32'd136314880;
      24188: inst = 32'd268468224;
      24189: inst = 32'd201348991;
      24190: inst = 32'd203451216;
      24191: inst = 32'd136314880;
      24192: inst = 32'd268468224;
      24193: inst = 32'd201348992;
      24194: inst = 32'd203451216;
      24195: inst = 32'd136314880;
      24196: inst = 32'd268468224;
      24197: inst = 32'd201348993;
      24198: inst = 32'd203451216;
      24199: inst = 32'd136314880;
      24200: inst = 32'd268468224;
      24201: inst = 32'd201348994;
      24202: inst = 32'd203451216;
      24203: inst = 32'd136314880;
      24204: inst = 32'd268468224;
      24205: inst = 32'd201348995;
      24206: inst = 32'd203451216;
      24207: inst = 32'd136314880;
      24208: inst = 32'd268468224;
      24209: inst = 32'd201348996;
      24210: inst = 32'd203451216;
      24211: inst = 32'd136314880;
      24212: inst = 32'd268468224;
      24213: inst = 32'd201348997;
      24214: inst = 32'd203451216;
      24215: inst = 32'd136314880;
      24216: inst = 32'd268468224;
      24217: inst = 32'd201348998;
      24218: inst = 32'd203451216;
      24219: inst = 32'd136314880;
      24220: inst = 32'd268468224;
      24221: inst = 32'd201348999;
      24222: inst = 32'd203451216;
      24223: inst = 32'd136314880;
      24224: inst = 32'd268468224;
      24225: inst = 32'd201349000;
      24226: inst = 32'd203451216;
      24227: inst = 32'd136314880;
      24228: inst = 32'd268468224;
      24229: inst = 32'd201349001;
      24230: inst = 32'd203451216;
      24231: inst = 32'd136314880;
      24232: inst = 32'd268468224;
      24233: inst = 32'd201349002;
      24234: inst = 32'd203451216;
      24235: inst = 32'd136314880;
      24236: inst = 32'd268468224;
      24237: inst = 32'd201349003;
      24238: inst = 32'd203451216;
      24239: inst = 32'd136314880;
      24240: inst = 32'd268468224;
      24241: inst = 32'd201349004;
      24242: inst = 32'd203451216;
      24243: inst = 32'd136314880;
      24244: inst = 32'd268468224;
      24245: inst = 32'd201349005;
      24246: inst = 32'd203451216;
      24247: inst = 32'd136314880;
      24248: inst = 32'd268468224;
      24249: inst = 32'd201349006;
      24250: inst = 32'd203451216;
      24251: inst = 32'd136314880;
      24252: inst = 32'd268468224;
      24253: inst = 32'd201349007;
      24254: inst = 32'd203451216;
      24255: inst = 32'd136314880;
      24256: inst = 32'd268468224;
      24257: inst = 32'd201349008;
      24258: inst = 32'd203449136;
      24259: inst = 32'd136314880;
      24260: inst = 32'd268468224;
      24261: inst = 32'd201349009;
      24262: inst = 32'd203451281;
      24263: inst = 32'd136314880;
      24264: inst = 32'd268468224;
      24265: inst = 32'd201349010;
      24266: inst = 32'd203455474;
      24267: inst = 32'd136314880;
      24268: inst = 32'd268468224;
      24269: inst = 32'd201349011;
      24270: inst = 32'd203457619;
      24271: inst = 32'd136314880;
      24272: inst = 32'd268468224;
      24273: inst = 32'd201349012;
      24274: inst = 32'd203459698;
      24275: inst = 32'd136314880;
      24276: inst = 32'd268468224;
      24277: inst = 32'd201349013;
      24278: inst = 32'd203459698;
      24279: inst = 32'd136314880;
      24280: inst = 32'd268468224;
      24281: inst = 32'd201349014;
      24282: inst = 32'd203459665;
      24283: inst = 32'd136314880;
      24284: inst = 32'd268468224;
      24285: inst = 32'd201349015;
      24286: inst = 32'd203459665;
      24287: inst = 32'd136314880;
      24288: inst = 32'd268468224;
      24289: inst = 32'd201349016;
      24290: inst = 32'd203461746;
      24291: inst = 32'd136314880;
      24292: inst = 32'd268468224;
      24293: inst = 32'd201349017;
      24294: inst = 32'd203459665;
      24295: inst = 32'd136314880;
      24296: inst = 32'd268468224;
      24297: inst = 32'd201349018;
      24298: inst = 32'd203459698;
      24299: inst = 32'd136314880;
      24300: inst = 32'd268468224;
      24301: inst = 32'd201349019;
      24302: inst = 32'd203459666;
      24303: inst = 32'd136314880;
      24304: inst = 32'd268468224;
      24305: inst = 32'd201349020;
      24306: inst = 32'd203459731;
      24307: inst = 32'd136314880;
      24308: inst = 32'd268468224;
      24309: inst = 32'd201349021;
      24310: inst = 32'd203457618;
      24311: inst = 32'd136314880;
      24312: inst = 32'd268468224;
      24313: inst = 32'd201349022;
      24314: inst = 32'd203457651;
      24315: inst = 32'd136314880;
      24316: inst = 32'd268468224;
      24317: inst = 32'd201349023;
      24318: inst = 32'd203457618;
      24319: inst = 32'd136314880;
      24320: inst = 32'd268468224;
      24321: inst = 32'd201349024;
      24322: inst = 32'd203459696;
      24323: inst = 32'd136314880;
      24324: inst = 32'd268468224;
      24325: inst = 32'd201349025;
      24326: inst = 32'd203459696;
      24327: inst = 32'd136314880;
      24328: inst = 32'd268468224;
      24329: inst = 32'd201349026;
      24330: inst = 32'd203461777;
      24331: inst = 32'd136314880;
      24332: inst = 32'd268468224;
      24333: inst = 32'd201349027;
      24334: inst = 32'd203459697;
      24335: inst = 32'd136314880;
      24336: inst = 32'd268468224;
      24337: inst = 32'd201349028;
      24338: inst = 32'd203459665;
      24339: inst = 32'd136314880;
      24340: inst = 32'd268468224;
      24341: inst = 32'd201349029;
      24342: inst = 32'd203461779;
      24343: inst = 32'd136314880;
      24344: inst = 32'd268468224;
      24345: inst = 32'd201349030;
      24346: inst = 32'd203459633;
      24347: inst = 32'd136314880;
      24348: inst = 32'd268468224;
      24349: inst = 32'd201349031;
      24350: inst = 32'd203447021;
      24351: inst = 32'd136314880;
      24352: inst = 32'd268468224;
      24353: inst = 32'd201349032;
      24354: inst = 32'd203444875;
      24355: inst = 32'd136314880;
      24356: inst = 32'd268468224;
      24357: inst = 32'd201349033;
      24358: inst = 32'd203442796;
      24359: inst = 32'd136314880;
      24360: inst = 32'd268468224;
      24361: inst = 32'd201349034;
      24362: inst = 32'd203451248;
      24363: inst = 32'd136314880;
      24364: inst = 32'd268468224;
      24365: inst = 32'd201349035;
      24366: inst = 32'd203449167;
      24367: inst = 32'd136314880;
      24368: inst = 32'd268468224;
      24369: inst = 32'd201349036;
      24370: inst = 32'd203449200;
      24371: inst = 32'd136314880;
      24372: inst = 32'd268468224;
      24373: inst = 32'd201349037;
      24374: inst = 32'd203449200;
      24375: inst = 32'd136314880;
      24376: inst = 32'd268468224;
      24377: inst = 32'd201349038;
      24378: inst = 32'd203449200;
      24379: inst = 32'd136314880;
      24380: inst = 32'd268468224;
      24381: inst = 32'd201349039;
      24382: inst = 32'd203447152;
      24383: inst = 32'd136314880;
      24384: inst = 32'd268468224;
      24385: inst = 32'd201349040;
      24386: inst = 32'd203447152;
      24387: inst = 32'd136314880;
      24388: inst = 32'd268468224;
      24389: inst = 32'd201349041;
      24390: inst = 32'd203449200;
      24391: inst = 32'd136314880;
      24392: inst = 32'd268468224;
      24393: inst = 32'd201349042;
      24394: inst = 32'd203449200;
      24395: inst = 32'd136314880;
      24396: inst = 32'd268468224;
      24397: inst = 32'd201349043;
      24398: inst = 32'd203449200;
      24399: inst = 32'd136314880;
      24400: inst = 32'd268468224;
      24401: inst = 32'd201349044;
      24402: inst = 32'd203449167;
      24403: inst = 32'd136314880;
      24404: inst = 32'd268468224;
      24405: inst = 32'd201349045;
      24406: inst = 32'd203451248;
      24407: inst = 32'd136314880;
      24408: inst = 32'd268468224;
      24409: inst = 32'd201349046;
      24410: inst = 32'd203442796;
      24411: inst = 32'd136314880;
      24412: inst = 32'd268468224;
      24413: inst = 32'd201349047;
      24414: inst = 32'd203444875;
      24415: inst = 32'd136314880;
      24416: inst = 32'd268468224;
      24417: inst = 32'd201349048;
      24418: inst = 32'd203449069;
      24419: inst = 32'd136314880;
      24420: inst = 32'd268468224;
      24421: inst = 32'd201349049;
      24422: inst = 32'd203457585;
      24423: inst = 32'd136314880;
      24424: inst = 32'd268468224;
      24425: inst = 32'd201349050;
      24426: inst = 32'd203461778;
      24427: inst = 32'd136314880;
      24428: inst = 32'd268468224;
      24429: inst = 32'd201349051;
      24430: inst = 32'd203459665;
      24431: inst = 32'd136314880;
      24432: inst = 32'd268468224;
      24433: inst = 32'd201349052;
      24434: inst = 32'd203459697;
      24435: inst = 32'd136314880;
      24436: inst = 32'd268468224;
      24437: inst = 32'd201349053;
      24438: inst = 32'd203459697;
      24439: inst = 32'd136314880;
      24440: inst = 32'd268468224;
      24441: inst = 32'd201349054;
      24442: inst = 32'd203459664;
      24443: inst = 32'd136314880;
      24444: inst = 32'd268468224;
      24445: inst = 32'd201349055;
      24446: inst = 32'd203459697;
      24447: inst = 32'd136314880;
      24448: inst = 32'd268468224;
      24449: inst = 32'd201349056;
      24450: inst = 32'd203459664;
      24451: inst = 32'd136314880;
      24452: inst = 32'd268468224;
      24453: inst = 32'd201349057;
      24454: inst = 32'd203459697;
      24455: inst = 32'd136314880;
      24456: inst = 32'd268468224;
      24457: inst = 32'd201349058;
      24458: inst = 32'd203459664;
      24459: inst = 32'd136314880;
      24460: inst = 32'd268468224;
      24461: inst = 32'd201349059;
      24462: inst = 32'd203461777;
      24463: inst = 32'd136314880;
      24464: inst = 32'd268468224;
      24465: inst = 32'd201349060;
      24466: inst = 32'd203457649;
      24467: inst = 32'd136314880;
      24468: inst = 32'd268468224;
      24469: inst = 32'd201349061;
      24470: inst = 32'd203459729;
      24471: inst = 32'd136314880;
      24472: inst = 32'd268468224;
      24473: inst = 32'd201349062;
      24474: inst = 32'd203459697;
      24475: inst = 32'd136314880;
      24476: inst = 32'd268468224;
      24477: inst = 32'd201349063;
      24478: inst = 32'd203459729;
      24479: inst = 32'd136314880;
      24480: inst = 32'd268468224;
      24481: inst = 32'd201349064;
      24482: inst = 32'd203459697;
      24483: inst = 32'd136314880;
      24484: inst = 32'd268468224;
      24485: inst = 32'd201349065;
      24486: inst = 32'd203459697;
      24487: inst = 32'd136314880;
      24488: inst = 32'd268468224;
      24489: inst = 32'd201349066;
      24490: inst = 32'd203459729;
      24491: inst = 32'd136314880;
      24492: inst = 32'd268468224;
      24493: inst = 32'd201349067;
      24494: inst = 32'd203459730;
      24495: inst = 32'd136314880;
      24496: inst = 32'd268468224;
      24497: inst = 32'd201349068;
      24498: inst = 32'd203457618;
      24499: inst = 32'd136314880;
      24500: inst = 32'd268468224;
      24501: inst = 32'd201349069;
      24502: inst = 32'd203453457;
      24503: inst = 32'd136314880;
      24504: inst = 32'd268468224;
      24505: inst = 32'd201349070;
      24506: inst = 32'd203449264;
      24507: inst = 32'd136314880;
      24508: inst = 32'd268468224;
      24509: inst = 32'd201349071;
      24510: inst = 32'd203447151;
      24511: inst = 32'd136314880;
      24512: inst = 32'd268468224;
      24513: inst = 32'd201349072;
      24514: inst = 32'd203451215;
      24515: inst = 32'd136314880;
      24516: inst = 32'd268468224;
      24517: inst = 32'd201349073;
      24518: inst = 32'd203451215;
      24519: inst = 32'd136314880;
      24520: inst = 32'd268468224;
      24521: inst = 32'd201349074;
      24522: inst = 32'd203451215;
      24523: inst = 32'd136314880;
      24524: inst = 32'd268468224;
      24525: inst = 32'd201349075;
      24526: inst = 32'd203451215;
      24527: inst = 32'd136314880;
      24528: inst = 32'd268468224;
      24529: inst = 32'd201349076;
      24530: inst = 32'd203451215;
      24531: inst = 32'd136314880;
      24532: inst = 32'd268468224;
      24533: inst = 32'd201349077;
      24534: inst = 32'd203451215;
      24535: inst = 32'd136314880;
      24536: inst = 32'd268468224;
      24537: inst = 32'd201349078;
      24538: inst = 32'd203451215;
      24539: inst = 32'd136314880;
      24540: inst = 32'd268468224;
      24541: inst = 32'd201349079;
      24542: inst = 32'd203451215;
      24543: inst = 32'd136314880;
      24544: inst = 32'd268468224;
      24545: inst = 32'd201349080;
      24546: inst = 32'd203451215;
      24547: inst = 32'd136314880;
      24548: inst = 32'd268468224;
      24549: inst = 32'd201349081;
      24550: inst = 32'd203451215;
      24551: inst = 32'd136314880;
      24552: inst = 32'd268468224;
      24553: inst = 32'd201349082;
      24554: inst = 32'd203451215;
      24555: inst = 32'd136314880;
      24556: inst = 32'd268468224;
      24557: inst = 32'd201349083;
      24558: inst = 32'd203451215;
      24559: inst = 32'd136314880;
      24560: inst = 32'd268468224;
      24561: inst = 32'd201349084;
      24562: inst = 32'd203451215;
      24563: inst = 32'd136314880;
      24564: inst = 32'd268468224;
      24565: inst = 32'd201349085;
      24566: inst = 32'd203451215;
      24567: inst = 32'd136314880;
      24568: inst = 32'd268468224;
      24569: inst = 32'd201349086;
      24570: inst = 32'd203451215;
      24571: inst = 32'd136314880;
      24572: inst = 32'd268468224;
      24573: inst = 32'd201349087;
      24574: inst = 32'd203451215;
      24575: inst = 32'd136314880;
    endcase
  end
endmodule
