`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Company: lirc572
// Engineer: lirc572
// 
// Create Date: 
// Design Name: NECPU
// Module Name: InstMem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module instMem (
    input  [31:0]  address,
    output reg [31:0] inst
  );
  always @ (address) begin
    inst = 32'd0;
    case (address)
      0: inst = 32'h10000000;
      1: inst = 32'hc000005;
      2: inst = 32'h13e00000;
      3: inst = 32'hfe00087;
      4: inst = 32'h5be00000;
      5: inst = 32'h1020007f;
      6: inst = 32'hc202815;
      7: inst = 32'h30210001;
      8: inst = 32'h13e00000;
      9: inst = 32'hfe00007;
      10: inst = 32'h1c200000;
      11: inst = 32'h5be00000;
      12: inst = 32'h10000000;
      13: inst = 32'hc000011;
      14: inst = 32'h13e00000;
      15: inst = 32'hfe048df;
      16: inst = 32'h5be00000;
      17: inst = 32'h1020007f;
      18: inst = 32'hc202815;
      19: inst = 32'h30210001;
      20: inst = 32'h13e00000;
      21: inst = 32'hfe00013;
      22: inst = 32'h1c200000;
      23: inst = 32'h5be00000;
      24: inst = 32'h10000000;
      25: inst = 32'hc000000;
      26: inst = 32'h10200000;
      27: inst = 32'hc20001f;
      28: inst = 32'h13e00000;
      29: inst = 32'hfe060f8;
      30: inst = 32'h5be00000;
      31: inst = 32'h10000000;
      32: inst = 32'hc000024;
      33: inst = 32'h13a00000;
      34: inst = 32'hfa00000;
      35: inst = 32'h13600000;
      36: inst = 32'hf600000;
      37: inst = 32'h13800000;
      38: inst = 32'hf800000;
      39: inst = 32'h10208000;
      40: inst = 32'hc200001;
      41: inst = 32'h4210000;
      42: inst = 32'h10400000;
      43: inst = 32'hc40001b;
      44: inst = 32'h34211000;
      45: inst = 32'h38211000;
      46: inst = 32'h13e00000;
      47: inst = 32'hfe00041;
      48: inst = 32'h20200010;
      49: inst = 32'h5be00000;
      50: inst = 32'h13e00000;
      51: inst = 32'hfe0004b;
      52: inst = 32'h20200008;
      53: inst = 32'h5be00000;
      54: inst = 32'h13e00000;
      55: inst = 32'hfe00055;
      56: inst = 32'h20200004;
      57: inst = 32'h5be00000;
      58: inst = 32'h13e00000;
      59: inst = 32'hfe0005f;
      60: inst = 32'h20200002;
      61: inst = 32'h5be00000;
      62: inst = 32'h13e00000;
      63: inst = 32'hfe00069;
      64: inst = 32'h5be00000;
      65: inst = 32'h339c0001;
      66: inst = 32'h13a00000;
      67: inst = 32'hfa00000;
      68: inst = 32'hca00001;
      69: inst = 32'h10c08000;
      70: inst = 32'hcc00000;
      71: inst = 32'h8a60000;
      72: inst = 32'h13e00000;
      73: inst = 32'hfe0006d;
      74: inst = 32'h5be00000;
      75: inst = 32'h2b7b0001;
      76: inst = 32'h13a00000;
      77: inst = 32'hfa00003;
      78: inst = 32'hca00002;
      79: inst = 32'h10c08000;
      80: inst = 32'hcc00000;
      81: inst = 32'h8a60000;
      82: inst = 32'h13e00000;
      83: inst = 32'hfe0006d;
      84: inst = 32'h5be00000;
      85: inst = 32'h337b0001;
      86: inst = 32'h13a00000;
      87: inst = 32'hfa00001;
      88: inst = 32'hca00004;
      89: inst = 32'h10c08000;
      90: inst = 32'hcc00000;
      91: inst = 32'h8a60000;
      92: inst = 32'h13e00000;
      93: inst = 32'hfe0006d;
      94: inst = 32'h5be00000;
      95: inst = 32'h2b9c0001;
      96: inst = 32'h13a00000;
      97: inst = 32'hfa00005;
      98: inst = 32'hca00008;
      99: inst = 32'h10c08000;
      100: inst = 32'hcc00000;
      101: inst = 32'h8a60000;
      102: inst = 32'h13e00000;
      103: inst = 32'hfe0006d;
      104: inst = 32'h5be00000;
      105: inst = 32'hca00010;
      106: inst = 32'h10c08000;
      107: inst = 32'hcc00000;
      108: inst = 32'h8a60000;
      109: inst = 32'h10000000;
      110: inst = 32'hc000072;
      111: inst = 32'h13e00000;
      112: inst = 32'hfe06102;
      113: inst = 32'h5be00000;
      114: inst = 32'h283d0000;
      115: inst = 32'h285b0000;
      116: inst = 32'h287c0000;
      117: inst = 32'h10000000;
      118: inst = 32'hc00007a;
      119: inst = 32'h13e00000;
      120: inst = 32'hfe05130;
      121: inst = 32'h5be00000;
      122: inst = 32'h10200002;
      123: inst = 32'hc208b0a;
      124: inst = 32'h30210001;
      125: inst = 32'h13e00000;
      126: inst = 32'hfe0007c;
      127: inst = 32'h1c200000;
      128: inst = 32'h5be00000;
      129: inst = 32'h13e00000;
      130: inst = 32'hfe00027;
      131: inst = 32'h5be00000;
      132: inst = 32'h13e00000;
      133: inst = 32'hfe0a9f4;
      134: inst = 32'h5be00000;
      135: inst = 32'hc20eeb6;
      136: inst = 32'h10408000;
      137: inst = 32'hc403fe0;
      138: inst = 32'h8220000;
      139: inst = 32'h10408000;
      140: inst = 32'hc403fe1;
      141: inst = 32'h8220000;
      142: inst = 32'h10408000;
      143: inst = 32'hc403fe2;
      144: inst = 32'h8220000;
      145: inst = 32'h10408000;
      146: inst = 32'hc403fe3;
      147: inst = 32'h8220000;
      148: inst = 32'h10408000;
      149: inst = 32'hc403fe4;
      150: inst = 32'h8220000;
      151: inst = 32'h10408000;
      152: inst = 32'hc403fe5;
      153: inst = 32'h8220000;
      154: inst = 32'h10408000;
      155: inst = 32'hc403fe6;
      156: inst = 32'h8220000;
      157: inst = 32'h10408000;
      158: inst = 32'hc403fe7;
      159: inst = 32'h8220000;
      160: inst = 32'h10408000;
      161: inst = 32'hc403fe8;
      162: inst = 32'h8220000;
      163: inst = 32'h10408000;
      164: inst = 32'hc403fe9;
      165: inst = 32'h8220000;
      166: inst = 32'h10408000;
      167: inst = 32'hc403fea;
      168: inst = 32'h8220000;
      169: inst = 32'h10408000;
      170: inst = 32'hc403fec;
      171: inst = 32'h8220000;
      172: inst = 32'h10408000;
      173: inst = 32'hc403fed;
      174: inst = 32'h8220000;
      175: inst = 32'h10408000;
      176: inst = 32'hc403fee;
      177: inst = 32'h8220000;
      178: inst = 32'h10408000;
      179: inst = 32'hc403fef;
      180: inst = 32'h8220000;
      181: inst = 32'h10408000;
      182: inst = 32'hc403ff0;
      183: inst = 32'h8220000;
      184: inst = 32'h10408000;
      185: inst = 32'hc403ff1;
      186: inst = 32'h8220000;
      187: inst = 32'h10408000;
      188: inst = 32'hc403ff2;
      189: inst = 32'h8220000;
      190: inst = 32'h10408000;
      191: inst = 32'hc403ff3;
      192: inst = 32'h8220000;
      193: inst = 32'h10408000;
      194: inst = 32'hc403ff4;
      195: inst = 32'h8220000;
      196: inst = 32'h10408000;
      197: inst = 32'hc403ff5;
      198: inst = 32'h8220000;
      199: inst = 32'h10408000;
      200: inst = 32'hc403ff6;
      201: inst = 32'h8220000;
      202: inst = 32'h10408000;
      203: inst = 32'hc403ff7;
      204: inst = 32'h8220000;
      205: inst = 32'h10408000;
      206: inst = 32'hc403ff8;
      207: inst = 32'h8220000;
      208: inst = 32'h10408000;
      209: inst = 32'hc403ff9;
      210: inst = 32'h8220000;
      211: inst = 32'h10408000;
      212: inst = 32'hc403ffa;
      213: inst = 32'h8220000;
      214: inst = 32'h10408000;
      215: inst = 32'hc403ffb;
      216: inst = 32'h8220000;
      217: inst = 32'h10408000;
      218: inst = 32'hc403ffc;
      219: inst = 32'h8220000;
      220: inst = 32'h10408000;
      221: inst = 32'hc403ffd;
      222: inst = 32'h8220000;
      223: inst = 32'h10408000;
      224: inst = 32'hc403ffe;
      225: inst = 32'h8220000;
      226: inst = 32'h10408000;
      227: inst = 32'hc403fff;
      228: inst = 32'h8220000;
      229: inst = 32'h10408000;
      230: inst = 32'hc404000;
      231: inst = 32'h8220000;
      232: inst = 32'h10408000;
      233: inst = 32'hc404001;
      234: inst = 32'h8220000;
      235: inst = 32'h10408000;
      236: inst = 32'hc404002;
      237: inst = 32'h8220000;
      238: inst = 32'h10408000;
      239: inst = 32'hc404003;
      240: inst = 32'h8220000;
      241: inst = 32'h10408000;
      242: inst = 32'hc404004;
      243: inst = 32'h8220000;
      244: inst = 32'h10408000;
      245: inst = 32'hc404005;
      246: inst = 32'h8220000;
      247: inst = 32'h10408000;
      248: inst = 32'hc404006;
      249: inst = 32'h8220000;
      250: inst = 32'h10408000;
      251: inst = 32'hc404007;
      252: inst = 32'h8220000;
      253: inst = 32'h10408000;
      254: inst = 32'hc404008;
      255: inst = 32'h8220000;
      256: inst = 32'h10408000;
      257: inst = 32'hc404009;
      258: inst = 32'h8220000;
      259: inst = 32'h10408000;
      260: inst = 32'hc40400a;
      261: inst = 32'h8220000;
      262: inst = 32'h10408000;
      263: inst = 32'hc40400b;
      264: inst = 32'h8220000;
      265: inst = 32'h10408000;
      266: inst = 32'hc40400c;
      267: inst = 32'h8220000;
      268: inst = 32'h10408000;
      269: inst = 32'hc40400d;
      270: inst = 32'h8220000;
      271: inst = 32'h10408000;
      272: inst = 32'hc40400e;
      273: inst = 32'h8220000;
      274: inst = 32'h10408000;
      275: inst = 32'hc40400f;
      276: inst = 32'h8220000;
      277: inst = 32'h10408000;
      278: inst = 32'hc404010;
      279: inst = 32'h8220000;
      280: inst = 32'h10408000;
      281: inst = 32'hc404011;
      282: inst = 32'h8220000;
      283: inst = 32'h10408000;
      284: inst = 32'hc404012;
      285: inst = 32'h8220000;
      286: inst = 32'h10408000;
      287: inst = 32'hc404013;
      288: inst = 32'h8220000;
      289: inst = 32'h10408000;
      290: inst = 32'hc404014;
      291: inst = 32'h8220000;
      292: inst = 32'h10408000;
      293: inst = 32'hc404015;
      294: inst = 32'h8220000;
      295: inst = 32'h10408000;
      296: inst = 32'hc404016;
      297: inst = 32'h8220000;
      298: inst = 32'h10408000;
      299: inst = 32'hc404017;
      300: inst = 32'h8220000;
      301: inst = 32'h10408000;
      302: inst = 32'hc404018;
      303: inst = 32'h8220000;
      304: inst = 32'h10408000;
      305: inst = 32'hc404019;
      306: inst = 32'h8220000;
      307: inst = 32'h10408000;
      308: inst = 32'hc40401a;
      309: inst = 32'h8220000;
      310: inst = 32'h10408000;
      311: inst = 32'hc40401b;
      312: inst = 32'h8220000;
      313: inst = 32'h10408000;
      314: inst = 32'hc40401c;
      315: inst = 32'h8220000;
      316: inst = 32'h10408000;
      317: inst = 32'hc40401d;
      318: inst = 32'h8220000;
      319: inst = 32'h10408000;
      320: inst = 32'hc40401e;
      321: inst = 32'h8220000;
      322: inst = 32'h10408000;
      323: inst = 32'hc40401f;
      324: inst = 32'h8220000;
      325: inst = 32'h10408000;
      326: inst = 32'hc404020;
      327: inst = 32'h8220000;
      328: inst = 32'h10408000;
      329: inst = 32'hc404021;
      330: inst = 32'h8220000;
      331: inst = 32'h10408000;
      332: inst = 32'hc404022;
      333: inst = 32'h8220000;
      334: inst = 32'h10408000;
      335: inst = 32'hc404023;
      336: inst = 32'h8220000;
      337: inst = 32'h10408000;
      338: inst = 32'hc404024;
      339: inst = 32'h8220000;
      340: inst = 32'h10408000;
      341: inst = 32'hc404025;
      342: inst = 32'h8220000;
      343: inst = 32'h10408000;
      344: inst = 32'hc404026;
      345: inst = 32'h8220000;
      346: inst = 32'h10408000;
      347: inst = 32'hc404027;
      348: inst = 32'h8220000;
      349: inst = 32'h10408000;
      350: inst = 32'hc404028;
      351: inst = 32'h8220000;
      352: inst = 32'h10408000;
      353: inst = 32'hc404029;
      354: inst = 32'h8220000;
      355: inst = 32'h10408000;
      356: inst = 32'hc40402a;
      357: inst = 32'h8220000;
      358: inst = 32'h10408000;
      359: inst = 32'hc40402b;
      360: inst = 32'h8220000;
      361: inst = 32'h10408000;
      362: inst = 32'hc40402c;
      363: inst = 32'h8220000;
      364: inst = 32'h10408000;
      365: inst = 32'hc40402d;
      366: inst = 32'h8220000;
      367: inst = 32'h10408000;
      368: inst = 32'hc40402e;
      369: inst = 32'h8220000;
      370: inst = 32'h10408000;
      371: inst = 32'hc40402f;
      372: inst = 32'h8220000;
      373: inst = 32'h10408000;
      374: inst = 32'hc404030;
      375: inst = 32'h8220000;
      376: inst = 32'h10408000;
      377: inst = 32'hc404031;
      378: inst = 32'h8220000;
      379: inst = 32'h10408000;
      380: inst = 32'hc404032;
      381: inst = 32'h8220000;
      382: inst = 32'h10408000;
      383: inst = 32'hc404033;
      384: inst = 32'h8220000;
      385: inst = 32'h10408000;
      386: inst = 32'hc404034;
      387: inst = 32'h8220000;
      388: inst = 32'h10408000;
      389: inst = 32'hc404035;
      390: inst = 32'h8220000;
      391: inst = 32'h10408000;
      392: inst = 32'hc404036;
      393: inst = 32'h8220000;
      394: inst = 32'h10408000;
      395: inst = 32'hc404037;
      396: inst = 32'h8220000;
      397: inst = 32'h10408000;
      398: inst = 32'hc404038;
      399: inst = 32'h8220000;
      400: inst = 32'h10408000;
      401: inst = 32'hc404039;
      402: inst = 32'h8220000;
      403: inst = 32'h10408000;
      404: inst = 32'hc40403a;
      405: inst = 32'h8220000;
      406: inst = 32'h10408000;
      407: inst = 32'hc40403b;
      408: inst = 32'h8220000;
      409: inst = 32'h10408000;
      410: inst = 32'hc40403c;
      411: inst = 32'h8220000;
      412: inst = 32'h10408000;
      413: inst = 32'hc40403d;
      414: inst = 32'h8220000;
      415: inst = 32'h10408000;
      416: inst = 32'hc40403e;
      417: inst = 32'h8220000;
      418: inst = 32'h10408000;
      419: inst = 32'hc40403f;
      420: inst = 32'h8220000;
      421: inst = 32'h10408000;
      422: inst = 32'hc404040;
      423: inst = 32'h8220000;
      424: inst = 32'h10408000;
      425: inst = 32'hc404041;
      426: inst = 32'h8220000;
      427: inst = 32'h10408000;
      428: inst = 32'hc404042;
      429: inst = 32'h8220000;
      430: inst = 32'h10408000;
      431: inst = 32'hc404043;
      432: inst = 32'h8220000;
      433: inst = 32'h10408000;
      434: inst = 32'hc404044;
      435: inst = 32'h8220000;
      436: inst = 32'h10408000;
      437: inst = 32'hc404045;
      438: inst = 32'h8220000;
      439: inst = 32'h10408000;
      440: inst = 32'hc404046;
      441: inst = 32'h8220000;
      442: inst = 32'h10408000;
      443: inst = 32'hc404047;
      444: inst = 32'h8220000;
      445: inst = 32'h10408000;
      446: inst = 32'hc404048;
      447: inst = 32'h8220000;
      448: inst = 32'h10408000;
      449: inst = 32'hc404049;
      450: inst = 32'h8220000;
      451: inst = 32'h10408000;
      452: inst = 32'hc40404a;
      453: inst = 32'h8220000;
      454: inst = 32'h10408000;
      455: inst = 32'hc40404c;
      456: inst = 32'h8220000;
      457: inst = 32'h10408000;
      458: inst = 32'hc40404d;
      459: inst = 32'h8220000;
      460: inst = 32'h10408000;
      461: inst = 32'hc40404e;
      462: inst = 32'h8220000;
      463: inst = 32'h10408000;
      464: inst = 32'hc40404f;
      465: inst = 32'h8220000;
      466: inst = 32'h10408000;
      467: inst = 32'hc404050;
      468: inst = 32'h8220000;
      469: inst = 32'h10408000;
      470: inst = 32'hc404051;
      471: inst = 32'h8220000;
      472: inst = 32'h10408000;
      473: inst = 32'hc404052;
      474: inst = 32'h8220000;
      475: inst = 32'h10408000;
      476: inst = 32'hc404053;
      477: inst = 32'h8220000;
      478: inst = 32'h10408000;
      479: inst = 32'hc404054;
      480: inst = 32'h8220000;
      481: inst = 32'h10408000;
      482: inst = 32'hc404055;
      483: inst = 32'h8220000;
      484: inst = 32'h10408000;
      485: inst = 32'hc404056;
      486: inst = 32'h8220000;
      487: inst = 32'h10408000;
      488: inst = 32'hc404057;
      489: inst = 32'h8220000;
      490: inst = 32'h10408000;
      491: inst = 32'hc404058;
      492: inst = 32'h8220000;
      493: inst = 32'h10408000;
      494: inst = 32'hc404059;
      495: inst = 32'h8220000;
      496: inst = 32'h10408000;
      497: inst = 32'hc40405a;
      498: inst = 32'h8220000;
      499: inst = 32'h10408000;
      500: inst = 32'hc40405b;
      501: inst = 32'h8220000;
      502: inst = 32'h10408000;
      503: inst = 32'hc40405c;
      504: inst = 32'h8220000;
      505: inst = 32'h10408000;
      506: inst = 32'hc40405d;
      507: inst = 32'h8220000;
      508: inst = 32'h10408000;
      509: inst = 32'hc40405e;
      510: inst = 32'h8220000;
      511: inst = 32'h10408000;
      512: inst = 32'hc40405f;
      513: inst = 32'h8220000;
      514: inst = 32'h10408000;
      515: inst = 32'hc404060;
      516: inst = 32'h8220000;
      517: inst = 32'h10408000;
      518: inst = 32'hc404061;
      519: inst = 32'h8220000;
      520: inst = 32'h10408000;
      521: inst = 32'hc404062;
      522: inst = 32'h8220000;
      523: inst = 32'h10408000;
      524: inst = 32'hc404063;
      525: inst = 32'h8220000;
      526: inst = 32'h10408000;
      527: inst = 32'hc404064;
      528: inst = 32'h8220000;
      529: inst = 32'h10408000;
      530: inst = 32'hc404065;
      531: inst = 32'h8220000;
      532: inst = 32'h10408000;
      533: inst = 32'hc404066;
      534: inst = 32'h8220000;
      535: inst = 32'h10408000;
      536: inst = 32'hc404067;
      537: inst = 32'h8220000;
      538: inst = 32'h10408000;
      539: inst = 32'hc404068;
      540: inst = 32'h8220000;
      541: inst = 32'h10408000;
      542: inst = 32'hc404069;
      543: inst = 32'h8220000;
      544: inst = 32'h10408000;
      545: inst = 32'hc40406a;
      546: inst = 32'h8220000;
      547: inst = 32'h10408000;
      548: inst = 32'hc40406b;
      549: inst = 32'h8220000;
      550: inst = 32'h10408000;
      551: inst = 32'hc40406c;
      552: inst = 32'h8220000;
      553: inst = 32'h10408000;
      554: inst = 32'hc40406d;
      555: inst = 32'h8220000;
      556: inst = 32'h10408000;
      557: inst = 32'hc40406e;
      558: inst = 32'h8220000;
      559: inst = 32'h10408000;
      560: inst = 32'hc40406f;
      561: inst = 32'h8220000;
      562: inst = 32'h10408000;
      563: inst = 32'hc404070;
      564: inst = 32'h8220000;
      565: inst = 32'h10408000;
      566: inst = 32'hc404071;
      567: inst = 32'h8220000;
      568: inst = 32'h10408000;
      569: inst = 32'hc404072;
      570: inst = 32'h8220000;
      571: inst = 32'h10408000;
      572: inst = 32'hc404073;
      573: inst = 32'h8220000;
      574: inst = 32'h10408000;
      575: inst = 32'hc404074;
      576: inst = 32'h8220000;
      577: inst = 32'h10408000;
      578: inst = 32'hc404075;
      579: inst = 32'h8220000;
      580: inst = 32'h10408000;
      581: inst = 32'hc404076;
      582: inst = 32'h8220000;
      583: inst = 32'h10408000;
      584: inst = 32'hc404077;
      585: inst = 32'h8220000;
      586: inst = 32'h10408000;
      587: inst = 32'hc404078;
      588: inst = 32'h8220000;
      589: inst = 32'h10408000;
      590: inst = 32'hc404079;
      591: inst = 32'h8220000;
      592: inst = 32'h10408000;
      593: inst = 32'hc40407a;
      594: inst = 32'h8220000;
      595: inst = 32'h10408000;
      596: inst = 32'hc40407b;
      597: inst = 32'h8220000;
      598: inst = 32'h10408000;
      599: inst = 32'hc40407c;
      600: inst = 32'h8220000;
      601: inst = 32'h10408000;
      602: inst = 32'hc40407d;
      603: inst = 32'h8220000;
      604: inst = 32'h10408000;
      605: inst = 32'hc40407e;
      606: inst = 32'h8220000;
      607: inst = 32'h10408000;
      608: inst = 32'hc40407f;
      609: inst = 32'h8220000;
      610: inst = 32'h10408000;
      611: inst = 32'hc404080;
      612: inst = 32'h8220000;
      613: inst = 32'h10408000;
      614: inst = 32'hc404081;
      615: inst = 32'h8220000;
      616: inst = 32'h10408000;
      617: inst = 32'hc404082;
      618: inst = 32'h8220000;
      619: inst = 32'h10408000;
      620: inst = 32'hc404083;
      621: inst = 32'h8220000;
      622: inst = 32'h10408000;
      623: inst = 32'hc404084;
      624: inst = 32'h8220000;
      625: inst = 32'h10408000;
      626: inst = 32'hc404085;
      627: inst = 32'h8220000;
      628: inst = 32'h10408000;
      629: inst = 32'hc404086;
      630: inst = 32'h8220000;
      631: inst = 32'h10408000;
      632: inst = 32'hc404087;
      633: inst = 32'h8220000;
      634: inst = 32'h10408000;
      635: inst = 32'hc404088;
      636: inst = 32'h8220000;
      637: inst = 32'h10408000;
      638: inst = 32'hc404089;
      639: inst = 32'h8220000;
      640: inst = 32'h10408000;
      641: inst = 32'hc40408a;
      642: inst = 32'h8220000;
      643: inst = 32'h10408000;
      644: inst = 32'hc40408b;
      645: inst = 32'h8220000;
      646: inst = 32'h10408000;
      647: inst = 32'hc40408c;
      648: inst = 32'h8220000;
      649: inst = 32'h10408000;
      650: inst = 32'hc40408d;
      651: inst = 32'h8220000;
      652: inst = 32'h10408000;
      653: inst = 32'hc40408e;
      654: inst = 32'h8220000;
      655: inst = 32'h10408000;
      656: inst = 32'hc40408f;
      657: inst = 32'h8220000;
      658: inst = 32'h10408000;
      659: inst = 32'hc404090;
      660: inst = 32'h8220000;
      661: inst = 32'h10408000;
      662: inst = 32'hc404091;
      663: inst = 32'h8220000;
      664: inst = 32'h10408000;
      665: inst = 32'hc404092;
      666: inst = 32'h8220000;
      667: inst = 32'h10408000;
      668: inst = 32'hc404093;
      669: inst = 32'h8220000;
      670: inst = 32'h10408000;
      671: inst = 32'hc404094;
      672: inst = 32'h8220000;
      673: inst = 32'h10408000;
      674: inst = 32'hc404095;
      675: inst = 32'h8220000;
      676: inst = 32'h10408000;
      677: inst = 32'hc404096;
      678: inst = 32'h8220000;
      679: inst = 32'h10408000;
      680: inst = 32'hc404097;
      681: inst = 32'h8220000;
      682: inst = 32'h10408000;
      683: inst = 32'hc404098;
      684: inst = 32'h8220000;
      685: inst = 32'h10408000;
      686: inst = 32'hc404099;
      687: inst = 32'h8220000;
      688: inst = 32'h10408000;
      689: inst = 32'hc40409a;
      690: inst = 32'h8220000;
      691: inst = 32'h10408000;
      692: inst = 32'hc40409b;
      693: inst = 32'h8220000;
      694: inst = 32'h10408000;
      695: inst = 32'hc40409c;
      696: inst = 32'h8220000;
      697: inst = 32'h10408000;
      698: inst = 32'hc40409d;
      699: inst = 32'h8220000;
      700: inst = 32'h10408000;
      701: inst = 32'hc40409e;
      702: inst = 32'h8220000;
      703: inst = 32'h10408000;
      704: inst = 32'hc40409f;
      705: inst = 32'h8220000;
      706: inst = 32'h10408000;
      707: inst = 32'hc4040a0;
      708: inst = 32'h8220000;
      709: inst = 32'h10408000;
      710: inst = 32'hc4040a1;
      711: inst = 32'h8220000;
      712: inst = 32'h10408000;
      713: inst = 32'hc4040a2;
      714: inst = 32'h8220000;
      715: inst = 32'h10408000;
      716: inst = 32'hc4040a3;
      717: inst = 32'h8220000;
      718: inst = 32'h10408000;
      719: inst = 32'hc4040a4;
      720: inst = 32'h8220000;
      721: inst = 32'h10408000;
      722: inst = 32'hc4040a5;
      723: inst = 32'h8220000;
      724: inst = 32'h10408000;
      725: inst = 32'hc4040a6;
      726: inst = 32'h8220000;
      727: inst = 32'h10408000;
      728: inst = 32'hc4040a7;
      729: inst = 32'h8220000;
      730: inst = 32'h10408000;
      731: inst = 32'hc4040a8;
      732: inst = 32'h8220000;
      733: inst = 32'h10408000;
      734: inst = 32'hc4040a9;
      735: inst = 32'h8220000;
      736: inst = 32'h10408000;
      737: inst = 32'hc4040aa;
      738: inst = 32'h8220000;
      739: inst = 32'h10408000;
      740: inst = 32'hc4040ac;
      741: inst = 32'h8220000;
      742: inst = 32'h10408000;
      743: inst = 32'hc4040ad;
      744: inst = 32'h8220000;
      745: inst = 32'h10408000;
      746: inst = 32'hc4040ae;
      747: inst = 32'h8220000;
      748: inst = 32'h10408000;
      749: inst = 32'hc4040af;
      750: inst = 32'h8220000;
      751: inst = 32'h10408000;
      752: inst = 32'hc4040b0;
      753: inst = 32'h8220000;
      754: inst = 32'h10408000;
      755: inst = 32'hc4040b1;
      756: inst = 32'h8220000;
      757: inst = 32'h10408000;
      758: inst = 32'hc4040b2;
      759: inst = 32'h8220000;
      760: inst = 32'h10408000;
      761: inst = 32'hc4040b3;
      762: inst = 32'h8220000;
      763: inst = 32'h10408000;
      764: inst = 32'hc4040b4;
      765: inst = 32'h8220000;
      766: inst = 32'h10408000;
      767: inst = 32'hc4040b5;
      768: inst = 32'h8220000;
      769: inst = 32'h10408000;
      770: inst = 32'hc4040b6;
      771: inst = 32'h8220000;
      772: inst = 32'h10408000;
      773: inst = 32'hc4040b7;
      774: inst = 32'h8220000;
      775: inst = 32'h10408000;
      776: inst = 32'hc4040b8;
      777: inst = 32'h8220000;
      778: inst = 32'h10408000;
      779: inst = 32'hc4040b9;
      780: inst = 32'h8220000;
      781: inst = 32'h10408000;
      782: inst = 32'hc4040ba;
      783: inst = 32'h8220000;
      784: inst = 32'h10408000;
      785: inst = 32'hc4040bb;
      786: inst = 32'h8220000;
      787: inst = 32'h10408000;
      788: inst = 32'hc4040bc;
      789: inst = 32'h8220000;
      790: inst = 32'h10408000;
      791: inst = 32'hc4040bd;
      792: inst = 32'h8220000;
      793: inst = 32'h10408000;
      794: inst = 32'hc4040be;
      795: inst = 32'h8220000;
      796: inst = 32'h10408000;
      797: inst = 32'hc4040bf;
      798: inst = 32'h8220000;
      799: inst = 32'h10408000;
      800: inst = 32'hc4040c0;
      801: inst = 32'h8220000;
      802: inst = 32'h10408000;
      803: inst = 32'hc4040c1;
      804: inst = 32'h8220000;
      805: inst = 32'h10408000;
      806: inst = 32'hc4040c2;
      807: inst = 32'h8220000;
      808: inst = 32'h10408000;
      809: inst = 32'hc4040c3;
      810: inst = 32'h8220000;
      811: inst = 32'h10408000;
      812: inst = 32'hc4040c4;
      813: inst = 32'h8220000;
      814: inst = 32'h10408000;
      815: inst = 32'hc4040c5;
      816: inst = 32'h8220000;
      817: inst = 32'h10408000;
      818: inst = 32'hc4040c6;
      819: inst = 32'h8220000;
      820: inst = 32'h10408000;
      821: inst = 32'hc4040c7;
      822: inst = 32'h8220000;
      823: inst = 32'h10408000;
      824: inst = 32'hc4040c8;
      825: inst = 32'h8220000;
      826: inst = 32'h10408000;
      827: inst = 32'hc4040c9;
      828: inst = 32'h8220000;
      829: inst = 32'h10408000;
      830: inst = 32'hc4040ca;
      831: inst = 32'h8220000;
      832: inst = 32'h10408000;
      833: inst = 32'hc4040cb;
      834: inst = 32'h8220000;
      835: inst = 32'h10408000;
      836: inst = 32'hc4040cc;
      837: inst = 32'h8220000;
      838: inst = 32'h10408000;
      839: inst = 32'hc4040cd;
      840: inst = 32'h8220000;
      841: inst = 32'h10408000;
      842: inst = 32'hc4040ce;
      843: inst = 32'h8220000;
      844: inst = 32'h10408000;
      845: inst = 32'hc4040cf;
      846: inst = 32'h8220000;
      847: inst = 32'h10408000;
      848: inst = 32'hc4040d0;
      849: inst = 32'h8220000;
      850: inst = 32'h10408000;
      851: inst = 32'hc4040d1;
      852: inst = 32'h8220000;
      853: inst = 32'h10408000;
      854: inst = 32'hc4040d2;
      855: inst = 32'h8220000;
      856: inst = 32'h10408000;
      857: inst = 32'hc4040d3;
      858: inst = 32'h8220000;
      859: inst = 32'h10408000;
      860: inst = 32'hc4040d4;
      861: inst = 32'h8220000;
      862: inst = 32'h10408000;
      863: inst = 32'hc4040d5;
      864: inst = 32'h8220000;
      865: inst = 32'h10408000;
      866: inst = 32'hc4040d6;
      867: inst = 32'h8220000;
      868: inst = 32'h10408000;
      869: inst = 32'hc4040d7;
      870: inst = 32'h8220000;
      871: inst = 32'h10408000;
      872: inst = 32'hc4040d8;
      873: inst = 32'h8220000;
      874: inst = 32'h10408000;
      875: inst = 32'hc4040d9;
      876: inst = 32'h8220000;
      877: inst = 32'h10408000;
      878: inst = 32'hc4040da;
      879: inst = 32'h8220000;
      880: inst = 32'h10408000;
      881: inst = 32'hc4040db;
      882: inst = 32'h8220000;
      883: inst = 32'h10408000;
      884: inst = 32'hc4040dc;
      885: inst = 32'h8220000;
      886: inst = 32'h10408000;
      887: inst = 32'hc4040dd;
      888: inst = 32'h8220000;
      889: inst = 32'h10408000;
      890: inst = 32'hc4040de;
      891: inst = 32'h8220000;
      892: inst = 32'h10408000;
      893: inst = 32'hc4040df;
      894: inst = 32'h8220000;
      895: inst = 32'h10408000;
      896: inst = 32'hc4040e0;
      897: inst = 32'h8220000;
      898: inst = 32'h10408000;
      899: inst = 32'hc4040e1;
      900: inst = 32'h8220000;
      901: inst = 32'h10408000;
      902: inst = 32'hc4040e2;
      903: inst = 32'h8220000;
      904: inst = 32'h10408000;
      905: inst = 32'hc4040e3;
      906: inst = 32'h8220000;
      907: inst = 32'h10408000;
      908: inst = 32'hc4040e4;
      909: inst = 32'h8220000;
      910: inst = 32'h10408000;
      911: inst = 32'hc4040e5;
      912: inst = 32'h8220000;
      913: inst = 32'h10408000;
      914: inst = 32'hc4040e6;
      915: inst = 32'h8220000;
      916: inst = 32'h10408000;
      917: inst = 32'hc4040e7;
      918: inst = 32'h8220000;
      919: inst = 32'h10408000;
      920: inst = 32'hc4040e8;
      921: inst = 32'h8220000;
      922: inst = 32'h10408000;
      923: inst = 32'hc4040e9;
      924: inst = 32'h8220000;
      925: inst = 32'h10408000;
      926: inst = 32'hc4040ea;
      927: inst = 32'h8220000;
      928: inst = 32'h10408000;
      929: inst = 32'hc4040eb;
      930: inst = 32'h8220000;
      931: inst = 32'h10408000;
      932: inst = 32'hc4040ec;
      933: inst = 32'h8220000;
      934: inst = 32'h10408000;
      935: inst = 32'hc4040ed;
      936: inst = 32'h8220000;
      937: inst = 32'h10408000;
      938: inst = 32'hc4040ee;
      939: inst = 32'h8220000;
      940: inst = 32'h10408000;
      941: inst = 32'hc4040ef;
      942: inst = 32'h8220000;
      943: inst = 32'h10408000;
      944: inst = 32'hc4040f0;
      945: inst = 32'h8220000;
      946: inst = 32'h10408000;
      947: inst = 32'hc4040f1;
      948: inst = 32'h8220000;
      949: inst = 32'h10408000;
      950: inst = 32'hc4040f2;
      951: inst = 32'h8220000;
      952: inst = 32'h10408000;
      953: inst = 32'hc4040f3;
      954: inst = 32'h8220000;
      955: inst = 32'h10408000;
      956: inst = 32'hc4040f4;
      957: inst = 32'h8220000;
      958: inst = 32'h10408000;
      959: inst = 32'hc4040f5;
      960: inst = 32'h8220000;
      961: inst = 32'h10408000;
      962: inst = 32'hc4040f6;
      963: inst = 32'h8220000;
      964: inst = 32'h10408000;
      965: inst = 32'hc4040f7;
      966: inst = 32'h8220000;
      967: inst = 32'h10408000;
      968: inst = 32'hc4040f8;
      969: inst = 32'h8220000;
      970: inst = 32'h10408000;
      971: inst = 32'hc4040f9;
      972: inst = 32'h8220000;
      973: inst = 32'h10408000;
      974: inst = 32'hc4040fa;
      975: inst = 32'h8220000;
      976: inst = 32'h10408000;
      977: inst = 32'hc4040fb;
      978: inst = 32'h8220000;
      979: inst = 32'h10408000;
      980: inst = 32'hc4040fc;
      981: inst = 32'h8220000;
      982: inst = 32'h10408000;
      983: inst = 32'hc4040fd;
      984: inst = 32'h8220000;
      985: inst = 32'h10408000;
      986: inst = 32'hc4040fe;
      987: inst = 32'h8220000;
      988: inst = 32'h10408000;
      989: inst = 32'hc4040ff;
      990: inst = 32'h8220000;
      991: inst = 32'h10408000;
      992: inst = 32'hc404100;
      993: inst = 32'h8220000;
      994: inst = 32'h10408000;
      995: inst = 32'hc404101;
      996: inst = 32'h8220000;
      997: inst = 32'h10408000;
      998: inst = 32'hc404102;
      999: inst = 32'h8220000;
      1000: inst = 32'h10408000;
      1001: inst = 32'hc404103;
      1002: inst = 32'h8220000;
      1003: inst = 32'h10408000;
      1004: inst = 32'hc404104;
      1005: inst = 32'h8220000;
      1006: inst = 32'h10408000;
      1007: inst = 32'hc404105;
      1008: inst = 32'h8220000;
      1009: inst = 32'h10408000;
      1010: inst = 32'hc404106;
      1011: inst = 32'h8220000;
      1012: inst = 32'h10408000;
      1013: inst = 32'hc404107;
      1014: inst = 32'h8220000;
      1015: inst = 32'h10408000;
      1016: inst = 32'hc404108;
      1017: inst = 32'h8220000;
      1018: inst = 32'h10408000;
      1019: inst = 32'hc404109;
      1020: inst = 32'h8220000;
      1021: inst = 32'h10408000;
      1022: inst = 32'hc40410a;
      1023: inst = 32'h8220000;
      1024: inst = 32'h10408000;
      1025: inst = 32'hc40410c;
      1026: inst = 32'h8220000;
      1027: inst = 32'h10408000;
      1028: inst = 32'hc40410d;
      1029: inst = 32'h8220000;
      1030: inst = 32'h10408000;
      1031: inst = 32'hc40410e;
      1032: inst = 32'h8220000;
      1033: inst = 32'h10408000;
      1034: inst = 32'hc40410f;
      1035: inst = 32'h8220000;
      1036: inst = 32'h10408000;
      1037: inst = 32'hc404110;
      1038: inst = 32'h8220000;
      1039: inst = 32'h10408000;
      1040: inst = 32'hc404111;
      1041: inst = 32'h8220000;
      1042: inst = 32'h10408000;
      1043: inst = 32'hc404112;
      1044: inst = 32'h8220000;
      1045: inst = 32'h10408000;
      1046: inst = 32'hc404113;
      1047: inst = 32'h8220000;
      1048: inst = 32'h10408000;
      1049: inst = 32'hc404114;
      1050: inst = 32'h8220000;
      1051: inst = 32'h10408000;
      1052: inst = 32'hc404115;
      1053: inst = 32'h8220000;
      1054: inst = 32'h10408000;
      1055: inst = 32'hc404116;
      1056: inst = 32'h8220000;
      1057: inst = 32'h10408000;
      1058: inst = 32'hc404117;
      1059: inst = 32'h8220000;
      1060: inst = 32'h10408000;
      1061: inst = 32'hc404118;
      1062: inst = 32'h8220000;
      1063: inst = 32'h10408000;
      1064: inst = 32'hc404119;
      1065: inst = 32'h8220000;
      1066: inst = 32'h10408000;
      1067: inst = 32'hc40411a;
      1068: inst = 32'h8220000;
      1069: inst = 32'h10408000;
      1070: inst = 32'hc40411b;
      1071: inst = 32'h8220000;
      1072: inst = 32'h10408000;
      1073: inst = 32'hc40411c;
      1074: inst = 32'h8220000;
      1075: inst = 32'h10408000;
      1076: inst = 32'hc40411d;
      1077: inst = 32'h8220000;
      1078: inst = 32'h10408000;
      1079: inst = 32'hc40411e;
      1080: inst = 32'h8220000;
      1081: inst = 32'h10408000;
      1082: inst = 32'hc40411f;
      1083: inst = 32'h8220000;
      1084: inst = 32'h10408000;
      1085: inst = 32'hc404120;
      1086: inst = 32'h8220000;
      1087: inst = 32'h10408000;
      1088: inst = 32'hc404121;
      1089: inst = 32'h8220000;
      1090: inst = 32'h10408000;
      1091: inst = 32'hc404122;
      1092: inst = 32'h8220000;
      1093: inst = 32'h10408000;
      1094: inst = 32'hc404123;
      1095: inst = 32'h8220000;
      1096: inst = 32'h10408000;
      1097: inst = 32'hc404124;
      1098: inst = 32'h8220000;
      1099: inst = 32'h10408000;
      1100: inst = 32'hc404125;
      1101: inst = 32'h8220000;
      1102: inst = 32'h10408000;
      1103: inst = 32'hc404126;
      1104: inst = 32'h8220000;
      1105: inst = 32'h10408000;
      1106: inst = 32'hc404127;
      1107: inst = 32'h8220000;
      1108: inst = 32'h10408000;
      1109: inst = 32'hc404128;
      1110: inst = 32'h8220000;
      1111: inst = 32'h10408000;
      1112: inst = 32'hc404129;
      1113: inst = 32'h8220000;
      1114: inst = 32'h10408000;
      1115: inst = 32'hc40412a;
      1116: inst = 32'h8220000;
      1117: inst = 32'h10408000;
      1118: inst = 32'hc40412b;
      1119: inst = 32'h8220000;
      1120: inst = 32'h10408000;
      1121: inst = 32'hc40412c;
      1122: inst = 32'h8220000;
      1123: inst = 32'h10408000;
      1124: inst = 32'hc40412d;
      1125: inst = 32'h8220000;
      1126: inst = 32'h10408000;
      1127: inst = 32'hc40412e;
      1128: inst = 32'h8220000;
      1129: inst = 32'h10408000;
      1130: inst = 32'hc40412f;
      1131: inst = 32'h8220000;
      1132: inst = 32'h10408000;
      1133: inst = 32'hc404130;
      1134: inst = 32'h8220000;
      1135: inst = 32'h10408000;
      1136: inst = 32'hc404131;
      1137: inst = 32'h8220000;
      1138: inst = 32'h10408000;
      1139: inst = 32'hc404132;
      1140: inst = 32'h8220000;
      1141: inst = 32'h10408000;
      1142: inst = 32'hc404133;
      1143: inst = 32'h8220000;
      1144: inst = 32'h10408000;
      1145: inst = 32'hc404134;
      1146: inst = 32'h8220000;
      1147: inst = 32'h10408000;
      1148: inst = 32'hc404135;
      1149: inst = 32'h8220000;
      1150: inst = 32'h10408000;
      1151: inst = 32'hc404136;
      1152: inst = 32'h8220000;
      1153: inst = 32'h10408000;
      1154: inst = 32'hc404137;
      1155: inst = 32'h8220000;
      1156: inst = 32'h10408000;
      1157: inst = 32'hc404138;
      1158: inst = 32'h8220000;
      1159: inst = 32'h10408000;
      1160: inst = 32'hc404139;
      1161: inst = 32'h8220000;
      1162: inst = 32'h10408000;
      1163: inst = 32'hc40413a;
      1164: inst = 32'h8220000;
      1165: inst = 32'h10408000;
      1166: inst = 32'hc40413b;
      1167: inst = 32'h8220000;
      1168: inst = 32'h10408000;
      1169: inst = 32'hc40413c;
      1170: inst = 32'h8220000;
      1171: inst = 32'h10408000;
      1172: inst = 32'hc40413d;
      1173: inst = 32'h8220000;
      1174: inst = 32'h10408000;
      1175: inst = 32'hc40413e;
      1176: inst = 32'h8220000;
      1177: inst = 32'h10408000;
      1178: inst = 32'hc40413f;
      1179: inst = 32'h8220000;
      1180: inst = 32'h10408000;
      1181: inst = 32'hc404140;
      1182: inst = 32'h8220000;
      1183: inst = 32'h10408000;
      1184: inst = 32'hc404141;
      1185: inst = 32'h8220000;
      1186: inst = 32'h10408000;
      1187: inst = 32'hc404142;
      1188: inst = 32'h8220000;
      1189: inst = 32'h10408000;
      1190: inst = 32'hc404143;
      1191: inst = 32'h8220000;
      1192: inst = 32'h10408000;
      1193: inst = 32'hc404144;
      1194: inst = 32'h8220000;
      1195: inst = 32'h10408000;
      1196: inst = 32'hc404145;
      1197: inst = 32'h8220000;
      1198: inst = 32'h10408000;
      1199: inst = 32'hc404146;
      1200: inst = 32'h8220000;
      1201: inst = 32'h10408000;
      1202: inst = 32'hc404147;
      1203: inst = 32'h8220000;
      1204: inst = 32'h10408000;
      1205: inst = 32'hc404148;
      1206: inst = 32'h8220000;
      1207: inst = 32'h10408000;
      1208: inst = 32'hc404149;
      1209: inst = 32'h8220000;
      1210: inst = 32'h10408000;
      1211: inst = 32'hc40414a;
      1212: inst = 32'h8220000;
      1213: inst = 32'h10408000;
      1214: inst = 32'hc40414b;
      1215: inst = 32'h8220000;
      1216: inst = 32'h10408000;
      1217: inst = 32'hc40414c;
      1218: inst = 32'h8220000;
      1219: inst = 32'h10408000;
      1220: inst = 32'hc40414d;
      1221: inst = 32'h8220000;
      1222: inst = 32'h10408000;
      1223: inst = 32'hc40414e;
      1224: inst = 32'h8220000;
      1225: inst = 32'h10408000;
      1226: inst = 32'hc40414f;
      1227: inst = 32'h8220000;
      1228: inst = 32'h10408000;
      1229: inst = 32'hc404150;
      1230: inst = 32'h8220000;
      1231: inst = 32'h10408000;
      1232: inst = 32'hc404151;
      1233: inst = 32'h8220000;
      1234: inst = 32'h10408000;
      1235: inst = 32'hc404152;
      1236: inst = 32'h8220000;
      1237: inst = 32'h10408000;
      1238: inst = 32'hc404153;
      1239: inst = 32'h8220000;
      1240: inst = 32'h10408000;
      1241: inst = 32'hc404154;
      1242: inst = 32'h8220000;
      1243: inst = 32'h10408000;
      1244: inst = 32'hc404155;
      1245: inst = 32'h8220000;
      1246: inst = 32'h10408000;
      1247: inst = 32'hc404156;
      1248: inst = 32'h8220000;
      1249: inst = 32'h10408000;
      1250: inst = 32'hc404157;
      1251: inst = 32'h8220000;
      1252: inst = 32'h10408000;
      1253: inst = 32'hc404158;
      1254: inst = 32'h8220000;
      1255: inst = 32'h10408000;
      1256: inst = 32'hc404159;
      1257: inst = 32'h8220000;
      1258: inst = 32'h10408000;
      1259: inst = 32'hc40415a;
      1260: inst = 32'h8220000;
      1261: inst = 32'h10408000;
      1262: inst = 32'hc40415b;
      1263: inst = 32'h8220000;
      1264: inst = 32'h10408000;
      1265: inst = 32'hc40415c;
      1266: inst = 32'h8220000;
      1267: inst = 32'h10408000;
      1268: inst = 32'hc40415d;
      1269: inst = 32'h8220000;
      1270: inst = 32'h10408000;
      1271: inst = 32'hc40415e;
      1272: inst = 32'h8220000;
      1273: inst = 32'h10408000;
      1274: inst = 32'hc40415f;
      1275: inst = 32'h8220000;
      1276: inst = 32'h10408000;
      1277: inst = 32'hc404160;
      1278: inst = 32'h8220000;
      1279: inst = 32'h10408000;
      1280: inst = 32'hc404161;
      1281: inst = 32'h8220000;
      1282: inst = 32'h10408000;
      1283: inst = 32'hc404162;
      1284: inst = 32'h8220000;
      1285: inst = 32'h10408000;
      1286: inst = 32'hc404163;
      1287: inst = 32'h8220000;
      1288: inst = 32'h10408000;
      1289: inst = 32'hc404164;
      1290: inst = 32'h8220000;
      1291: inst = 32'h10408000;
      1292: inst = 32'hc404165;
      1293: inst = 32'h8220000;
      1294: inst = 32'h10408000;
      1295: inst = 32'hc404166;
      1296: inst = 32'h8220000;
      1297: inst = 32'h10408000;
      1298: inst = 32'hc404167;
      1299: inst = 32'h8220000;
      1300: inst = 32'h10408000;
      1301: inst = 32'hc404168;
      1302: inst = 32'h8220000;
      1303: inst = 32'h10408000;
      1304: inst = 32'hc404169;
      1305: inst = 32'h8220000;
      1306: inst = 32'h10408000;
      1307: inst = 32'hc40416a;
      1308: inst = 32'h8220000;
      1309: inst = 32'h10408000;
      1310: inst = 32'hc40416c;
      1311: inst = 32'h8220000;
      1312: inst = 32'h10408000;
      1313: inst = 32'hc40416d;
      1314: inst = 32'h8220000;
      1315: inst = 32'h10408000;
      1316: inst = 32'hc40416e;
      1317: inst = 32'h8220000;
      1318: inst = 32'h10408000;
      1319: inst = 32'hc40416f;
      1320: inst = 32'h8220000;
      1321: inst = 32'h10408000;
      1322: inst = 32'hc404170;
      1323: inst = 32'h8220000;
      1324: inst = 32'h10408000;
      1325: inst = 32'hc404171;
      1326: inst = 32'h8220000;
      1327: inst = 32'h10408000;
      1328: inst = 32'hc404172;
      1329: inst = 32'h8220000;
      1330: inst = 32'h10408000;
      1331: inst = 32'hc404173;
      1332: inst = 32'h8220000;
      1333: inst = 32'h10408000;
      1334: inst = 32'hc404174;
      1335: inst = 32'h8220000;
      1336: inst = 32'h10408000;
      1337: inst = 32'hc404175;
      1338: inst = 32'h8220000;
      1339: inst = 32'h10408000;
      1340: inst = 32'hc404176;
      1341: inst = 32'h8220000;
      1342: inst = 32'h10408000;
      1343: inst = 32'hc404177;
      1344: inst = 32'h8220000;
      1345: inst = 32'h10408000;
      1346: inst = 32'hc404178;
      1347: inst = 32'h8220000;
      1348: inst = 32'h10408000;
      1349: inst = 32'hc404179;
      1350: inst = 32'h8220000;
      1351: inst = 32'h10408000;
      1352: inst = 32'hc40417a;
      1353: inst = 32'h8220000;
      1354: inst = 32'h10408000;
      1355: inst = 32'hc40417b;
      1356: inst = 32'h8220000;
      1357: inst = 32'h10408000;
      1358: inst = 32'hc40417c;
      1359: inst = 32'h8220000;
      1360: inst = 32'h10408000;
      1361: inst = 32'hc40417d;
      1362: inst = 32'h8220000;
      1363: inst = 32'h10408000;
      1364: inst = 32'hc40417e;
      1365: inst = 32'h8220000;
      1366: inst = 32'h10408000;
      1367: inst = 32'hc40417f;
      1368: inst = 32'h8220000;
      1369: inst = 32'h10408000;
      1370: inst = 32'hc404180;
      1371: inst = 32'h8220000;
      1372: inst = 32'h10408000;
      1373: inst = 32'hc404181;
      1374: inst = 32'h8220000;
      1375: inst = 32'h10408000;
      1376: inst = 32'hc404182;
      1377: inst = 32'h8220000;
      1378: inst = 32'h10408000;
      1379: inst = 32'hc404183;
      1380: inst = 32'h8220000;
      1381: inst = 32'h10408000;
      1382: inst = 32'hc404184;
      1383: inst = 32'h8220000;
      1384: inst = 32'h10408000;
      1385: inst = 32'hc404185;
      1386: inst = 32'h8220000;
      1387: inst = 32'h10408000;
      1388: inst = 32'hc404186;
      1389: inst = 32'h8220000;
      1390: inst = 32'h10408000;
      1391: inst = 32'hc404187;
      1392: inst = 32'h8220000;
      1393: inst = 32'h10408000;
      1394: inst = 32'hc404188;
      1395: inst = 32'h8220000;
      1396: inst = 32'h10408000;
      1397: inst = 32'hc404189;
      1398: inst = 32'h8220000;
      1399: inst = 32'h10408000;
      1400: inst = 32'hc40418a;
      1401: inst = 32'h8220000;
      1402: inst = 32'h10408000;
      1403: inst = 32'hc40418b;
      1404: inst = 32'h8220000;
      1405: inst = 32'h10408000;
      1406: inst = 32'hc40418c;
      1407: inst = 32'h8220000;
      1408: inst = 32'h10408000;
      1409: inst = 32'hc40418d;
      1410: inst = 32'h8220000;
      1411: inst = 32'h10408000;
      1412: inst = 32'hc40418e;
      1413: inst = 32'h8220000;
      1414: inst = 32'h10408000;
      1415: inst = 32'hc40418f;
      1416: inst = 32'h8220000;
      1417: inst = 32'h10408000;
      1418: inst = 32'hc404190;
      1419: inst = 32'h8220000;
      1420: inst = 32'h10408000;
      1421: inst = 32'hc404191;
      1422: inst = 32'h8220000;
      1423: inst = 32'h10408000;
      1424: inst = 32'hc404192;
      1425: inst = 32'h8220000;
      1426: inst = 32'h10408000;
      1427: inst = 32'hc404193;
      1428: inst = 32'h8220000;
      1429: inst = 32'h10408000;
      1430: inst = 32'hc404194;
      1431: inst = 32'h8220000;
      1432: inst = 32'h10408000;
      1433: inst = 32'hc404195;
      1434: inst = 32'h8220000;
      1435: inst = 32'h10408000;
      1436: inst = 32'hc404196;
      1437: inst = 32'h8220000;
      1438: inst = 32'h10408000;
      1439: inst = 32'hc404197;
      1440: inst = 32'h8220000;
      1441: inst = 32'h10408000;
      1442: inst = 32'hc404198;
      1443: inst = 32'h8220000;
      1444: inst = 32'h10408000;
      1445: inst = 32'hc404199;
      1446: inst = 32'h8220000;
      1447: inst = 32'h10408000;
      1448: inst = 32'hc40419a;
      1449: inst = 32'h8220000;
      1450: inst = 32'h10408000;
      1451: inst = 32'hc40419b;
      1452: inst = 32'h8220000;
      1453: inst = 32'h10408000;
      1454: inst = 32'hc40419c;
      1455: inst = 32'h8220000;
      1456: inst = 32'h10408000;
      1457: inst = 32'hc40419d;
      1458: inst = 32'h8220000;
      1459: inst = 32'h10408000;
      1460: inst = 32'hc40419e;
      1461: inst = 32'h8220000;
      1462: inst = 32'h10408000;
      1463: inst = 32'hc40419f;
      1464: inst = 32'h8220000;
      1465: inst = 32'h10408000;
      1466: inst = 32'hc4041a0;
      1467: inst = 32'h8220000;
      1468: inst = 32'h10408000;
      1469: inst = 32'hc4041a1;
      1470: inst = 32'h8220000;
      1471: inst = 32'h10408000;
      1472: inst = 32'hc4041a2;
      1473: inst = 32'h8220000;
      1474: inst = 32'h10408000;
      1475: inst = 32'hc4041a3;
      1476: inst = 32'h8220000;
      1477: inst = 32'h10408000;
      1478: inst = 32'hc4041a4;
      1479: inst = 32'h8220000;
      1480: inst = 32'h10408000;
      1481: inst = 32'hc4041a5;
      1482: inst = 32'h8220000;
      1483: inst = 32'h10408000;
      1484: inst = 32'hc4041a6;
      1485: inst = 32'h8220000;
      1486: inst = 32'h10408000;
      1487: inst = 32'hc4041a7;
      1488: inst = 32'h8220000;
      1489: inst = 32'h10408000;
      1490: inst = 32'hc4041a8;
      1491: inst = 32'h8220000;
      1492: inst = 32'h10408000;
      1493: inst = 32'hc4041a9;
      1494: inst = 32'h8220000;
      1495: inst = 32'h10408000;
      1496: inst = 32'hc4041aa;
      1497: inst = 32'h8220000;
      1498: inst = 32'h10408000;
      1499: inst = 32'hc4041ab;
      1500: inst = 32'h8220000;
      1501: inst = 32'h10408000;
      1502: inst = 32'hc4041ac;
      1503: inst = 32'h8220000;
      1504: inst = 32'h10408000;
      1505: inst = 32'hc4041ad;
      1506: inst = 32'h8220000;
      1507: inst = 32'h10408000;
      1508: inst = 32'hc4041ae;
      1509: inst = 32'h8220000;
      1510: inst = 32'h10408000;
      1511: inst = 32'hc4041af;
      1512: inst = 32'h8220000;
      1513: inst = 32'h10408000;
      1514: inst = 32'hc4041b0;
      1515: inst = 32'h8220000;
      1516: inst = 32'h10408000;
      1517: inst = 32'hc4041b1;
      1518: inst = 32'h8220000;
      1519: inst = 32'h10408000;
      1520: inst = 32'hc4041b2;
      1521: inst = 32'h8220000;
      1522: inst = 32'h10408000;
      1523: inst = 32'hc4041b3;
      1524: inst = 32'h8220000;
      1525: inst = 32'h10408000;
      1526: inst = 32'hc4041b4;
      1527: inst = 32'h8220000;
      1528: inst = 32'h10408000;
      1529: inst = 32'hc4041b5;
      1530: inst = 32'h8220000;
      1531: inst = 32'h10408000;
      1532: inst = 32'hc4041b6;
      1533: inst = 32'h8220000;
      1534: inst = 32'h10408000;
      1535: inst = 32'hc4041b7;
      1536: inst = 32'h8220000;
      1537: inst = 32'h10408000;
      1538: inst = 32'hc4041b8;
      1539: inst = 32'h8220000;
      1540: inst = 32'h10408000;
      1541: inst = 32'hc4041b9;
      1542: inst = 32'h8220000;
      1543: inst = 32'h10408000;
      1544: inst = 32'hc4041ba;
      1545: inst = 32'h8220000;
      1546: inst = 32'h10408000;
      1547: inst = 32'hc4041bb;
      1548: inst = 32'h8220000;
      1549: inst = 32'h10408000;
      1550: inst = 32'hc4041bc;
      1551: inst = 32'h8220000;
      1552: inst = 32'h10408000;
      1553: inst = 32'hc4041bd;
      1554: inst = 32'h8220000;
      1555: inst = 32'h10408000;
      1556: inst = 32'hc4041be;
      1557: inst = 32'h8220000;
      1558: inst = 32'h10408000;
      1559: inst = 32'hc4041bf;
      1560: inst = 32'h8220000;
      1561: inst = 32'h10408000;
      1562: inst = 32'hc4041c0;
      1563: inst = 32'h8220000;
      1564: inst = 32'h10408000;
      1565: inst = 32'hc4041c1;
      1566: inst = 32'h8220000;
      1567: inst = 32'h10408000;
      1568: inst = 32'hc4041c2;
      1569: inst = 32'h8220000;
      1570: inst = 32'h10408000;
      1571: inst = 32'hc4041c3;
      1572: inst = 32'h8220000;
      1573: inst = 32'h10408000;
      1574: inst = 32'hc4041c4;
      1575: inst = 32'h8220000;
      1576: inst = 32'h10408000;
      1577: inst = 32'hc4041c5;
      1578: inst = 32'h8220000;
      1579: inst = 32'h10408000;
      1580: inst = 32'hc4041c6;
      1581: inst = 32'h8220000;
      1582: inst = 32'h10408000;
      1583: inst = 32'hc4041c7;
      1584: inst = 32'h8220000;
      1585: inst = 32'h10408000;
      1586: inst = 32'hc4041c8;
      1587: inst = 32'h8220000;
      1588: inst = 32'h10408000;
      1589: inst = 32'hc4041c9;
      1590: inst = 32'h8220000;
      1591: inst = 32'h10408000;
      1592: inst = 32'hc4041ca;
      1593: inst = 32'h8220000;
      1594: inst = 32'h10408000;
      1595: inst = 32'hc4041cc;
      1596: inst = 32'h8220000;
      1597: inst = 32'h10408000;
      1598: inst = 32'hc4041cd;
      1599: inst = 32'h8220000;
      1600: inst = 32'h10408000;
      1601: inst = 32'hc4041ce;
      1602: inst = 32'h8220000;
      1603: inst = 32'h10408000;
      1604: inst = 32'hc4041cf;
      1605: inst = 32'h8220000;
      1606: inst = 32'h10408000;
      1607: inst = 32'hc4041d0;
      1608: inst = 32'h8220000;
      1609: inst = 32'h10408000;
      1610: inst = 32'hc4041d1;
      1611: inst = 32'h8220000;
      1612: inst = 32'h10408000;
      1613: inst = 32'hc4041d2;
      1614: inst = 32'h8220000;
      1615: inst = 32'h10408000;
      1616: inst = 32'hc4041d3;
      1617: inst = 32'h8220000;
      1618: inst = 32'h10408000;
      1619: inst = 32'hc4041d4;
      1620: inst = 32'h8220000;
      1621: inst = 32'h10408000;
      1622: inst = 32'hc4041d5;
      1623: inst = 32'h8220000;
      1624: inst = 32'h10408000;
      1625: inst = 32'hc4041d6;
      1626: inst = 32'h8220000;
      1627: inst = 32'h10408000;
      1628: inst = 32'hc4041d7;
      1629: inst = 32'h8220000;
      1630: inst = 32'h10408000;
      1631: inst = 32'hc4041d8;
      1632: inst = 32'h8220000;
      1633: inst = 32'h10408000;
      1634: inst = 32'hc4041d9;
      1635: inst = 32'h8220000;
      1636: inst = 32'h10408000;
      1637: inst = 32'hc404206;
      1638: inst = 32'h8220000;
      1639: inst = 32'h10408000;
      1640: inst = 32'hc404207;
      1641: inst = 32'h8220000;
      1642: inst = 32'h10408000;
      1643: inst = 32'hc404208;
      1644: inst = 32'h8220000;
      1645: inst = 32'h10408000;
      1646: inst = 32'hc404209;
      1647: inst = 32'h8220000;
      1648: inst = 32'h10408000;
      1649: inst = 32'hc40420a;
      1650: inst = 32'h8220000;
      1651: inst = 32'h10408000;
      1652: inst = 32'hc40420b;
      1653: inst = 32'h8220000;
      1654: inst = 32'h10408000;
      1655: inst = 32'hc40420c;
      1656: inst = 32'h8220000;
      1657: inst = 32'h10408000;
      1658: inst = 32'hc40420d;
      1659: inst = 32'h8220000;
      1660: inst = 32'h10408000;
      1661: inst = 32'hc40420e;
      1662: inst = 32'h8220000;
      1663: inst = 32'h10408000;
      1664: inst = 32'hc40420f;
      1665: inst = 32'h8220000;
      1666: inst = 32'h10408000;
      1667: inst = 32'hc404210;
      1668: inst = 32'h8220000;
      1669: inst = 32'h10408000;
      1670: inst = 32'hc404211;
      1671: inst = 32'h8220000;
      1672: inst = 32'h10408000;
      1673: inst = 32'hc404212;
      1674: inst = 32'h8220000;
      1675: inst = 32'h10408000;
      1676: inst = 32'hc404213;
      1677: inst = 32'h8220000;
      1678: inst = 32'h10408000;
      1679: inst = 32'hc404214;
      1680: inst = 32'h8220000;
      1681: inst = 32'h10408000;
      1682: inst = 32'hc404215;
      1683: inst = 32'h8220000;
      1684: inst = 32'h10408000;
      1685: inst = 32'hc404216;
      1686: inst = 32'h8220000;
      1687: inst = 32'h10408000;
      1688: inst = 32'hc404217;
      1689: inst = 32'h8220000;
      1690: inst = 32'h10408000;
      1691: inst = 32'hc404218;
      1692: inst = 32'h8220000;
      1693: inst = 32'h10408000;
      1694: inst = 32'hc404219;
      1695: inst = 32'h8220000;
      1696: inst = 32'h10408000;
      1697: inst = 32'hc40421a;
      1698: inst = 32'h8220000;
      1699: inst = 32'h10408000;
      1700: inst = 32'hc40421b;
      1701: inst = 32'h8220000;
      1702: inst = 32'h10408000;
      1703: inst = 32'hc40421c;
      1704: inst = 32'h8220000;
      1705: inst = 32'h10408000;
      1706: inst = 32'hc40421d;
      1707: inst = 32'h8220000;
      1708: inst = 32'h10408000;
      1709: inst = 32'hc40421e;
      1710: inst = 32'h8220000;
      1711: inst = 32'h10408000;
      1712: inst = 32'hc40421f;
      1713: inst = 32'h8220000;
      1714: inst = 32'h10408000;
      1715: inst = 32'hc404220;
      1716: inst = 32'h8220000;
      1717: inst = 32'h10408000;
      1718: inst = 32'hc404221;
      1719: inst = 32'h8220000;
      1720: inst = 32'h10408000;
      1721: inst = 32'hc404222;
      1722: inst = 32'h8220000;
      1723: inst = 32'h10408000;
      1724: inst = 32'hc404223;
      1725: inst = 32'h8220000;
      1726: inst = 32'h10408000;
      1727: inst = 32'hc404224;
      1728: inst = 32'h8220000;
      1729: inst = 32'h10408000;
      1730: inst = 32'hc404225;
      1731: inst = 32'h8220000;
      1732: inst = 32'h10408000;
      1733: inst = 32'hc404226;
      1734: inst = 32'h8220000;
      1735: inst = 32'h10408000;
      1736: inst = 32'hc404227;
      1737: inst = 32'h8220000;
      1738: inst = 32'h10408000;
      1739: inst = 32'hc404228;
      1740: inst = 32'h8220000;
      1741: inst = 32'h10408000;
      1742: inst = 32'hc404229;
      1743: inst = 32'h8220000;
      1744: inst = 32'h10408000;
      1745: inst = 32'hc40422a;
      1746: inst = 32'h8220000;
      1747: inst = 32'h10408000;
      1748: inst = 32'hc40422c;
      1749: inst = 32'h8220000;
      1750: inst = 32'h10408000;
      1751: inst = 32'hc40422d;
      1752: inst = 32'h8220000;
      1753: inst = 32'h10408000;
      1754: inst = 32'hc40422e;
      1755: inst = 32'h8220000;
      1756: inst = 32'h10408000;
      1757: inst = 32'hc40422f;
      1758: inst = 32'h8220000;
      1759: inst = 32'h10408000;
      1760: inst = 32'hc404230;
      1761: inst = 32'h8220000;
      1762: inst = 32'h10408000;
      1763: inst = 32'hc404231;
      1764: inst = 32'h8220000;
      1765: inst = 32'h10408000;
      1766: inst = 32'hc404232;
      1767: inst = 32'h8220000;
      1768: inst = 32'h10408000;
      1769: inst = 32'hc404233;
      1770: inst = 32'h8220000;
      1771: inst = 32'h10408000;
      1772: inst = 32'hc404234;
      1773: inst = 32'h8220000;
      1774: inst = 32'h10408000;
      1775: inst = 32'hc404235;
      1776: inst = 32'h8220000;
      1777: inst = 32'h10408000;
      1778: inst = 32'hc404236;
      1779: inst = 32'h8220000;
      1780: inst = 32'h10408000;
      1781: inst = 32'hc404237;
      1782: inst = 32'h8220000;
      1783: inst = 32'h10408000;
      1784: inst = 32'hc404238;
      1785: inst = 32'h8220000;
      1786: inst = 32'h10408000;
      1787: inst = 32'hc404239;
      1788: inst = 32'h8220000;
      1789: inst = 32'h10408000;
      1790: inst = 32'hc40423a;
      1791: inst = 32'h8220000;
      1792: inst = 32'h10408000;
      1793: inst = 32'hc40423b;
      1794: inst = 32'h8220000;
      1795: inst = 32'h10408000;
      1796: inst = 32'hc404264;
      1797: inst = 32'h8220000;
      1798: inst = 32'h10408000;
      1799: inst = 32'hc404265;
      1800: inst = 32'h8220000;
      1801: inst = 32'h10408000;
      1802: inst = 32'hc404266;
      1803: inst = 32'h8220000;
      1804: inst = 32'h10408000;
      1805: inst = 32'hc404267;
      1806: inst = 32'h8220000;
      1807: inst = 32'h10408000;
      1808: inst = 32'hc404268;
      1809: inst = 32'h8220000;
      1810: inst = 32'h10408000;
      1811: inst = 32'hc404269;
      1812: inst = 32'h8220000;
      1813: inst = 32'h10408000;
      1814: inst = 32'hc40426a;
      1815: inst = 32'h8220000;
      1816: inst = 32'h10408000;
      1817: inst = 32'hc40426b;
      1818: inst = 32'h8220000;
      1819: inst = 32'h10408000;
      1820: inst = 32'hc40426c;
      1821: inst = 32'h8220000;
      1822: inst = 32'h10408000;
      1823: inst = 32'hc40426d;
      1824: inst = 32'h8220000;
      1825: inst = 32'h10408000;
      1826: inst = 32'hc40426e;
      1827: inst = 32'h8220000;
      1828: inst = 32'h10408000;
      1829: inst = 32'hc40426f;
      1830: inst = 32'h8220000;
      1831: inst = 32'h10408000;
      1832: inst = 32'hc404270;
      1833: inst = 32'h8220000;
      1834: inst = 32'h10408000;
      1835: inst = 32'hc404271;
      1836: inst = 32'h8220000;
      1837: inst = 32'h10408000;
      1838: inst = 32'hc404272;
      1839: inst = 32'h8220000;
      1840: inst = 32'h10408000;
      1841: inst = 32'hc404273;
      1842: inst = 32'h8220000;
      1843: inst = 32'h10408000;
      1844: inst = 32'hc404274;
      1845: inst = 32'h8220000;
      1846: inst = 32'h10408000;
      1847: inst = 32'hc404275;
      1848: inst = 32'h8220000;
      1849: inst = 32'h10408000;
      1850: inst = 32'hc404276;
      1851: inst = 32'h8220000;
      1852: inst = 32'h10408000;
      1853: inst = 32'hc404277;
      1854: inst = 32'h8220000;
      1855: inst = 32'h10408000;
      1856: inst = 32'hc404278;
      1857: inst = 32'h8220000;
      1858: inst = 32'h10408000;
      1859: inst = 32'hc404279;
      1860: inst = 32'h8220000;
      1861: inst = 32'h10408000;
      1862: inst = 32'hc40427a;
      1863: inst = 32'h8220000;
      1864: inst = 32'h10408000;
      1865: inst = 32'hc40427b;
      1866: inst = 32'h8220000;
      1867: inst = 32'h10408000;
      1868: inst = 32'hc40427c;
      1869: inst = 32'h8220000;
      1870: inst = 32'h10408000;
      1871: inst = 32'hc40427d;
      1872: inst = 32'h8220000;
      1873: inst = 32'h10408000;
      1874: inst = 32'hc40427e;
      1875: inst = 32'h8220000;
      1876: inst = 32'h10408000;
      1877: inst = 32'hc40427f;
      1878: inst = 32'h8220000;
      1879: inst = 32'h10408000;
      1880: inst = 32'hc404280;
      1881: inst = 32'h8220000;
      1882: inst = 32'h10408000;
      1883: inst = 32'hc404281;
      1884: inst = 32'h8220000;
      1885: inst = 32'h10408000;
      1886: inst = 32'hc404282;
      1887: inst = 32'h8220000;
      1888: inst = 32'h10408000;
      1889: inst = 32'hc404283;
      1890: inst = 32'h8220000;
      1891: inst = 32'h10408000;
      1892: inst = 32'hc404284;
      1893: inst = 32'h8220000;
      1894: inst = 32'h10408000;
      1895: inst = 32'hc404285;
      1896: inst = 32'h8220000;
      1897: inst = 32'h10408000;
      1898: inst = 32'hc404286;
      1899: inst = 32'h8220000;
      1900: inst = 32'h10408000;
      1901: inst = 32'hc404287;
      1902: inst = 32'h8220000;
      1903: inst = 32'h10408000;
      1904: inst = 32'hc404288;
      1905: inst = 32'h8220000;
      1906: inst = 32'h10408000;
      1907: inst = 32'hc404289;
      1908: inst = 32'h8220000;
      1909: inst = 32'h10408000;
      1910: inst = 32'hc40428a;
      1911: inst = 32'h8220000;
      1912: inst = 32'h10408000;
      1913: inst = 32'hc40428c;
      1914: inst = 32'h8220000;
      1915: inst = 32'h10408000;
      1916: inst = 32'hc40428d;
      1917: inst = 32'h8220000;
      1918: inst = 32'h10408000;
      1919: inst = 32'hc40428e;
      1920: inst = 32'h8220000;
      1921: inst = 32'h10408000;
      1922: inst = 32'hc40428f;
      1923: inst = 32'h8220000;
      1924: inst = 32'h10408000;
      1925: inst = 32'hc404290;
      1926: inst = 32'h8220000;
      1927: inst = 32'h10408000;
      1928: inst = 32'hc404291;
      1929: inst = 32'h8220000;
      1930: inst = 32'h10408000;
      1931: inst = 32'hc404292;
      1932: inst = 32'h8220000;
      1933: inst = 32'h10408000;
      1934: inst = 32'hc404293;
      1935: inst = 32'h8220000;
      1936: inst = 32'h10408000;
      1937: inst = 32'hc404294;
      1938: inst = 32'h8220000;
      1939: inst = 32'h10408000;
      1940: inst = 32'hc404295;
      1941: inst = 32'h8220000;
      1942: inst = 32'h10408000;
      1943: inst = 32'hc404296;
      1944: inst = 32'h8220000;
      1945: inst = 32'h10408000;
      1946: inst = 32'hc404297;
      1947: inst = 32'h8220000;
      1948: inst = 32'h10408000;
      1949: inst = 32'hc404298;
      1950: inst = 32'h8220000;
      1951: inst = 32'h10408000;
      1952: inst = 32'hc404299;
      1953: inst = 32'h8220000;
      1954: inst = 32'h10408000;
      1955: inst = 32'hc40429a;
      1956: inst = 32'h8220000;
      1957: inst = 32'h10408000;
      1958: inst = 32'hc40429b;
      1959: inst = 32'h8220000;
      1960: inst = 32'h10408000;
      1961: inst = 32'hc4042c4;
      1962: inst = 32'h8220000;
      1963: inst = 32'h10408000;
      1964: inst = 32'hc4042c5;
      1965: inst = 32'h8220000;
      1966: inst = 32'h10408000;
      1967: inst = 32'hc4042c6;
      1968: inst = 32'h8220000;
      1969: inst = 32'h10408000;
      1970: inst = 32'hc4042c7;
      1971: inst = 32'h8220000;
      1972: inst = 32'h10408000;
      1973: inst = 32'hc4042c8;
      1974: inst = 32'h8220000;
      1975: inst = 32'h10408000;
      1976: inst = 32'hc4042c9;
      1977: inst = 32'h8220000;
      1978: inst = 32'h10408000;
      1979: inst = 32'hc4042ca;
      1980: inst = 32'h8220000;
      1981: inst = 32'h10408000;
      1982: inst = 32'hc4042cb;
      1983: inst = 32'h8220000;
      1984: inst = 32'h10408000;
      1985: inst = 32'hc4042cc;
      1986: inst = 32'h8220000;
      1987: inst = 32'h10408000;
      1988: inst = 32'hc4042cd;
      1989: inst = 32'h8220000;
      1990: inst = 32'h10408000;
      1991: inst = 32'hc4042ce;
      1992: inst = 32'h8220000;
      1993: inst = 32'h10408000;
      1994: inst = 32'hc4042cf;
      1995: inst = 32'h8220000;
      1996: inst = 32'h10408000;
      1997: inst = 32'hc4042d0;
      1998: inst = 32'h8220000;
      1999: inst = 32'h10408000;
      2000: inst = 32'hc4042d1;
      2001: inst = 32'h8220000;
      2002: inst = 32'h10408000;
      2003: inst = 32'hc4042d2;
      2004: inst = 32'h8220000;
      2005: inst = 32'h10408000;
      2006: inst = 32'hc4042d3;
      2007: inst = 32'h8220000;
      2008: inst = 32'h10408000;
      2009: inst = 32'hc4042d4;
      2010: inst = 32'h8220000;
      2011: inst = 32'h10408000;
      2012: inst = 32'hc4042d5;
      2013: inst = 32'h8220000;
      2014: inst = 32'h10408000;
      2015: inst = 32'hc4042d6;
      2016: inst = 32'h8220000;
      2017: inst = 32'h10408000;
      2018: inst = 32'hc4042d7;
      2019: inst = 32'h8220000;
      2020: inst = 32'h10408000;
      2021: inst = 32'hc4042d8;
      2022: inst = 32'h8220000;
      2023: inst = 32'h10408000;
      2024: inst = 32'hc4042d9;
      2025: inst = 32'h8220000;
      2026: inst = 32'h10408000;
      2027: inst = 32'hc4042da;
      2028: inst = 32'h8220000;
      2029: inst = 32'h10408000;
      2030: inst = 32'hc4042db;
      2031: inst = 32'h8220000;
      2032: inst = 32'h10408000;
      2033: inst = 32'hc4042dc;
      2034: inst = 32'h8220000;
      2035: inst = 32'h10408000;
      2036: inst = 32'hc4042dd;
      2037: inst = 32'h8220000;
      2038: inst = 32'h10408000;
      2039: inst = 32'hc4042de;
      2040: inst = 32'h8220000;
      2041: inst = 32'h10408000;
      2042: inst = 32'hc4042df;
      2043: inst = 32'h8220000;
      2044: inst = 32'h10408000;
      2045: inst = 32'hc4042e0;
      2046: inst = 32'h8220000;
      2047: inst = 32'h10408000;
      2048: inst = 32'hc4042e1;
      2049: inst = 32'h8220000;
      2050: inst = 32'h10408000;
      2051: inst = 32'hc4042e2;
      2052: inst = 32'h8220000;
      2053: inst = 32'h10408000;
      2054: inst = 32'hc4042e3;
      2055: inst = 32'h8220000;
      2056: inst = 32'h10408000;
      2057: inst = 32'hc4042e4;
      2058: inst = 32'h8220000;
      2059: inst = 32'h10408000;
      2060: inst = 32'hc4042e5;
      2061: inst = 32'h8220000;
      2062: inst = 32'h10408000;
      2063: inst = 32'hc4042e6;
      2064: inst = 32'h8220000;
      2065: inst = 32'h10408000;
      2066: inst = 32'hc4042e7;
      2067: inst = 32'h8220000;
      2068: inst = 32'h10408000;
      2069: inst = 32'hc4042e8;
      2070: inst = 32'h8220000;
      2071: inst = 32'h10408000;
      2072: inst = 32'hc4042e9;
      2073: inst = 32'h8220000;
      2074: inst = 32'h10408000;
      2075: inst = 32'hc4042ee;
      2076: inst = 32'h8220000;
      2077: inst = 32'h10408000;
      2078: inst = 32'hc4042ef;
      2079: inst = 32'h8220000;
      2080: inst = 32'h10408000;
      2081: inst = 32'hc4042f0;
      2082: inst = 32'h8220000;
      2083: inst = 32'h10408000;
      2084: inst = 32'hc4042f1;
      2085: inst = 32'h8220000;
      2086: inst = 32'h10408000;
      2087: inst = 32'hc4042f2;
      2088: inst = 32'h8220000;
      2089: inst = 32'h10408000;
      2090: inst = 32'hc4042f3;
      2091: inst = 32'h8220000;
      2092: inst = 32'h10408000;
      2093: inst = 32'hc4042f4;
      2094: inst = 32'h8220000;
      2095: inst = 32'h10408000;
      2096: inst = 32'hc4042f5;
      2097: inst = 32'h8220000;
      2098: inst = 32'h10408000;
      2099: inst = 32'hc4042f6;
      2100: inst = 32'h8220000;
      2101: inst = 32'h10408000;
      2102: inst = 32'hc4042f7;
      2103: inst = 32'h8220000;
      2104: inst = 32'h10408000;
      2105: inst = 32'hc4042f8;
      2106: inst = 32'h8220000;
      2107: inst = 32'h10408000;
      2108: inst = 32'hc4042f9;
      2109: inst = 32'h8220000;
      2110: inst = 32'h10408000;
      2111: inst = 32'hc4042fa;
      2112: inst = 32'h8220000;
      2113: inst = 32'h10408000;
      2114: inst = 32'hc4042fb;
      2115: inst = 32'h8220000;
      2116: inst = 32'h10408000;
      2117: inst = 32'hc404324;
      2118: inst = 32'h8220000;
      2119: inst = 32'h10408000;
      2120: inst = 32'hc404325;
      2121: inst = 32'h8220000;
      2122: inst = 32'h10408000;
      2123: inst = 32'hc404326;
      2124: inst = 32'h8220000;
      2125: inst = 32'h10408000;
      2126: inst = 32'hc404327;
      2127: inst = 32'h8220000;
      2128: inst = 32'h10408000;
      2129: inst = 32'hc404328;
      2130: inst = 32'h8220000;
      2131: inst = 32'h10408000;
      2132: inst = 32'hc404329;
      2133: inst = 32'h8220000;
      2134: inst = 32'h10408000;
      2135: inst = 32'hc40432a;
      2136: inst = 32'h8220000;
      2137: inst = 32'h10408000;
      2138: inst = 32'hc40432b;
      2139: inst = 32'h8220000;
      2140: inst = 32'h10408000;
      2141: inst = 32'hc40432c;
      2142: inst = 32'h8220000;
      2143: inst = 32'h10408000;
      2144: inst = 32'hc40432d;
      2145: inst = 32'h8220000;
      2146: inst = 32'h10408000;
      2147: inst = 32'hc40432e;
      2148: inst = 32'h8220000;
      2149: inst = 32'h10408000;
      2150: inst = 32'hc40432f;
      2151: inst = 32'h8220000;
      2152: inst = 32'h10408000;
      2153: inst = 32'hc404330;
      2154: inst = 32'h8220000;
      2155: inst = 32'h10408000;
      2156: inst = 32'hc404331;
      2157: inst = 32'h8220000;
      2158: inst = 32'h10408000;
      2159: inst = 32'hc404332;
      2160: inst = 32'h8220000;
      2161: inst = 32'h10408000;
      2162: inst = 32'hc404333;
      2163: inst = 32'h8220000;
      2164: inst = 32'h10408000;
      2165: inst = 32'hc404334;
      2166: inst = 32'h8220000;
      2167: inst = 32'h10408000;
      2168: inst = 32'hc404335;
      2169: inst = 32'h8220000;
      2170: inst = 32'h10408000;
      2171: inst = 32'hc404336;
      2172: inst = 32'h8220000;
      2173: inst = 32'h10408000;
      2174: inst = 32'hc404337;
      2175: inst = 32'h8220000;
      2176: inst = 32'h10408000;
      2177: inst = 32'hc404338;
      2178: inst = 32'h8220000;
      2179: inst = 32'h10408000;
      2180: inst = 32'hc404339;
      2181: inst = 32'h8220000;
      2182: inst = 32'h10408000;
      2183: inst = 32'hc40433a;
      2184: inst = 32'h8220000;
      2185: inst = 32'h10408000;
      2186: inst = 32'hc40433b;
      2187: inst = 32'h8220000;
      2188: inst = 32'h10408000;
      2189: inst = 32'hc40433c;
      2190: inst = 32'h8220000;
      2191: inst = 32'h10408000;
      2192: inst = 32'hc40433d;
      2193: inst = 32'h8220000;
      2194: inst = 32'h10408000;
      2195: inst = 32'hc40433e;
      2196: inst = 32'h8220000;
      2197: inst = 32'h10408000;
      2198: inst = 32'hc40433f;
      2199: inst = 32'h8220000;
      2200: inst = 32'h10408000;
      2201: inst = 32'hc404340;
      2202: inst = 32'h8220000;
      2203: inst = 32'h10408000;
      2204: inst = 32'hc404341;
      2205: inst = 32'h8220000;
      2206: inst = 32'h10408000;
      2207: inst = 32'hc404342;
      2208: inst = 32'h8220000;
      2209: inst = 32'h10408000;
      2210: inst = 32'hc404343;
      2211: inst = 32'h8220000;
      2212: inst = 32'h10408000;
      2213: inst = 32'hc404344;
      2214: inst = 32'h8220000;
      2215: inst = 32'h10408000;
      2216: inst = 32'hc404345;
      2217: inst = 32'h8220000;
      2218: inst = 32'h10408000;
      2219: inst = 32'hc404346;
      2220: inst = 32'h8220000;
      2221: inst = 32'h10408000;
      2222: inst = 32'hc404347;
      2223: inst = 32'h8220000;
      2224: inst = 32'h10408000;
      2225: inst = 32'hc404348;
      2226: inst = 32'h8220000;
      2227: inst = 32'h10408000;
      2228: inst = 32'hc40434f;
      2229: inst = 32'h8220000;
      2230: inst = 32'h10408000;
      2231: inst = 32'hc404350;
      2232: inst = 32'h8220000;
      2233: inst = 32'h10408000;
      2234: inst = 32'hc404351;
      2235: inst = 32'h8220000;
      2236: inst = 32'h10408000;
      2237: inst = 32'hc404352;
      2238: inst = 32'h8220000;
      2239: inst = 32'h10408000;
      2240: inst = 32'hc404353;
      2241: inst = 32'h8220000;
      2242: inst = 32'h10408000;
      2243: inst = 32'hc404354;
      2244: inst = 32'h8220000;
      2245: inst = 32'h10408000;
      2246: inst = 32'hc404355;
      2247: inst = 32'h8220000;
      2248: inst = 32'h10408000;
      2249: inst = 32'hc404356;
      2250: inst = 32'h8220000;
      2251: inst = 32'h10408000;
      2252: inst = 32'hc404357;
      2253: inst = 32'h8220000;
      2254: inst = 32'h10408000;
      2255: inst = 32'hc404358;
      2256: inst = 32'h8220000;
      2257: inst = 32'h10408000;
      2258: inst = 32'hc404359;
      2259: inst = 32'h8220000;
      2260: inst = 32'h10408000;
      2261: inst = 32'hc40435a;
      2262: inst = 32'h8220000;
      2263: inst = 32'h10408000;
      2264: inst = 32'hc40435b;
      2265: inst = 32'h8220000;
      2266: inst = 32'h10408000;
      2267: inst = 32'hc404384;
      2268: inst = 32'h8220000;
      2269: inst = 32'h10408000;
      2270: inst = 32'hc404385;
      2271: inst = 32'h8220000;
      2272: inst = 32'h10408000;
      2273: inst = 32'hc404386;
      2274: inst = 32'h8220000;
      2275: inst = 32'h10408000;
      2276: inst = 32'hc404387;
      2277: inst = 32'h8220000;
      2278: inst = 32'h10408000;
      2279: inst = 32'hc404388;
      2280: inst = 32'h8220000;
      2281: inst = 32'h10408000;
      2282: inst = 32'hc404389;
      2283: inst = 32'h8220000;
      2284: inst = 32'h10408000;
      2285: inst = 32'hc40438a;
      2286: inst = 32'h8220000;
      2287: inst = 32'h10408000;
      2288: inst = 32'hc40438b;
      2289: inst = 32'h8220000;
      2290: inst = 32'h10408000;
      2291: inst = 32'hc40438c;
      2292: inst = 32'h8220000;
      2293: inst = 32'h10408000;
      2294: inst = 32'hc40438d;
      2295: inst = 32'h8220000;
      2296: inst = 32'h10408000;
      2297: inst = 32'hc40438e;
      2298: inst = 32'h8220000;
      2299: inst = 32'h10408000;
      2300: inst = 32'hc40438f;
      2301: inst = 32'h8220000;
      2302: inst = 32'h10408000;
      2303: inst = 32'hc404390;
      2304: inst = 32'h8220000;
      2305: inst = 32'h10408000;
      2306: inst = 32'hc404391;
      2307: inst = 32'h8220000;
      2308: inst = 32'h10408000;
      2309: inst = 32'hc404392;
      2310: inst = 32'h8220000;
      2311: inst = 32'h10408000;
      2312: inst = 32'hc404393;
      2313: inst = 32'h8220000;
      2314: inst = 32'h10408000;
      2315: inst = 32'hc404394;
      2316: inst = 32'h8220000;
      2317: inst = 32'h10408000;
      2318: inst = 32'hc404395;
      2319: inst = 32'h8220000;
      2320: inst = 32'h10408000;
      2321: inst = 32'hc404396;
      2322: inst = 32'h8220000;
      2323: inst = 32'h10408000;
      2324: inst = 32'hc404397;
      2325: inst = 32'h8220000;
      2326: inst = 32'h10408000;
      2327: inst = 32'hc404398;
      2328: inst = 32'h8220000;
      2329: inst = 32'h10408000;
      2330: inst = 32'hc404399;
      2331: inst = 32'h8220000;
      2332: inst = 32'h10408000;
      2333: inst = 32'hc40439a;
      2334: inst = 32'h8220000;
      2335: inst = 32'h10408000;
      2336: inst = 32'hc40439b;
      2337: inst = 32'h8220000;
      2338: inst = 32'h10408000;
      2339: inst = 32'hc40439c;
      2340: inst = 32'h8220000;
      2341: inst = 32'h10408000;
      2342: inst = 32'hc40439d;
      2343: inst = 32'h8220000;
      2344: inst = 32'h10408000;
      2345: inst = 32'hc40439e;
      2346: inst = 32'h8220000;
      2347: inst = 32'h10408000;
      2348: inst = 32'hc40439f;
      2349: inst = 32'h8220000;
      2350: inst = 32'h10408000;
      2351: inst = 32'hc4043a0;
      2352: inst = 32'h8220000;
      2353: inst = 32'h10408000;
      2354: inst = 32'hc4043a1;
      2355: inst = 32'h8220000;
      2356: inst = 32'h10408000;
      2357: inst = 32'hc4043a2;
      2358: inst = 32'h8220000;
      2359: inst = 32'h10408000;
      2360: inst = 32'hc4043a3;
      2361: inst = 32'h8220000;
      2362: inst = 32'h10408000;
      2363: inst = 32'hc4043a4;
      2364: inst = 32'h8220000;
      2365: inst = 32'h10408000;
      2366: inst = 32'hc4043a5;
      2367: inst = 32'h8220000;
      2368: inst = 32'h10408000;
      2369: inst = 32'hc4043a6;
      2370: inst = 32'h8220000;
      2371: inst = 32'h10408000;
      2372: inst = 32'hc4043b1;
      2373: inst = 32'h8220000;
      2374: inst = 32'h10408000;
      2375: inst = 32'hc4043b2;
      2376: inst = 32'h8220000;
      2377: inst = 32'h10408000;
      2378: inst = 32'hc4043b3;
      2379: inst = 32'h8220000;
      2380: inst = 32'h10408000;
      2381: inst = 32'hc4043b4;
      2382: inst = 32'h8220000;
      2383: inst = 32'h10408000;
      2384: inst = 32'hc4043b5;
      2385: inst = 32'h8220000;
      2386: inst = 32'h10408000;
      2387: inst = 32'hc4043b6;
      2388: inst = 32'h8220000;
      2389: inst = 32'h10408000;
      2390: inst = 32'hc4043b7;
      2391: inst = 32'h8220000;
      2392: inst = 32'h10408000;
      2393: inst = 32'hc4043b8;
      2394: inst = 32'h8220000;
      2395: inst = 32'h10408000;
      2396: inst = 32'hc4043b9;
      2397: inst = 32'h8220000;
      2398: inst = 32'h10408000;
      2399: inst = 32'hc4043ba;
      2400: inst = 32'h8220000;
      2401: inst = 32'h10408000;
      2402: inst = 32'hc4043bb;
      2403: inst = 32'h8220000;
      2404: inst = 32'h10408000;
      2405: inst = 32'hc4043e4;
      2406: inst = 32'h8220000;
      2407: inst = 32'h10408000;
      2408: inst = 32'hc4043e5;
      2409: inst = 32'h8220000;
      2410: inst = 32'h10408000;
      2411: inst = 32'hc4043e6;
      2412: inst = 32'h8220000;
      2413: inst = 32'h10408000;
      2414: inst = 32'hc4043e7;
      2415: inst = 32'h8220000;
      2416: inst = 32'h10408000;
      2417: inst = 32'hc4043e8;
      2418: inst = 32'h8220000;
      2419: inst = 32'h10408000;
      2420: inst = 32'hc4043e9;
      2421: inst = 32'h8220000;
      2422: inst = 32'h10408000;
      2423: inst = 32'hc4043ea;
      2424: inst = 32'h8220000;
      2425: inst = 32'h10408000;
      2426: inst = 32'hc4043eb;
      2427: inst = 32'h8220000;
      2428: inst = 32'h10408000;
      2429: inst = 32'hc4043ec;
      2430: inst = 32'h8220000;
      2431: inst = 32'h10408000;
      2432: inst = 32'hc4043ed;
      2433: inst = 32'h8220000;
      2434: inst = 32'h10408000;
      2435: inst = 32'hc4043ee;
      2436: inst = 32'h8220000;
      2437: inst = 32'h10408000;
      2438: inst = 32'hc4043ef;
      2439: inst = 32'h8220000;
      2440: inst = 32'h10408000;
      2441: inst = 32'hc4043f0;
      2442: inst = 32'h8220000;
      2443: inst = 32'h10408000;
      2444: inst = 32'hc4043f1;
      2445: inst = 32'h8220000;
      2446: inst = 32'h10408000;
      2447: inst = 32'hc4043f2;
      2448: inst = 32'h8220000;
      2449: inst = 32'h10408000;
      2450: inst = 32'hc4043f3;
      2451: inst = 32'h8220000;
      2452: inst = 32'h10408000;
      2453: inst = 32'hc4043f4;
      2454: inst = 32'h8220000;
      2455: inst = 32'h10408000;
      2456: inst = 32'hc4043f5;
      2457: inst = 32'h8220000;
      2458: inst = 32'h10408000;
      2459: inst = 32'hc4043f6;
      2460: inst = 32'h8220000;
      2461: inst = 32'h10408000;
      2462: inst = 32'hc4043f7;
      2463: inst = 32'h8220000;
      2464: inst = 32'h10408000;
      2465: inst = 32'hc4043f8;
      2466: inst = 32'h8220000;
      2467: inst = 32'h10408000;
      2468: inst = 32'hc4043f9;
      2469: inst = 32'h8220000;
      2470: inst = 32'h10408000;
      2471: inst = 32'hc4043fa;
      2472: inst = 32'h8220000;
      2473: inst = 32'h10408000;
      2474: inst = 32'hc4043fb;
      2475: inst = 32'h8220000;
      2476: inst = 32'h10408000;
      2477: inst = 32'hc4043fc;
      2478: inst = 32'h8220000;
      2479: inst = 32'h10408000;
      2480: inst = 32'hc4043fd;
      2481: inst = 32'h8220000;
      2482: inst = 32'h10408000;
      2483: inst = 32'hc4043fe;
      2484: inst = 32'h8220000;
      2485: inst = 32'h10408000;
      2486: inst = 32'hc4043ff;
      2487: inst = 32'h8220000;
      2488: inst = 32'h10408000;
      2489: inst = 32'hc404400;
      2490: inst = 32'h8220000;
      2491: inst = 32'h10408000;
      2492: inst = 32'hc404401;
      2493: inst = 32'h8220000;
      2494: inst = 32'h10408000;
      2495: inst = 32'hc404402;
      2496: inst = 32'h8220000;
      2497: inst = 32'h10408000;
      2498: inst = 32'hc404403;
      2499: inst = 32'h8220000;
      2500: inst = 32'h10408000;
      2501: inst = 32'hc404404;
      2502: inst = 32'h8220000;
      2503: inst = 32'h10408000;
      2504: inst = 32'hc404405;
      2505: inst = 32'h8220000;
      2506: inst = 32'h10408000;
      2507: inst = 32'hc404412;
      2508: inst = 32'h8220000;
      2509: inst = 32'h10408000;
      2510: inst = 32'hc404413;
      2511: inst = 32'h8220000;
      2512: inst = 32'h10408000;
      2513: inst = 32'hc404414;
      2514: inst = 32'h8220000;
      2515: inst = 32'h10408000;
      2516: inst = 32'hc404415;
      2517: inst = 32'h8220000;
      2518: inst = 32'h10408000;
      2519: inst = 32'hc404416;
      2520: inst = 32'h8220000;
      2521: inst = 32'h10408000;
      2522: inst = 32'hc404417;
      2523: inst = 32'h8220000;
      2524: inst = 32'h10408000;
      2525: inst = 32'hc404418;
      2526: inst = 32'h8220000;
      2527: inst = 32'h10408000;
      2528: inst = 32'hc404419;
      2529: inst = 32'h8220000;
      2530: inst = 32'h10408000;
      2531: inst = 32'hc40441a;
      2532: inst = 32'h8220000;
      2533: inst = 32'h10408000;
      2534: inst = 32'hc40441b;
      2535: inst = 32'h8220000;
      2536: inst = 32'h10408000;
      2537: inst = 32'hc404444;
      2538: inst = 32'h8220000;
      2539: inst = 32'h10408000;
      2540: inst = 32'hc404445;
      2541: inst = 32'h8220000;
      2542: inst = 32'h10408000;
      2543: inst = 32'hc404446;
      2544: inst = 32'h8220000;
      2545: inst = 32'h10408000;
      2546: inst = 32'hc404447;
      2547: inst = 32'h8220000;
      2548: inst = 32'h10408000;
      2549: inst = 32'hc404448;
      2550: inst = 32'h8220000;
      2551: inst = 32'h10408000;
      2552: inst = 32'hc404449;
      2553: inst = 32'h8220000;
      2554: inst = 32'h10408000;
      2555: inst = 32'hc40444a;
      2556: inst = 32'h8220000;
      2557: inst = 32'h10408000;
      2558: inst = 32'hc40444b;
      2559: inst = 32'h8220000;
      2560: inst = 32'h10408000;
      2561: inst = 32'hc40444c;
      2562: inst = 32'h8220000;
      2563: inst = 32'h10408000;
      2564: inst = 32'hc40444d;
      2565: inst = 32'h8220000;
      2566: inst = 32'h10408000;
      2567: inst = 32'hc40444e;
      2568: inst = 32'h8220000;
      2569: inst = 32'h10408000;
      2570: inst = 32'hc40444f;
      2571: inst = 32'h8220000;
      2572: inst = 32'h10408000;
      2573: inst = 32'hc404450;
      2574: inst = 32'h8220000;
      2575: inst = 32'h10408000;
      2576: inst = 32'hc404451;
      2577: inst = 32'h8220000;
      2578: inst = 32'h10408000;
      2579: inst = 32'hc404452;
      2580: inst = 32'h8220000;
      2581: inst = 32'h10408000;
      2582: inst = 32'hc404453;
      2583: inst = 32'h8220000;
      2584: inst = 32'h10408000;
      2585: inst = 32'hc404454;
      2586: inst = 32'h8220000;
      2587: inst = 32'h10408000;
      2588: inst = 32'hc404455;
      2589: inst = 32'h8220000;
      2590: inst = 32'h10408000;
      2591: inst = 32'hc404456;
      2592: inst = 32'h8220000;
      2593: inst = 32'h10408000;
      2594: inst = 32'hc404457;
      2595: inst = 32'h8220000;
      2596: inst = 32'h10408000;
      2597: inst = 32'hc404458;
      2598: inst = 32'h8220000;
      2599: inst = 32'h10408000;
      2600: inst = 32'hc404459;
      2601: inst = 32'h8220000;
      2602: inst = 32'h10408000;
      2603: inst = 32'hc40445a;
      2604: inst = 32'h8220000;
      2605: inst = 32'h10408000;
      2606: inst = 32'hc40445b;
      2607: inst = 32'h8220000;
      2608: inst = 32'h10408000;
      2609: inst = 32'hc40445c;
      2610: inst = 32'h8220000;
      2611: inst = 32'h10408000;
      2612: inst = 32'hc40445d;
      2613: inst = 32'h8220000;
      2614: inst = 32'h10408000;
      2615: inst = 32'hc40445e;
      2616: inst = 32'h8220000;
      2617: inst = 32'h10408000;
      2618: inst = 32'hc40445f;
      2619: inst = 32'h8220000;
      2620: inst = 32'h10408000;
      2621: inst = 32'hc404460;
      2622: inst = 32'h8220000;
      2623: inst = 32'h10408000;
      2624: inst = 32'hc404461;
      2625: inst = 32'h8220000;
      2626: inst = 32'h10408000;
      2627: inst = 32'hc404462;
      2628: inst = 32'h8220000;
      2629: inst = 32'h10408000;
      2630: inst = 32'hc404463;
      2631: inst = 32'h8220000;
      2632: inst = 32'h10408000;
      2633: inst = 32'hc404464;
      2634: inst = 32'h8220000;
      2635: inst = 32'h10408000;
      2636: inst = 32'hc404465;
      2637: inst = 32'h8220000;
      2638: inst = 32'h10408000;
      2639: inst = 32'hc404466;
      2640: inst = 32'h8220000;
      2641: inst = 32'h10408000;
      2642: inst = 32'hc404467;
      2643: inst = 32'h8220000;
      2644: inst = 32'h10408000;
      2645: inst = 32'hc404468;
      2646: inst = 32'h8220000;
      2647: inst = 32'h10408000;
      2648: inst = 32'hc404469;
      2649: inst = 32'h8220000;
      2650: inst = 32'h10408000;
      2651: inst = 32'hc40446e;
      2652: inst = 32'h8220000;
      2653: inst = 32'h10408000;
      2654: inst = 32'hc40446f;
      2655: inst = 32'h8220000;
      2656: inst = 32'h10408000;
      2657: inst = 32'hc404470;
      2658: inst = 32'h8220000;
      2659: inst = 32'h10408000;
      2660: inst = 32'hc404471;
      2661: inst = 32'h8220000;
      2662: inst = 32'h10408000;
      2663: inst = 32'hc404472;
      2664: inst = 32'h8220000;
      2665: inst = 32'h10408000;
      2666: inst = 32'hc404473;
      2667: inst = 32'h8220000;
      2668: inst = 32'h10408000;
      2669: inst = 32'hc404474;
      2670: inst = 32'h8220000;
      2671: inst = 32'h10408000;
      2672: inst = 32'hc404475;
      2673: inst = 32'h8220000;
      2674: inst = 32'h10408000;
      2675: inst = 32'hc404476;
      2676: inst = 32'h8220000;
      2677: inst = 32'h10408000;
      2678: inst = 32'hc404477;
      2679: inst = 32'h8220000;
      2680: inst = 32'h10408000;
      2681: inst = 32'hc404478;
      2682: inst = 32'h8220000;
      2683: inst = 32'h10408000;
      2684: inst = 32'hc404479;
      2685: inst = 32'h8220000;
      2686: inst = 32'h10408000;
      2687: inst = 32'hc40447a;
      2688: inst = 32'h8220000;
      2689: inst = 32'h10408000;
      2690: inst = 32'hc40447b;
      2691: inst = 32'h8220000;
      2692: inst = 32'h10408000;
      2693: inst = 32'hc4044a4;
      2694: inst = 32'h8220000;
      2695: inst = 32'h10408000;
      2696: inst = 32'hc4044a5;
      2697: inst = 32'h8220000;
      2698: inst = 32'h10408000;
      2699: inst = 32'hc4044a6;
      2700: inst = 32'h8220000;
      2701: inst = 32'h10408000;
      2702: inst = 32'hc4044a7;
      2703: inst = 32'h8220000;
      2704: inst = 32'h10408000;
      2705: inst = 32'hc4044a8;
      2706: inst = 32'h8220000;
      2707: inst = 32'h10408000;
      2708: inst = 32'hc4044a9;
      2709: inst = 32'h8220000;
      2710: inst = 32'h10408000;
      2711: inst = 32'hc4044aa;
      2712: inst = 32'h8220000;
      2713: inst = 32'h10408000;
      2714: inst = 32'hc4044ab;
      2715: inst = 32'h8220000;
      2716: inst = 32'h10408000;
      2717: inst = 32'hc4044ac;
      2718: inst = 32'h8220000;
      2719: inst = 32'h10408000;
      2720: inst = 32'hc4044ad;
      2721: inst = 32'h8220000;
      2722: inst = 32'h10408000;
      2723: inst = 32'hc4044ae;
      2724: inst = 32'h8220000;
      2725: inst = 32'h10408000;
      2726: inst = 32'hc4044af;
      2727: inst = 32'h8220000;
      2728: inst = 32'h10408000;
      2729: inst = 32'hc4044b0;
      2730: inst = 32'h8220000;
      2731: inst = 32'h10408000;
      2732: inst = 32'hc4044b1;
      2733: inst = 32'h8220000;
      2734: inst = 32'h10408000;
      2735: inst = 32'hc4044b6;
      2736: inst = 32'h8220000;
      2737: inst = 32'h10408000;
      2738: inst = 32'hc4044b7;
      2739: inst = 32'h8220000;
      2740: inst = 32'h10408000;
      2741: inst = 32'hc4044b8;
      2742: inst = 32'h8220000;
      2743: inst = 32'h10408000;
      2744: inst = 32'hc4044b9;
      2745: inst = 32'h8220000;
      2746: inst = 32'h10408000;
      2747: inst = 32'hc4044ba;
      2748: inst = 32'h8220000;
      2749: inst = 32'h10408000;
      2750: inst = 32'hc4044bb;
      2751: inst = 32'h8220000;
      2752: inst = 32'h10408000;
      2753: inst = 32'hc4044bc;
      2754: inst = 32'h8220000;
      2755: inst = 32'h10408000;
      2756: inst = 32'hc4044bd;
      2757: inst = 32'h8220000;
      2758: inst = 32'h10408000;
      2759: inst = 32'hc4044be;
      2760: inst = 32'h8220000;
      2761: inst = 32'h10408000;
      2762: inst = 32'hc4044bf;
      2763: inst = 32'h8220000;
      2764: inst = 32'h10408000;
      2765: inst = 32'hc4044c0;
      2766: inst = 32'h8220000;
      2767: inst = 32'h10408000;
      2768: inst = 32'hc4044c1;
      2769: inst = 32'h8220000;
      2770: inst = 32'h10408000;
      2771: inst = 32'hc4044c2;
      2772: inst = 32'h8220000;
      2773: inst = 32'h10408000;
      2774: inst = 32'hc4044c3;
      2775: inst = 32'h8220000;
      2776: inst = 32'h10408000;
      2777: inst = 32'hc4044c4;
      2778: inst = 32'h8220000;
      2779: inst = 32'h10408000;
      2780: inst = 32'hc4044c5;
      2781: inst = 32'h8220000;
      2782: inst = 32'h10408000;
      2783: inst = 32'hc4044c6;
      2784: inst = 32'h8220000;
      2785: inst = 32'h10408000;
      2786: inst = 32'hc4044c7;
      2787: inst = 32'h8220000;
      2788: inst = 32'h10408000;
      2789: inst = 32'hc4044c8;
      2790: inst = 32'h8220000;
      2791: inst = 32'h10408000;
      2792: inst = 32'hc4044c9;
      2793: inst = 32'h8220000;
      2794: inst = 32'h10408000;
      2795: inst = 32'hc4044ca;
      2796: inst = 32'h8220000;
      2797: inst = 32'h10408000;
      2798: inst = 32'hc4044cd;
      2799: inst = 32'h8220000;
      2800: inst = 32'h10408000;
      2801: inst = 32'hc4044ce;
      2802: inst = 32'h8220000;
      2803: inst = 32'h10408000;
      2804: inst = 32'hc4044cf;
      2805: inst = 32'h8220000;
      2806: inst = 32'h10408000;
      2807: inst = 32'hc4044d0;
      2808: inst = 32'h8220000;
      2809: inst = 32'h10408000;
      2810: inst = 32'hc4044d1;
      2811: inst = 32'h8220000;
      2812: inst = 32'h10408000;
      2813: inst = 32'hc4044d2;
      2814: inst = 32'h8220000;
      2815: inst = 32'h10408000;
      2816: inst = 32'hc4044d3;
      2817: inst = 32'h8220000;
      2818: inst = 32'h10408000;
      2819: inst = 32'hc4044d4;
      2820: inst = 32'h8220000;
      2821: inst = 32'h10408000;
      2822: inst = 32'hc4044d5;
      2823: inst = 32'h8220000;
      2824: inst = 32'h10408000;
      2825: inst = 32'hc4044d6;
      2826: inst = 32'h8220000;
      2827: inst = 32'h10408000;
      2828: inst = 32'hc4044d7;
      2829: inst = 32'h8220000;
      2830: inst = 32'h10408000;
      2831: inst = 32'hc4044d8;
      2832: inst = 32'h8220000;
      2833: inst = 32'h10408000;
      2834: inst = 32'hc4044d9;
      2835: inst = 32'h8220000;
      2836: inst = 32'h10408000;
      2837: inst = 32'hc4044da;
      2838: inst = 32'h8220000;
      2839: inst = 32'h10408000;
      2840: inst = 32'hc4044db;
      2841: inst = 32'h8220000;
      2842: inst = 32'h10408000;
      2843: inst = 32'hc404504;
      2844: inst = 32'h8220000;
      2845: inst = 32'h10408000;
      2846: inst = 32'hc404505;
      2847: inst = 32'h8220000;
      2848: inst = 32'h10408000;
      2849: inst = 32'hc404506;
      2850: inst = 32'h8220000;
      2851: inst = 32'h10408000;
      2852: inst = 32'hc404507;
      2853: inst = 32'h8220000;
      2854: inst = 32'h10408000;
      2855: inst = 32'hc404508;
      2856: inst = 32'h8220000;
      2857: inst = 32'h10408000;
      2858: inst = 32'hc404509;
      2859: inst = 32'h8220000;
      2860: inst = 32'h10408000;
      2861: inst = 32'hc40450a;
      2862: inst = 32'h8220000;
      2863: inst = 32'h10408000;
      2864: inst = 32'hc40450b;
      2865: inst = 32'h8220000;
      2866: inst = 32'h10408000;
      2867: inst = 32'hc40450c;
      2868: inst = 32'h8220000;
      2869: inst = 32'h10408000;
      2870: inst = 32'hc40450d;
      2871: inst = 32'h8220000;
      2872: inst = 32'h10408000;
      2873: inst = 32'hc40450e;
      2874: inst = 32'h8220000;
      2875: inst = 32'h10408000;
      2876: inst = 32'hc40450f;
      2877: inst = 32'h8220000;
      2878: inst = 32'h10408000;
      2879: inst = 32'hc404510;
      2880: inst = 32'h8220000;
      2881: inst = 32'h10408000;
      2882: inst = 32'hc404511;
      2883: inst = 32'h8220000;
      2884: inst = 32'h10408000;
      2885: inst = 32'hc404512;
      2886: inst = 32'h8220000;
      2887: inst = 32'h10408000;
      2888: inst = 32'hc404515;
      2889: inst = 32'h8220000;
      2890: inst = 32'h10408000;
      2891: inst = 32'hc404516;
      2892: inst = 32'h8220000;
      2893: inst = 32'h10408000;
      2894: inst = 32'hc404517;
      2895: inst = 32'h8220000;
      2896: inst = 32'h10408000;
      2897: inst = 32'hc404518;
      2898: inst = 32'h8220000;
      2899: inst = 32'h10408000;
      2900: inst = 32'hc404519;
      2901: inst = 32'h8220000;
      2902: inst = 32'h10408000;
      2903: inst = 32'hc40451a;
      2904: inst = 32'h8220000;
      2905: inst = 32'h10408000;
      2906: inst = 32'hc40451b;
      2907: inst = 32'h8220000;
      2908: inst = 32'h10408000;
      2909: inst = 32'hc40451c;
      2910: inst = 32'h8220000;
      2911: inst = 32'h10408000;
      2912: inst = 32'hc40451d;
      2913: inst = 32'h8220000;
      2914: inst = 32'h10408000;
      2915: inst = 32'hc40451e;
      2916: inst = 32'h8220000;
      2917: inst = 32'h10408000;
      2918: inst = 32'hc40451f;
      2919: inst = 32'h8220000;
      2920: inst = 32'h10408000;
      2921: inst = 32'hc404520;
      2922: inst = 32'h8220000;
      2923: inst = 32'h10408000;
      2924: inst = 32'hc404521;
      2925: inst = 32'h8220000;
      2926: inst = 32'h10408000;
      2927: inst = 32'hc404522;
      2928: inst = 32'h8220000;
      2929: inst = 32'h10408000;
      2930: inst = 32'hc404523;
      2931: inst = 32'h8220000;
      2932: inst = 32'h10408000;
      2933: inst = 32'hc404524;
      2934: inst = 32'h8220000;
      2935: inst = 32'h10408000;
      2936: inst = 32'hc404525;
      2937: inst = 32'h8220000;
      2938: inst = 32'h10408000;
      2939: inst = 32'hc404526;
      2940: inst = 32'h8220000;
      2941: inst = 32'h10408000;
      2942: inst = 32'hc404527;
      2943: inst = 32'h8220000;
      2944: inst = 32'h10408000;
      2945: inst = 32'hc404528;
      2946: inst = 32'h8220000;
      2947: inst = 32'h10408000;
      2948: inst = 32'hc404529;
      2949: inst = 32'h8220000;
      2950: inst = 32'h10408000;
      2951: inst = 32'hc40452a;
      2952: inst = 32'h8220000;
      2953: inst = 32'h10408000;
      2954: inst = 32'hc40452b;
      2955: inst = 32'h8220000;
      2956: inst = 32'h10408000;
      2957: inst = 32'hc40452c;
      2958: inst = 32'h8220000;
      2959: inst = 32'h10408000;
      2960: inst = 32'hc40452d;
      2961: inst = 32'h8220000;
      2962: inst = 32'h10408000;
      2963: inst = 32'hc40452e;
      2964: inst = 32'h8220000;
      2965: inst = 32'h10408000;
      2966: inst = 32'hc40452f;
      2967: inst = 32'h8220000;
      2968: inst = 32'h10408000;
      2969: inst = 32'hc404530;
      2970: inst = 32'h8220000;
      2971: inst = 32'h10408000;
      2972: inst = 32'hc404531;
      2973: inst = 32'h8220000;
      2974: inst = 32'h10408000;
      2975: inst = 32'hc404532;
      2976: inst = 32'h8220000;
      2977: inst = 32'h10408000;
      2978: inst = 32'hc404533;
      2979: inst = 32'h8220000;
      2980: inst = 32'h10408000;
      2981: inst = 32'hc404534;
      2982: inst = 32'h8220000;
      2983: inst = 32'h10408000;
      2984: inst = 32'hc404535;
      2985: inst = 32'h8220000;
      2986: inst = 32'h10408000;
      2987: inst = 32'hc404536;
      2988: inst = 32'h8220000;
      2989: inst = 32'h10408000;
      2990: inst = 32'hc404537;
      2991: inst = 32'h8220000;
      2992: inst = 32'h10408000;
      2993: inst = 32'hc404538;
      2994: inst = 32'h8220000;
      2995: inst = 32'h10408000;
      2996: inst = 32'hc404539;
      2997: inst = 32'h8220000;
      2998: inst = 32'h10408000;
      2999: inst = 32'hc40453a;
      3000: inst = 32'h8220000;
      3001: inst = 32'h10408000;
      3002: inst = 32'hc40453b;
      3003: inst = 32'h8220000;
      3004: inst = 32'h10408000;
      3005: inst = 32'hc404564;
      3006: inst = 32'h8220000;
      3007: inst = 32'h10408000;
      3008: inst = 32'hc404565;
      3009: inst = 32'h8220000;
      3010: inst = 32'h10408000;
      3011: inst = 32'hc404566;
      3012: inst = 32'h8220000;
      3013: inst = 32'h10408000;
      3014: inst = 32'hc404567;
      3015: inst = 32'h8220000;
      3016: inst = 32'h10408000;
      3017: inst = 32'hc404568;
      3018: inst = 32'h8220000;
      3019: inst = 32'h10408000;
      3020: inst = 32'hc404569;
      3021: inst = 32'h8220000;
      3022: inst = 32'h10408000;
      3023: inst = 32'hc40456a;
      3024: inst = 32'h8220000;
      3025: inst = 32'h10408000;
      3026: inst = 32'hc40456b;
      3027: inst = 32'h8220000;
      3028: inst = 32'h10408000;
      3029: inst = 32'hc40456c;
      3030: inst = 32'h8220000;
      3031: inst = 32'h10408000;
      3032: inst = 32'hc40456d;
      3033: inst = 32'h8220000;
      3034: inst = 32'h10408000;
      3035: inst = 32'hc40456e;
      3036: inst = 32'h8220000;
      3037: inst = 32'h10408000;
      3038: inst = 32'hc40456f;
      3039: inst = 32'h8220000;
      3040: inst = 32'h10408000;
      3041: inst = 32'hc404570;
      3042: inst = 32'h8220000;
      3043: inst = 32'h10408000;
      3044: inst = 32'hc404571;
      3045: inst = 32'h8220000;
      3046: inst = 32'h10408000;
      3047: inst = 32'hc404572;
      3048: inst = 32'h8220000;
      3049: inst = 32'h10408000;
      3050: inst = 32'hc404573;
      3051: inst = 32'h8220000;
      3052: inst = 32'h10408000;
      3053: inst = 32'hc404574;
      3054: inst = 32'h8220000;
      3055: inst = 32'h10408000;
      3056: inst = 32'hc404575;
      3057: inst = 32'h8220000;
      3058: inst = 32'h10408000;
      3059: inst = 32'hc404576;
      3060: inst = 32'h8220000;
      3061: inst = 32'h10408000;
      3062: inst = 32'hc404577;
      3063: inst = 32'h8220000;
      3064: inst = 32'h10408000;
      3065: inst = 32'hc404578;
      3066: inst = 32'h8220000;
      3067: inst = 32'h10408000;
      3068: inst = 32'hc404579;
      3069: inst = 32'h8220000;
      3070: inst = 32'h10408000;
      3071: inst = 32'hc40457a;
      3072: inst = 32'h8220000;
      3073: inst = 32'h10408000;
      3074: inst = 32'hc40457b;
      3075: inst = 32'h8220000;
      3076: inst = 32'h10408000;
      3077: inst = 32'hc40457c;
      3078: inst = 32'h8220000;
      3079: inst = 32'h10408000;
      3080: inst = 32'hc40457d;
      3081: inst = 32'h8220000;
      3082: inst = 32'h10408000;
      3083: inst = 32'hc40457e;
      3084: inst = 32'h8220000;
      3085: inst = 32'h10408000;
      3086: inst = 32'hc40457f;
      3087: inst = 32'h8220000;
      3088: inst = 32'h10408000;
      3089: inst = 32'hc404580;
      3090: inst = 32'h8220000;
      3091: inst = 32'h10408000;
      3092: inst = 32'hc404581;
      3093: inst = 32'h8220000;
      3094: inst = 32'h10408000;
      3095: inst = 32'hc404582;
      3096: inst = 32'h8220000;
      3097: inst = 32'h10408000;
      3098: inst = 32'hc404583;
      3099: inst = 32'h8220000;
      3100: inst = 32'h10408000;
      3101: inst = 32'hc404584;
      3102: inst = 32'h8220000;
      3103: inst = 32'h10408000;
      3104: inst = 32'hc404585;
      3105: inst = 32'h8220000;
      3106: inst = 32'h10408000;
      3107: inst = 32'hc404586;
      3108: inst = 32'h8220000;
      3109: inst = 32'h10408000;
      3110: inst = 32'hc404587;
      3111: inst = 32'h8220000;
      3112: inst = 32'h10408000;
      3113: inst = 32'hc404588;
      3114: inst = 32'h8220000;
      3115: inst = 32'h10408000;
      3116: inst = 32'hc404589;
      3117: inst = 32'h8220000;
      3118: inst = 32'h10408000;
      3119: inst = 32'hc40458a;
      3120: inst = 32'h8220000;
      3121: inst = 32'h10408000;
      3122: inst = 32'hc40458b;
      3123: inst = 32'h8220000;
      3124: inst = 32'h10408000;
      3125: inst = 32'hc40458c;
      3126: inst = 32'h8220000;
      3127: inst = 32'h10408000;
      3128: inst = 32'hc40458d;
      3129: inst = 32'h8220000;
      3130: inst = 32'h10408000;
      3131: inst = 32'hc40458e;
      3132: inst = 32'h8220000;
      3133: inst = 32'h10408000;
      3134: inst = 32'hc40458f;
      3135: inst = 32'h8220000;
      3136: inst = 32'h10408000;
      3137: inst = 32'hc404590;
      3138: inst = 32'h8220000;
      3139: inst = 32'h10408000;
      3140: inst = 32'hc404591;
      3141: inst = 32'h8220000;
      3142: inst = 32'h10408000;
      3143: inst = 32'hc404592;
      3144: inst = 32'h8220000;
      3145: inst = 32'h10408000;
      3146: inst = 32'hc404593;
      3147: inst = 32'h8220000;
      3148: inst = 32'h10408000;
      3149: inst = 32'hc404594;
      3150: inst = 32'h8220000;
      3151: inst = 32'h10408000;
      3152: inst = 32'hc404595;
      3153: inst = 32'h8220000;
      3154: inst = 32'h10408000;
      3155: inst = 32'hc404596;
      3156: inst = 32'h8220000;
      3157: inst = 32'h10408000;
      3158: inst = 32'hc404597;
      3159: inst = 32'h8220000;
      3160: inst = 32'h10408000;
      3161: inst = 32'hc404598;
      3162: inst = 32'h8220000;
      3163: inst = 32'h10408000;
      3164: inst = 32'hc404599;
      3165: inst = 32'h8220000;
      3166: inst = 32'h10408000;
      3167: inst = 32'hc40459a;
      3168: inst = 32'h8220000;
      3169: inst = 32'h10408000;
      3170: inst = 32'hc40459b;
      3171: inst = 32'h8220000;
      3172: inst = 32'h10408000;
      3173: inst = 32'hc4045c4;
      3174: inst = 32'h8220000;
      3175: inst = 32'h10408000;
      3176: inst = 32'hc4045c5;
      3177: inst = 32'h8220000;
      3178: inst = 32'h10408000;
      3179: inst = 32'hc4045c6;
      3180: inst = 32'h8220000;
      3181: inst = 32'h10408000;
      3182: inst = 32'hc4045c7;
      3183: inst = 32'h8220000;
      3184: inst = 32'h10408000;
      3185: inst = 32'hc4045c8;
      3186: inst = 32'h8220000;
      3187: inst = 32'h10408000;
      3188: inst = 32'hc4045c9;
      3189: inst = 32'h8220000;
      3190: inst = 32'h10408000;
      3191: inst = 32'hc4045ca;
      3192: inst = 32'h8220000;
      3193: inst = 32'h10408000;
      3194: inst = 32'hc4045cb;
      3195: inst = 32'h8220000;
      3196: inst = 32'h10408000;
      3197: inst = 32'hc4045cc;
      3198: inst = 32'h8220000;
      3199: inst = 32'h10408000;
      3200: inst = 32'hc4045cd;
      3201: inst = 32'h8220000;
      3202: inst = 32'h10408000;
      3203: inst = 32'hc4045ce;
      3204: inst = 32'h8220000;
      3205: inst = 32'h10408000;
      3206: inst = 32'hc4045cf;
      3207: inst = 32'h8220000;
      3208: inst = 32'h10408000;
      3209: inst = 32'hc4045d0;
      3210: inst = 32'h8220000;
      3211: inst = 32'h10408000;
      3212: inst = 32'hc4045d1;
      3213: inst = 32'h8220000;
      3214: inst = 32'h10408000;
      3215: inst = 32'hc4045d2;
      3216: inst = 32'h8220000;
      3217: inst = 32'h10408000;
      3218: inst = 32'hc4045d3;
      3219: inst = 32'h8220000;
      3220: inst = 32'h10408000;
      3221: inst = 32'hc4045d4;
      3222: inst = 32'h8220000;
      3223: inst = 32'h10408000;
      3224: inst = 32'hc4045d5;
      3225: inst = 32'h8220000;
      3226: inst = 32'h10408000;
      3227: inst = 32'hc4045d6;
      3228: inst = 32'h8220000;
      3229: inst = 32'h10408000;
      3230: inst = 32'hc4045d7;
      3231: inst = 32'h8220000;
      3232: inst = 32'h10408000;
      3233: inst = 32'hc4045d8;
      3234: inst = 32'h8220000;
      3235: inst = 32'h10408000;
      3236: inst = 32'hc4045d9;
      3237: inst = 32'h8220000;
      3238: inst = 32'h10408000;
      3239: inst = 32'hc4045da;
      3240: inst = 32'h8220000;
      3241: inst = 32'h10408000;
      3242: inst = 32'hc4045db;
      3243: inst = 32'h8220000;
      3244: inst = 32'h10408000;
      3245: inst = 32'hc4045dc;
      3246: inst = 32'h8220000;
      3247: inst = 32'h10408000;
      3248: inst = 32'hc4045dd;
      3249: inst = 32'h8220000;
      3250: inst = 32'h10408000;
      3251: inst = 32'hc4045de;
      3252: inst = 32'h8220000;
      3253: inst = 32'h10408000;
      3254: inst = 32'hc4045df;
      3255: inst = 32'h8220000;
      3256: inst = 32'h10408000;
      3257: inst = 32'hc4045e0;
      3258: inst = 32'h8220000;
      3259: inst = 32'h10408000;
      3260: inst = 32'hc4045e1;
      3261: inst = 32'h8220000;
      3262: inst = 32'h10408000;
      3263: inst = 32'hc4045e2;
      3264: inst = 32'h8220000;
      3265: inst = 32'h10408000;
      3266: inst = 32'hc4045e3;
      3267: inst = 32'h8220000;
      3268: inst = 32'h10408000;
      3269: inst = 32'hc4045e4;
      3270: inst = 32'h8220000;
      3271: inst = 32'h10408000;
      3272: inst = 32'hc4045e5;
      3273: inst = 32'h8220000;
      3274: inst = 32'h10408000;
      3275: inst = 32'hc4045e6;
      3276: inst = 32'h8220000;
      3277: inst = 32'h10408000;
      3278: inst = 32'hc4045e7;
      3279: inst = 32'h8220000;
      3280: inst = 32'h10408000;
      3281: inst = 32'hc4045e8;
      3282: inst = 32'h8220000;
      3283: inst = 32'h10408000;
      3284: inst = 32'hc4045e9;
      3285: inst = 32'h8220000;
      3286: inst = 32'h10408000;
      3287: inst = 32'hc4045ea;
      3288: inst = 32'h8220000;
      3289: inst = 32'h10408000;
      3290: inst = 32'hc4045eb;
      3291: inst = 32'h8220000;
      3292: inst = 32'h10408000;
      3293: inst = 32'hc4045ec;
      3294: inst = 32'h8220000;
      3295: inst = 32'h10408000;
      3296: inst = 32'hc4045ed;
      3297: inst = 32'h8220000;
      3298: inst = 32'h10408000;
      3299: inst = 32'hc4045ee;
      3300: inst = 32'h8220000;
      3301: inst = 32'h10408000;
      3302: inst = 32'hc4045ef;
      3303: inst = 32'h8220000;
      3304: inst = 32'h10408000;
      3305: inst = 32'hc4045f0;
      3306: inst = 32'h8220000;
      3307: inst = 32'h10408000;
      3308: inst = 32'hc4045f1;
      3309: inst = 32'h8220000;
      3310: inst = 32'h10408000;
      3311: inst = 32'hc4045f2;
      3312: inst = 32'h8220000;
      3313: inst = 32'h10408000;
      3314: inst = 32'hc4045f3;
      3315: inst = 32'h8220000;
      3316: inst = 32'h10408000;
      3317: inst = 32'hc4045f4;
      3318: inst = 32'h8220000;
      3319: inst = 32'h10408000;
      3320: inst = 32'hc4045f5;
      3321: inst = 32'h8220000;
      3322: inst = 32'h10408000;
      3323: inst = 32'hc4045f6;
      3324: inst = 32'h8220000;
      3325: inst = 32'h10408000;
      3326: inst = 32'hc4045f7;
      3327: inst = 32'h8220000;
      3328: inst = 32'h10408000;
      3329: inst = 32'hc4045f8;
      3330: inst = 32'h8220000;
      3331: inst = 32'h10408000;
      3332: inst = 32'hc4045f9;
      3333: inst = 32'h8220000;
      3334: inst = 32'h10408000;
      3335: inst = 32'hc4045fa;
      3336: inst = 32'h8220000;
      3337: inst = 32'h10408000;
      3338: inst = 32'hc4045fb;
      3339: inst = 32'h8220000;
      3340: inst = 32'h10408000;
      3341: inst = 32'hc404624;
      3342: inst = 32'h8220000;
      3343: inst = 32'h10408000;
      3344: inst = 32'hc404625;
      3345: inst = 32'h8220000;
      3346: inst = 32'h10408000;
      3347: inst = 32'hc404626;
      3348: inst = 32'h8220000;
      3349: inst = 32'h10408000;
      3350: inst = 32'hc404627;
      3351: inst = 32'h8220000;
      3352: inst = 32'h10408000;
      3353: inst = 32'hc404628;
      3354: inst = 32'h8220000;
      3355: inst = 32'h10408000;
      3356: inst = 32'hc404629;
      3357: inst = 32'h8220000;
      3358: inst = 32'h10408000;
      3359: inst = 32'hc40462a;
      3360: inst = 32'h8220000;
      3361: inst = 32'h10408000;
      3362: inst = 32'hc40462b;
      3363: inst = 32'h8220000;
      3364: inst = 32'h10408000;
      3365: inst = 32'hc40462c;
      3366: inst = 32'h8220000;
      3367: inst = 32'h10408000;
      3368: inst = 32'hc40462d;
      3369: inst = 32'h8220000;
      3370: inst = 32'h10408000;
      3371: inst = 32'hc40462e;
      3372: inst = 32'h8220000;
      3373: inst = 32'h10408000;
      3374: inst = 32'hc40462f;
      3375: inst = 32'h8220000;
      3376: inst = 32'h10408000;
      3377: inst = 32'hc404630;
      3378: inst = 32'h8220000;
      3379: inst = 32'h10408000;
      3380: inst = 32'hc404631;
      3381: inst = 32'h8220000;
      3382: inst = 32'h10408000;
      3383: inst = 32'hc404632;
      3384: inst = 32'h8220000;
      3385: inst = 32'h10408000;
      3386: inst = 32'hc404633;
      3387: inst = 32'h8220000;
      3388: inst = 32'h10408000;
      3389: inst = 32'hc404634;
      3390: inst = 32'h8220000;
      3391: inst = 32'h10408000;
      3392: inst = 32'hc404635;
      3393: inst = 32'h8220000;
      3394: inst = 32'h10408000;
      3395: inst = 32'hc404636;
      3396: inst = 32'h8220000;
      3397: inst = 32'h10408000;
      3398: inst = 32'hc404637;
      3399: inst = 32'h8220000;
      3400: inst = 32'h10408000;
      3401: inst = 32'hc404638;
      3402: inst = 32'h8220000;
      3403: inst = 32'h10408000;
      3404: inst = 32'hc404639;
      3405: inst = 32'h8220000;
      3406: inst = 32'h10408000;
      3407: inst = 32'hc40463a;
      3408: inst = 32'h8220000;
      3409: inst = 32'h10408000;
      3410: inst = 32'hc40463b;
      3411: inst = 32'h8220000;
      3412: inst = 32'h10408000;
      3413: inst = 32'hc40463c;
      3414: inst = 32'h8220000;
      3415: inst = 32'h10408000;
      3416: inst = 32'hc40463d;
      3417: inst = 32'h8220000;
      3418: inst = 32'h10408000;
      3419: inst = 32'hc40463e;
      3420: inst = 32'h8220000;
      3421: inst = 32'h10408000;
      3422: inst = 32'hc40463f;
      3423: inst = 32'h8220000;
      3424: inst = 32'h10408000;
      3425: inst = 32'hc404640;
      3426: inst = 32'h8220000;
      3427: inst = 32'h10408000;
      3428: inst = 32'hc404641;
      3429: inst = 32'h8220000;
      3430: inst = 32'h10408000;
      3431: inst = 32'hc404642;
      3432: inst = 32'h8220000;
      3433: inst = 32'h10408000;
      3434: inst = 32'hc404643;
      3435: inst = 32'h8220000;
      3436: inst = 32'h10408000;
      3437: inst = 32'hc404644;
      3438: inst = 32'h8220000;
      3439: inst = 32'h10408000;
      3440: inst = 32'hc404645;
      3441: inst = 32'h8220000;
      3442: inst = 32'h10408000;
      3443: inst = 32'hc404646;
      3444: inst = 32'h8220000;
      3445: inst = 32'h10408000;
      3446: inst = 32'hc404647;
      3447: inst = 32'h8220000;
      3448: inst = 32'h10408000;
      3449: inst = 32'hc404648;
      3450: inst = 32'h8220000;
      3451: inst = 32'h10408000;
      3452: inst = 32'hc404649;
      3453: inst = 32'h8220000;
      3454: inst = 32'h10408000;
      3455: inst = 32'hc40464a;
      3456: inst = 32'h8220000;
      3457: inst = 32'h10408000;
      3458: inst = 32'hc40464b;
      3459: inst = 32'h8220000;
      3460: inst = 32'h10408000;
      3461: inst = 32'hc40464c;
      3462: inst = 32'h8220000;
      3463: inst = 32'h10408000;
      3464: inst = 32'hc40464d;
      3465: inst = 32'h8220000;
      3466: inst = 32'h10408000;
      3467: inst = 32'hc40464e;
      3468: inst = 32'h8220000;
      3469: inst = 32'h10408000;
      3470: inst = 32'hc40464f;
      3471: inst = 32'h8220000;
      3472: inst = 32'h10408000;
      3473: inst = 32'hc404650;
      3474: inst = 32'h8220000;
      3475: inst = 32'h10408000;
      3476: inst = 32'hc404651;
      3477: inst = 32'h8220000;
      3478: inst = 32'h10408000;
      3479: inst = 32'hc404652;
      3480: inst = 32'h8220000;
      3481: inst = 32'h10408000;
      3482: inst = 32'hc404653;
      3483: inst = 32'h8220000;
      3484: inst = 32'h10408000;
      3485: inst = 32'hc404654;
      3486: inst = 32'h8220000;
      3487: inst = 32'h10408000;
      3488: inst = 32'hc404655;
      3489: inst = 32'h8220000;
      3490: inst = 32'h10408000;
      3491: inst = 32'hc404656;
      3492: inst = 32'h8220000;
      3493: inst = 32'h10408000;
      3494: inst = 32'hc404657;
      3495: inst = 32'h8220000;
      3496: inst = 32'h10408000;
      3497: inst = 32'hc404658;
      3498: inst = 32'h8220000;
      3499: inst = 32'h10408000;
      3500: inst = 32'hc404659;
      3501: inst = 32'h8220000;
      3502: inst = 32'h10408000;
      3503: inst = 32'hc40465a;
      3504: inst = 32'h8220000;
      3505: inst = 32'h10408000;
      3506: inst = 32'hc40465b;
      3507: inst = 32'h8220000;
      3508: inst = 32'h10408000;
      3509: inst = 32'hc404684;
      3510: inst = 32'h8220000;
      3511: inst = 32'h10408000;
      3512: inst = 32'hc404685;
      3513: inst = 32'h8220000;
      3514: inst = 32'h10408000;
      3515: inst = 32'hc404686;
      3516: inst = 32'h8220000;
      3517: inst = 32'h10408000;
      3518: inst = 32'hc404687;
      3519: inst = 32'h8220000;
      3520: inst = 32'h10408000;
      3521: inst = 32'hc404688;
      3522: inst = 32'h8220000;
      3523: inst = 32'h10408000;
      3524: inst = 32'hc404689;
      3525: inst = 32'h8220000;
      3526: inst = 32'h10408000;
      3527: inst = 32'hc40468a;
      3528: inst = 32'h8220000;
      3529: inst = 32'h10408000;
      3530: inst = 32'hc40468b;
      3531: inst = 32'h8220000;
      3532: inst = 32'h10408000;
      3533: inst = 32'hc40468c;
      3534: inst = 32'h8220000;
      3535: inst = 32'h10408000;
      3536: inst = 32'hc40468d;
      3537: inst = 32'h8220000;
      3538: inst = 32'h10408000;
      3539: inst = 32'hc40468e;
      3540: inst = 32'h8220000;
      3541: inst = 32'h10408000;
      3542: inst = 32'hc40468f;
      3543: inst = 32'h8220000;
      3544: inst = 32'h10408000;
      3545: inst = 32'hc404690;
      3546: inst = 32'h8220000;
      3547: inst = 32'h10408000;
      3548: inst = 32'hc404691;
      3549: inst = 32'h8220000;
      3550: inst = 32'h10408000;
      3551: inst = 32'hc404692;
      3552: inst = 32'h8220000;
      3553: inst = 32'h10408000;
      3554: inst = 32'hc404693;
      3555: inst = 32'h8220000;
      3556: inst = 32'h10408000;
      3557: inst = 32'hc404694;
      3558: inst = 32'h8220000;
      3559: inst = 32'h10408000;
      3560: inst = 32'hc404695;
      3561: inst = 32'h8220000;
      3562: inst = 32'h10408000;
      3563: inst = 32'hc404696;
      3564: inst = 32'h8220000;
      3565: inst = 32'h10408000;
      3566: inst = 32'hc404697;
      3567: inst = 32'h8220000;
      3568: inst = 32'h10408000;
      3569: inst = 32'hc404698;
      3570: inst = 32'h8220000;
      3571: inst = 32'h10408000;
      3572: inst = 32'hc404699;
      3573: inst = 32'h8220000;
      3574: inst = 32'h10408000;
      3575: inst = 32'hc40469a;
      3576: inst = 32'h8220000;
      3577: inst = 32'h10408000;
      3578: inst = 32'hc40469b;
      3579: inst = 32'h8220000;
      3580: inst = 32'h10408000;
      3581: inst = 32'hc40469c;
      3582: inst = 32'h8220000;
      3583: inst = 32'h10408000;
      3584: inst = 32'hc40469d;
      3585: inst = 32'h8220000;
      3586: inst = 32'h10408000;
      3587: inst = 32'hc40469e;
      3588: inst = 32'h8220000;
      3589: inst = 32'h10408000;
      3590: inst = 32'hc40469f;
      3591: inst = 32'h8220000;
      3592: inst = 32'h10408000;
      3593: inst = 32'hc4046a0;
      3594: inst = 32'h8220000;
      3595: inst = 32'h10408000;
      3596: inst = 32'hc4046a1;
      3597: inst = 32'h8220000;
      3598: inst = 32'h10408000;
      3599: inst = 32'hc4046a2;
      3600: inst = 32'h8220000;
      3601: inst = 32'h10408000;
      3602: inst = 32'hc4046a3;
      3603: inst = 32'h8220000;
      3604: inst = 32'h10408000;
      3605: inst = 32'hc4046a4;
      3606: inst = 32'h8220000;
      3607: inst = 32'h10408000;
      3608: inst = 32'hc4046a5;
      3609: inst = 32'h8220000;
      3610: inst = 32'h10408000;
      3611: inst = 32'hc4046a6;
      3612: inst = 32'h8220000;
      3613: inst = 32'h10408000;
      3614: inst = 32'hc4046a7;
      3615: inst = 32'h8220000;
      3616: inst = 32'h10408000;
      3617: inst = 32'hc4046a8;
      3618: inst = 32'h8220000;
      3619: inst = 32'h10408000;
      3620: inst = 32'hc4046a9;
      3621: inst = 32'h8220000;
      3622: inst = 32'h10408000;
      3623: inst = 32'hc4046aa;
      3624: inst = 32'h8220000;
      3625: inst = 32'h10408000;
      3626: inst = 32'hc4046ab;
      3627: inst = 32'h8220000;
      3628: inst = 32'h10408000;
      3629: inst = 32'hc4046ac;
      3630: inst = 32'h8220000;
      3631: inst = 32'h10408000;
      3632: inst = 32'hc4046ad;
      3633: inst = 32'h8220000;
      3634: inst = 32'h10408000;
      3635: inst = 32'hc4046ae;
      3636: inst = 32'h8220000;
      3637: inst = 32'h10408000;
      3638: inst = 32'hc4046af;
      3639: inst = 32'h8220000;
      3640: inst = 32'h10408000;
      3641: inst = 32'hc4046b0;
      3642: inst = 32'h8220000;
      3643: inst = 32'h10408000;
      3644: inst = 32'hc4046b1;
      3645: inst = 32'h8220000;
      3646: inst = 32'h10408000;
      3647: inst = 32'hc4046b2;
      3648: inst = 32'h8220000;
      3649: inst = 32'h10408000;
      3650: inst = 32'hc4046b3;
      3651: inst = 32'h8220000;
      3652: inst = 32'h10408000;
      3653: inst = 32'hc4046b4;
      3654: inst = 32'h8220000;
      3655: inst = 32'h10408000;
      3656: inst = 32'hc4046b5;
      3657: inst = 32'h8220000;
      3658: inst = 32'h10408000;
      3659: inst = 32'hc4046b6;
      3660: inst = 32'h8220000;
      3661: inst = 32'h10408000;
      3662: inst = 32'hc4046b7;
      3663: inst = 32'h8220000;
      3664: inst = 32'h10408000;
      3665: inst = 32'hc4046b8;
      3666: inst = 32'h8220000;
      3667: inst = 32'h10408000;
      3668: inst = 32'hc4046b9;
      3669: inst = 32'h8220000;
      3670: inst = 32'h10408000;
      3671: inst = 32'hc4046ba;
      3672: inst = 32'h8220000;
      3673: inst = 32'h10408000;
      3674: inst = 32'hc4046bb;
      3675: inst = 32'h8220000;
      3676: inst = 32'h10408000;
      3677: inst = 32'hc4046e4;
      3678: inst = 32'h8220000;
      3679: inst = 32'h10408000;
      3680: inst = 32'hc4046e5;
      3681: inst = 32'h8220000;
      3682: inst = 32'h10408000;
      3683: inst = 32'hc4046e6;
      3684: inst = 32'h8220000;
      3685: inst = 32'h10408000;
      3686: inst = 32'hc4046e7;
      3687: inst = 32'h8220000;
      3688: inst = 32'h10408000;
      3689: inst = 32'hc4046e8;
      3690: inst = 32'h8220000;
      3691: inst = 32'h10408000;
      3692: inst = 32'hc4046e9;
      3693: inst = 32'h8220000;
      3694: inst = 32'h10408000;
      3695: inst = 32'hc4046ea;
      3696: inst = 32'h8220000;
      3697: inst = 32'h10408000;
      3698: inst = 32'hc4046eb;
      3699: inst = 32'h8220000;
      3700: inst = 32'h10408000;
      3701: inst = 32'hc4046ec;
      3702: inst = 32'h8220000;
      3703: inst = 32'h10408000;
      3704: inst = 32'hc4046ed;
      3705: inst = 32'h8220000;
      3706: inst = 32'h10408000;
      3707: inst = 32'hc4046ee;
      3708: inst = 32'h8220000;
      3709: inst = 32'h10408000;
      3710: inst = 32'hc404700;
      3711: inst = 32'h8220000;
      3712: inst = 32'h10408000;
      3713: inst = 32'hc404701;
      3714: inst = 32'h8220000;
      3715: inst = 32'h10408000;
      3716: inst = 32'hc404702;
      3717: inst = 32'h8220000;
      3718: inst = 32'h10408000;
      3719: inst = 32'hc404703;
      3720: inst = 32'h8220000;
      3721: inst = 32'h10408000;
      3722: inst = 32'hc404704;
      3723: inst = 32'h8220000;
      3724: inst = 32'h10408000;
      3725: inst = 32'hc404705;
      3726: inst = 32'h8220000;
      3727: inst = 32'h10408000;
      3728: inst = 32'hc404706;
      3729: inst = 32'h8220000;
      3730: inst = 32'h10408000;
      3731: inst = 32'hc404707;
      3732: inst = 32'h8220000;
      3733: inst = 32'h10408000;
      3734: inst = 32'hc404708;
      3735: inst = 32'h8220000;
      3736: inst = 32'h10408000;
      3737: inst = 32'hc404709;
      3738: inst = 32'h8220000;
      3739: inst = 32'h10408000;
      3740: inst = 32'hc40470a;
      3741: inst = 32'h8220000;
      3742: inst = 32'h10408000;
      3743: inst = 32'hc40470b;
      3744: inst = 32'h8220000;
      3745: inst = 32'h10408000;
      3746: inst = 32'hc40470c;
      3747: inst = 32'h8220000;
      3748: inst = 32'h10408000;
      3749: inst = 32'hc40470d;
      3750: inst = 32'h8220000;
      3751: inst = 32'h10408000;
      3752: inst = 32'hc40470e;
      3753: inst = 32'h8220000;
      3754: inst = 32'h10408000;
      3755: inst = 32'hc40470f;
      3756: inst = 32'h8220000;
      3757: inst = 32'h10408000;
      3758: inst = 32'hc404710;
      3759: inst = 32'h8220000;
      3760: inst = 32'h10408000;
      3761: inst = 32'hc404711;
      3762: inst = 32'h8220000;
      3763: inst = 32'h10408000;
      3764: inst = 32'hc404712;
      3765: inst = 32'h8220000;
      3766: inst = 32'h10408000;
      3767: inst = 32'hc404713;
      3768: inst = 32'h8220000;
      3769: inst = 32'h10408000;
      3770: inst = 32'hc404714;
      3771: inst = 32'h8220000;
      3772: inst = 32'h10408000;
      3773: inst = 32'hc404715;
      3774: inst = 32'h8220000;
      3775: inst = 32'h10408000;
      3776: inst = 32'hc404716;
      3777: inst = 32'h8220000;
      3778: inst = 32'h10408000;
      3779: inst = 32'hc404717;
      3780: inst = 32'h8220000;
      3781: inst = 32'h10408000;
      3782: inst = 32'hc404718;
      3783: inst = 32'h8220000;
      3784: inst = 32'h10408000;
      3785: inst = 32'hc404719;
      3786: inst = 32'h8220000;
      3787: inst = 32'h10408000;
      3788: inst = 32'hc40471a;
      3789: inst = 32'h8220000;
      3790: inst = 32'h10408000;
      3791: inst = 32'hc40471b;
      3792: inst = 32'h8220000;
      3793: inst = 32'h10408000;
      3794: inst = 32'hc404744;
      3795: inst = 32'h8220000;
      3796: inst = 32'h10408000;
      3797: inst = 32'hc404745;
      3798: inst = 32'h8220000;
      3799: inst = 32'h10408000;
      3800: inst = 32'hc404746;
      3801: inst = 32'h8220000;
      3802: inst = 32'h10408000;
      3803: inst = 32'hc404747;
      3804: inst = 32'h8220000;
      3805: inst = 32'h10408000;
      3806: inst = 32'hc404748;
      3807: inst = 32'h8220000;
      3808: inst = 32'h10408000;
      3809: inst = 32'hc404749;
      3810: inst = 32'h8220000;
      3811: inst = 32'h10408000;
      3812: inst = 32'hc40474a;
      3813: inst = 32'h8220000;
      3814: inst = 32'h10408000;
      3815: inst = 32'hc40474b;
      3816: inst = 32'h8220000;
      3817: inst = 32'h10408000;
      3818: inst = 32'hc40474c;
      3819: inst = 32'h8220000;
      3820: inst = 32'h10408000;
      3821: inst = 32'hc40474d;
      3822: inst = 32'h8220000;
      3823: inst = 32'h10408000;
      3824: inst = 32'hc40474e;
      3825: inst = 32'h8220000;
      3826: inst = 32'h10408000;
      3827: inst = 32'hc404760;
      3828: inst = 32'h8220000;
      3829: inst = 32'h10408000;
      3830: inst = 32'hc404761;
      3831: inst = 32'h8220000;
      3832: inst = 32'h10408000;
      3833: inst = 32'hc404762;
      3834: inst = 32'h8220000;
      3835: inst = 32'h10408000;
      3836: inst = 32'hc404763;
      3837: inst = 32'h8220000;
      3838: inst = 32'h10408000;
      3839: inst = 32'hc404764;
      3840: inst = 32'h8220000;
      3841: inst = 32'h10408000;
      3842: inst = 32'hc404765;
      3843: inst = 32'h8220000;
      3844: inst = 32'h10408000;
      3845: inst = 32'hc404766;
      3846: inst = 32'h8220000;
      3847: inst = 32'h10408000;
      3848: inst = 32'hc404767;
      3849: inst = 32'h8220000;
      3850: inst = 32'h10408000;
      3851: inst = 32'hc404768;
      3852: inst = 32'h8220000;
      3853: inst = 32'h10408000;
      3854: inst = 32'hc404769;
      3855: inst = 32'h8220000;
      3856: inst = 32'h10408000;
      3857: inst = 32'hc40476a;
      3858: inst = 32'h8220000;
      3859: inst = 32'h10408000;
      3860: inst = 32'hc40476b;
      3861: inst = 32'h8220000;
      3862: inst = 32'h10408000;
      3863: inst = 32'hc40476c;
      3864: inst = 32'h8220000;
      3865: inst = 32'h10408000;
      3866: inst = 32'hc40476d;
      3867: inst = 32'h8220000;
      3868: inst = 32'h10408000;
      3869: inst = 32'hc40476e;
      3870: inst = 32'h8220000;
      3871: inst = 32'h10408000;
      3872: inst = 32'hc40476f;
      3873: inst = 32'h8220000;
      3874: inst = 32'h10408000;
      3875: inst = 32'hc404770;
      3876: inst = 32'h8220000;
      3877: inst = 32'h10408000;
      3878: inst = 32'hc404771;
      3879: inst = 32'h8220000;
      3880: inst = 32'h10408000;
      3881: inst = 32'hc404772;
      3882: inst = 32'h8220000;
      3883: inst = 32'h10408000;
      3884: inst = 32'hc404773;
      3885: inst = 32'h8220000;
      3886: inst = 32'h10408000;
      3887: inst = 32'hc404774;
      3888: inst = 32'h8220000;
      3889: inst = 32'h10408000;
      3890: inst = 32'hc404775;
      3891: inst = 32'h8220000;
      3892: inst = 32'h10408000;
      3893: inst = 32'hc404776;
      3894: inst = 32'h8220000;
      3895: inst = 32'h10408000;
      3896: inst = 32'hc404777;
      3897: inst = 32'h8220000;
      3898: inst = 32'h10408000;
      3899: inst = 32'hc404778;
      3900: inst = 32'h8220000;
      3901: inst = 32'h10408000;
      3902: inst = 32'hc404779;
      3903: inst = 32'h8220000;
      3904: inst = 32'h10408000;
      3905: inst = 32'hc40477a;
      3906: inst = 32'h8220000;
      3907: inst = 32'h10408000;
      3908: inst = 32'hc40477b;
      3909: inst = 32'h8220000;
      3910: inst = 32'h10408000;
      3911: inst = 32'hc4047a4;
      3912: inst = 32'h8220000;
      3913: inst = 32'h10408000;
      3914: inst = 32'hc4047a5;
      3915: inst = 32'h8220000;
      3916: inst = 32'h10408000;
      3917: inst = 32'hc4047a6;
      3918: inst = 32'h8220000;
      3919: inst = 32'h10408000;
      3920: inst = 32'hc4047a7;
      3921: inst = 32'h8220000;
      3922: inst = 32'h10408000;
      3923: inst = 32'hc4047a8;
      3924: inst = 32'h8220000;
      3925: inst = 32'h10408000;
      3926: inst = 32'hc4047a9;
      3927: inst = 32'h8220000;
      3928: inst = 32'h10408000;
      3929: inst = 32'hc4047aa;
      3930: inst = 32'h8220000;
      3931: inst = 32'h10408000;
      3932: inst = 32'hc4047ab;
      3933: inst = 32'h8220000;
      3934: inst = 32'h10408000;
      3935: inst = 32'hc4047ac;
      3936: inst = 32'h8220000;
      3937: inst = 32'h10408000;
      3938: inst = 32'hc4047ad;
      3939: inst = 32'h8220000;
      3940: inst = 32'h10408000;
      3941: inst = 32'hc4047ae;
      3942: inst = 32'h8220000;
      3943: inst = 32'h10408000;
      3944: inst = 32'hc4047c0;
      3945: inst = 32'h8220000;
      3946: inst = 32'h10408000;
      3947: inst = 32'hc4047c1;
      3948: inst = 32'h8220000;
      3949: inst = 32'h10408000;
      3950: inst = 32'hc4047c2;
      3951: inst = 32'h8220000;
      3952: inst = 32'h10408000;
      3953: inst = 32'hc4047c3;
      3954: inst = 32'h8220000;
      3955: inst = 32'h10408000;
      3956: inst = 32'hc4047c4;
      3957: inst = 32'h8220000;
      3958: inst = 32'h10408000;
      3959: inst = 32'hc4047c5;
      3960: inst = 32'h8220000;
      3961: inst = 32'h10408000;
      3962: inst = 32'hc4047c6;
      3963: inst = 32'h8220000;
      3964: inst = 32'h10408000;
      3965: inst = 32'hc4047c7;
      3966: inst = 32'h8220000;
      3967: inst = 32'h10408000;
      3968: inst = 32'hc4047c8;
      3969: inst = 32'h8220000;
      3970: inst = 32'h10408000;
      3971: inst = 32'hc4047c9;
      3972: inst = 32'h8220000;
      3973: inst = 32'h10408000;
      3974: inst = 32'hc4047ca;
      3975: inst = 32'h8220000;
      3976: inst = 32'h10408000;
      3977: inst = 32'hc4047cb;
      3978: inst = 32'h8220000;
      3979: inst = 32'h10408000;
      3980: inst = 32'hc4047cc;
      3981: inst = 32'h8220000;
      3982: inst = 32'h10408000;
      3983: inst = 32'hc4047cd;
      3984: inst = 32'h8220000;
      3985: inst = 32'h10408000;
      3986: inst = 32'hc4047ce;
      3987: inst = 32'h8220000;
      3988: inst = 32'h10408000;
      3989: inst = 32'hc4047cf;
      3990: inst = 32'h8220000;
      3991: inst = 32'h10408000;
      3992: inst = 32'hc4047d0;
      3993: inst = 32'h8220000;
      3994: inst = 32'h10408000;
      3995: inst = 32'hc4047d1;
      3996: inst = 32'h8220000;
      3997: inst = 32'h10408000;
      3998: inst = 32'hc4047d2;
      3999: inst = 32'h8220000;
      4000: inst = 32'h10408000;
      4001: inst = 32'hc4047d3;
      4002: inst = 32'h8220000;
      4003: inst = 32'h10408000;
      4004: inst = 32'hc4047d4;
      4005: inst = 32'h8220000;
      4006: inst = 32'h10408000;
      4007: inst = 32'hc4047d5;
      4008: inst = 32'h8220000;
      4009: inst = 32'h10408000;
      4010: inst = 32'hc4047d6;
      4011: inst = 32'h8220000;
      4012: inst = 32'h10408000;
      4013: inst = 32'hc4047d7;
      4014: inst = 32'h8220000;
      4015: inst = 32'h10408000;
      4016: inst = 32'hc4047d8;
      4017: inst = 32'h8220000;
      4018: inst = 32'h10408000;
      4019: inst = 32'hc4047d9;
      4020: inst = 32'h8220000;
      4021: inst = 32'h10408000;
      4022: inst = 32'hc4047da;
      4023: inst = 32'h8220000;
      4024: inst = 32'h10408000;
      4025: inst = 32'hc4047db;
      4026: inst = 32'h8220000;
      4027: inst = 32'h10408000;
      4028: inst = 32'hc404804;
      4029: inst = 32'h8220000;
      4030: inst = 32'h10408000;
      4031: inst = 32'hc404805;
      4032: inst = 32'h8220000;
      4033: inst = 32'h10408000;
      4034: inst = 32'hc404806;
      4035: inst = 32'h8220000;
      4036: inst = 32'h10408000;
      4037: inst = 32'hc404807;
      4038: inst = 32'h8220000;
      4039: inst = 32'h10408000;
      4040: inst = 32'hc404808;
      4041: inst = 32'h8220000;
      4042: inst = 32'h10408000;
      4043: inst = 32'hc404809;
      4044: inst = 32'h8220000;
      4045: inst = 32'h10408000;
      4046: inst = 32'hc40480a;
      4047: inst = 32'h8220000;
      4048: inst = 32'h10408000;
      4049: inst = 32'hc40480b;
      4050: inst = 32'h8220000;
      4051: inst = 32'h10408000;
      4052: inst = 32'hc40480c;
      4053: inst = 32'h8220000;
      4054: inst = 32'h10408000;
      4055: inst = 32'hc40480d;
      4056: inst = 32'h8220000;
      4057: inst = 32'h10408000;
      4058: inst = 32'hc40480e;
      4059: inst = 32'h8220000;
      4060: inst = 32'h10408000;
      4061: inst = 32'hc404820;
      4062: inst = 32'h8220000;
      4063: inst = 32'h10408000;
      4064: inst = 32'hc404821;
      4065: inst = 32'h8220000;
      4066: inst = 32'h10408000;
      4067: inst = 32'hc404822;
      4068: inst = 32'h8220000;
      4069: inst = 32'h10408000;
      4070: inst = 32'hc404823;
      4071: inst = 32'h8220000;
      4072: inst = 32'h10408000;
      4073: inst = 32'hc404824;
      4074: inst = 32'h8220000;
      4075: inst = 32'h10408000;
      4076: inst = 32'hc404825;
      4077: inst = 32'h8220000;
      4078: inst = 32'h10408000;
      4079: inst = 32'hc404826;
      4080: inst = 32'h8220000;
      4081: inst = 32'h10408000;
      4082: inst = 32'hc404827;
      4083: inst = 32'h8220000;
      4084: inst = 32'h10408000;
      4085: inst = 32'hc404828;
      4086: inst = 32'h8220000;
      4087: inst = 32'h10408000;
      4088: inst = 32'hc404829;
      4089: inst = 32'h8220000;
      4090: inst = 32'h10408000;
      4091: inst = 32'hc40482a;
      4092: inst = 32'h8220000;
      4093: inst = 32'h10408000;
      4094: inst = 32'hc40482b;
      4095: inst = 32'h8220000;
      4096: inst = 32'h10408000;
      4097: inst = 32'hc40482c;
      4098: inst = 32'h8220000;
      4099: inst = 32'h10408000;
      4100: inst = 32'hc40482d;
      4101: inst = 32'h8220000;
      4102: inst = 32'h10408000;
      4103: inst = 32'hc40482e;
      4104: inst = 32'h8220000;
      4105: inst = 32'h10408000;
      4106: inst = 32'hc40482f;
      4107: inst = 32'h8220000;
      4108: inst = 32'h10408000;
      4109: inst = 32'hc404830;
      4110: inst = 32'h8220000;
      4111: inst = 32'h10408000;
      4112: inst = 32'hc404831;
      4113: inst = 32'h8220000;
      4114: inst = 32'h10408000;
      4115: inst = 32'hc404832;
      4116: inst = 32'h8220000;
      4117: inst = 32'h10408000;
      4118: inst = 32'hc404833;
      4119: inst = 32'h8220000;
      4120: inst = 32'h10408000;
      4121: inst = 32'hc404834;
      4122: inst = 32'h8220000;
      4123: inst = 32'h10408000;
      4124: inst = 32'hc404835;
      4125: inst = 32'h8220000;
      4126: inst = 32'h10408000;
      4127: inst = 32'hc404836;
      4128: inst = 32'h8220000;
      4129: inst = 32'h10408000;
      4130: inst = 32'hc404837;
      4131: inst = 32'h8220000;
      4132: inst = 32'h10408000;
      4133: inst = 32'hc404838;
      4134: inst = 32'h8220000;
      4135: inst = 32'h10408000;
      4136: inst = 32'hc404839;
      4137: inst = 32'h8220000;
      4138: inst = 32'h10408000;
      4139: inst = 32'hc40483a;
      4140: inst = 32'h8220000;
      4141: inst = 32'h10408000;
      4142: inst = 32'hc40483b;
      4143: inst = 32'h8220000;
      4144: inst = 32'h10408000;
      4145: inst = 32'hc404864;
      4146: inst = 32'h8220000;
      4147: inst = 32'h10408000;
      4148: inst = 32'hc404865;
      4149: inst = 32'h8220000;
      4150: inst = 32'h10408000;
      4151: inst = 32'hc404866;
      4152: inst = 32'h8220000;
      4153: inst = 32'h10408000;
      4154: inst = 32'hc404867;
      4155: inst = 32'h8220000;
      4156: inst = 32'h10408000;
      4157: inst = 32'hc404868;
      4158: inst = 32'h8220000;
      4159: inst = 32'h10408000;
      4160: inst = 32'hc404869;
      4161: inst = 32'h8220000;
      4162: inst = 32'h10408000;
      4163: inst = 32'hc40486a;
      4164: inst = 32'h8220000;
      4165: inst = 32'h10408000;
      4166: inst = 32'hc40486b;
      4167: inst = 32'h8220000;
      4168: inst = 32'h10408000;
      4169: inst = 32'hc40486c;
      4170: inst = 32'h8220000;
      4171: inst = 32'h10408000;
      4172: inst = 32'hc40486d;
      4173: inst = 32'h8220000;
      4174: inst = 32'h10408000;
      4175: inst = 32'hc40486e;
      4176: inst = 32'h8220000;
      4177: inst = 32'h10408000;
      4178: inst = 32'hc404880;
      4179: inst = 32'h8220000;
      4180: inst = 32'h10408000;
      4181: inst = 32'hc404881;
      4182: inst = 32'h8220000;
      4183: inst = 32'h10408000;
      4184: inst = 32'hc404882;
      4185: inst = 32'h8220000;
      4186: inst = 32'h10408000;
      4187: inst = 32'hc404883;
      4188: inst = 32'h8220000;
      4189: inst = 32'h10408000;
      4190: inst = 32'hc404884;
      4191: inst = 32'h8220000;
      4192: inst = 32'h10408000;
      4193: inst = 32'hc404885;
      4194: inst = 32'h8220000;
      4195: inst = 32'h10408000;
      4196: inst = 32'hc404886;
      4197: inst = 32'h8220000;
      4198: inst = 32'h10408000;
      4199: inst = 32'hc404887;
      4200: inst = 32'h8220000;
      4201: inst = 32'h10408000;
      4202: inst = 32'hc404888;
      4203: inst = 32'h8220000;
      4204: inst = 32'h10408000;
      4205: inst = 32'hc404889;
      4206: inst = 32'h8220000;
      4207: inst = 32'h10408000;
      4208: inst = 32'hc40488a;
      4209: inst = 32'h8220000;
      4210: inst = 32'h10408000;
      4211: inst = 32'hc40488b;
      4212: inst = 32'h8220000;
      4213: inst = 32'h10408000;
      4214: inst = 32'hc40488c;
      4215: inst = 32'h8220000;
      4216: inst = 32'h10408000;
      4217: inst = 32'hc40488d;
      4218: inst = 32'h8220000;
      4219: inst = 32'h10408000;
      4220: inst = 32'hc40488e;
      4221: inst = 32'h8220000;
      4222: inst = 32'h10408000;
      4223: inst = 32'hc40488f;
      4224: inst = 32'h8220000;
      4225: inst = 32'h10408000;
      4226: inst = 32'hc404890;
      4227: inst = 32'h8220000;
      4228: inst = 32'h10408000;
      4229: inst = 32'hc404891;
      4230: inst = 32'h8220000;
      4231: inst = 32'h10408000;
      4232: inst = 32'hc404892;
      4233: inst = 32'h8220000;
      4234: inst = 32'h10408000;
      4235: inst = 32'hc404893;
      4236: inst = 32'h8220000;
      4237: inst = 32'h10408000;
      4238: inst = 32'hc404894;
      4239: inst = 32'h8220000;
      4240: inst = 32'h10408000;
      4241: inst = 32'hc404895;
      4242: inst = 32'h8220000;
      4243: inst = 32'h10408000;
      4244: inst = 32'hc404896;
      4245: inst = 32'h8220000;
      4246: inst = 32'h10408000;
      4247: inst = 32'hc404897;
      4248: inst = 32'h8220000;
      4249: inst = 32'h10408000;
      4250: inst = 32'hc404898;
      4251: inst = 32'h8220000;
      4252: inst = 32'h10408000;
      4253: inst = 32'hc404899;
      4254: inst = 32'h8220000;
      4255: inst = 32'h10408000;
      4256: inst = 32'hc40489a;
      4257: inst = 32'h8220000;
      4258: inst = 32'h10408000;
      4259: inst = 32'hc40489b;
      4260: inst = 32'h8220000;
      4261: inst = 32'h10408000;
      4262: inst = 32'hc4048c4;
      4263: inst = 32'h8220000;
      4264: inst = 32'h10408000;
      4265: inst = 32'hc4048c5;
      4266: inst = 32'h8220000;
      4267: inst = 32'h10408000;
      4268: inst = 32'hc4048c6;
      4269: inst = 32'h8220000;
      4270: inst = 32'h10408000;
      4271: inst = 32'hc4048c7;
      4272: inst = 32'h8220000;
      4273: inst = 32'h10408000;
      4274: inst = 32'hc4048c8;
      4275: inst = 32'h8220000;
      4276: inst = 32'h10408000;
      4277: inst = 32'hc4048c9;
      4278: inst = 32'h8220000;
      4279: inst = 32'h10408000;
      4280: inst = 32'hc4048ca;
      4281: inst = 32'h8220000;
      4282: inst = 32'h10408000;
      4283: inst = 32'hc4048cb;
      4284: inst = 32'h8220000;
      4285: inst = 32'h10408000;
      4286: inst = 32'hc4048cc;
      4287: inst = 32'h8220000;
      4288: inst = 32'h10408000;
      4289: inst = 32'hc4048cd;
      4290: inst = 32'h8220000;
      4291: inst = 32'h10408000;
      4292: inst = 32'hc4048ce;
      4293: inst = 32'h8220000;
      4294: inst = 32'h10408000;
      4295: inst = 32'hc4048e0;
      4296: inst = 32'h8220000;
      4297: inst = 32'h10408000;
      4298: inst = 32'hc4048e1;
      4299: inst = 32'h8220000;
      4300: inst = 32'h10408000;
      4301: inst = 32'hc4048e2;
      4302: inst = 32'h8220000;
      4303: inst = 32'h10408000;
      4304: inst = 32'hc4048e3;
      4305: inst = 32'h8220000;
      4306: inst = 32'h10408000;
      4307: inst = 32'hc4048e4;
      4308: inst = 32'h8220000;
      4309: inst = 32'h10408000;
      4310: inst = 32'hc4048e5;
      4311: inst = 32'h8220000;
      4312: inst = 32'h10408000;
      4313: inst = 32'hc4048e6;
      4314: inst = 32'h8220000;
      4315: inst = 32'h10408000;
      4316: inst = 32'hc4048e7;
      4317: inst = 32'h8220000;
      4318: inst = 32'h10408000;
      4319: inst = 32'hc4048e8;
      4320: inst = 32'h8220000;
      4321: inst = 32'h10408000;
      4322: inst = 32'hc4048e9;
      4323: inst = 32'h8220000;
      4324: inst = 32'h10408000;
      4325: inst = 32'hc4048ea;
      4326: inst = 32'h8220000;
      4327: inst = 32'h10408000;
      4328: inst = 32'hc4048eb;
      4329: inst = 32'h8220000;
      4330: inst = 32'h10408000;
      4331: inst = 32'hc4048ec;
      4332: inst = 32'h8220000;
      4333: inst = 32'h10408000;
      4334: inst = 32'hc4048ed;
      4335: inst = 32'h8220000;
      4336: inst = 32'h10408000;
      4337: inst = 32'hc4048ee;
      4338: inst = 32'h8220000;
      4339: inst = 32'h10408000;
      4340: inst = 32'hc4048ef;
      4341: inst = 32'h8220000;
      4342: inst = 32'h10408000;
      4343: inst = 32'hc4048f0;
      4344: inst = 32'h8220000;
      4345: inst = 32'h10408000;
      4346: inst = 32'hc4048f1;
      4347: inst = 32'h8220000;
      4348: inst = 32'h10408000;
      4349: inst = 32'hc4048f2;
      4350: inst = 32'h8220000;
      4351: inst = 32'h10408000;
      4352: inst = 32'hc4048f3;
      4353: inst = 32'h8220000;
      4354: inst = 32'h10408000;
      4355: inst = 32'hc4048f4;
      4356: inst = 32'h8220000;
      4357: inst = 32'h10408000;
      4358: inst = 32'hc4048f5;
      4359: inst = 32'h8220000;
      4360: inst = 32'h10408000;
      4361: inst = 32'hc4048f6;
      4362: inst = 32'h8220000;
      4363: inst = 32'h10408000;
      4364: inst = 32'hc4048f7;
      4365: inst = 32'h8220000;
      4366: inst = 32'h10408000;
      4367: inst = 32'hc4048f8;
      4368: inst = 32'h8220000;
      4369: inst = 32'h10408000;
      4370: inst = 32'hc4048f9;
      4371: inst = 32'h8220000;
      4372: inst = 32'h10408000;
      4373: inst = 32'hc4048fa;
      4374: inst = 32'h8220000;
      4375: inst = 32'h10408000;
      4376: inst = 32'hc4048fb;
      4377: inst = 32'h8220000;
      4378: inst = 32'h10408000;
      4379: inst = 32'hc404924;
      4380: inst = 32'h8220000;
      4381: inst = 32'h10408000;
      4382: inst = 32'hc404925;
      4383: inst = 32'h8220000;
      4384: inst = 32'h10408000;
      4385: inst = 32'hc404926;
      4386: inst = 32'h8220000;
      4387: inst = 32'h10408000;
      4388: inst = 32'hc404927;
      4389: inst = 32'h8220000;
      4390: inst = 32'h10408000;
      4391: inst = 32'hc404928;
      4392: inst = 32'h8220000;
      4393: inst = 32'h10408000;
      4394: inst = 32'hc404929;
      4395: inst = 32'h8220000;
      4396: inst = 32'h10408000;
      4397: inst = 32'hc40492a;
      4398: inst = 32'h8220000;
      4399: inst = 32'h10408000;
      4400: inst = 32'hc40492b;
      4401: inst = 32'h8220000;
      4402: inst = 32'h10408000;
      4403: inst = 32'hc40492c;
      4404: inst = 32'h8220000;
      4405: inst = 32'h10408000;
      4406: inst = 32'hc40492d;
      4407: inst = 32'h8220000;
      4408: inst = 32'h10408000;
      4409: inst = 32'hc40492e;
      4410: inst = 32'h8220000;
      4411: inst = 32'h10408000;
      4412: inst = 32'hc404940;
      4413: inst = 32'h8220000;
      4414: inst = 32'h10408000;
      4415: inst = 32'hc404941;
      4416: inst = 32'h8220000;
      4417: inst = 32'h10408000;
      4418: inst = 32'hc404942;
      4419: inst = 32'h8220000;
      4420: inst = 32'h10408000;
      4421: inst = 32'hc404943;
      4422: inst = 32'h8220000;
      4423: inst = 32'h10408000;
      4424: inst = 32'hc404944;
      4425: inst = 32'h8220000;
      4426: inst = 32'h10408000;
      4427: inst = 32'hc404945;
      4428: inst = 32'h8220000;
      4429: inst = 32'h10408000;
      4430: inst = 32'hc404946;
      4431: inst = 32'h8220000;
      4432: inst = 32'h10408000;
      4433: inst = 32'hc404947;
      4434: inst = 32'h8220000;
      4435: inst = 32'h10408000;
      4436: inst = 32'hc404948;
      4437: inst = 32'h8220000;
      4438: inst = 32'h10408000;
      4439: inst = 32'hc404949;
      4440: inst = 32'h8220000;
      4441: inst = 32'h10408000;
      4442: inst = 32'hc40494a;
      4443: inst = 32'h8220000;
      4444: inst = 32'h10408000;
      4445: inst = 32'hc40494b;
      4446: inst = 32'h8220000;
      4447: inst = 32'h10408000;
      4448: inst = 32'hc40494c;
      4449: inst = 32'h8220000;
      4450: inst = 32'h10408000;
      4451: inst = 32'hc40494d;
      4452: inst = 32'h8220000;
      4453: inst = 32'h10408000;
      4454: inst = 32'hc40494e;
      4455: inst = 32'h8220000;
      4456: inst = 32'h10408000;
      4457: inst = 32'hc40494f;
      4458: inst = 32'h8220000;
      4459: inst = 32'h10408000;
      4460: inst = 32'hc404950;
      4461: inst = 32'h8220000;
      4462: inst = 32'h10408000;
      4463: inst = 32'hc404951;
      4464: inst = 32'h8220000;
      4465: inst = 32'h10408000;
      4466: inst = 32'hc404952;
      4467: inst = 32'h8220000;
      4468: inst = 32'h10408000;
      4469: inst = 32'hc404953;
      4470: inst = 32'h8220000;
      4471: inst = 32'h10408000;
      4472: inst = 32'hc404954;
      4473: inst = 32'h8220000;
      4474: inst = 32'h10408000;
      4475: inst = 32'hc404955;
      4476: inst = 32'h8220000;
      4477: inst = 32'h10408000;
      4478: inst = 32'hc404956;
      4479: inst = 32'h8220000;
      4480: inst = 32'h10408000;
      4481: inst = 32'hc404957;
      4482: inst = 32'h8220000;
      4483: inst = 32'h10408000;
      4484: inst = 32'hc404958;
      4485: inst = 32'h8220000;
      4486: inst = 32'h10408000;
      4487: inst = 32'hc404959;
      4488: inst = 32'h8220000;
      4489: inst = 32'h10408000;
      4490: inst = 32'hc40495a;
      4491: inst = 32'h8220000;
      4492: inst = 32'h10408000;
      4493: inst = 32'hc40495b;
      4494: inst = 32'h8220000;
      4495: inst = 32'h10408000;
      4496: inst = 32'hc404984;
      4497: inst = 32'h8220000;
      4498: inst = 32'h10408000;
      4499: inst = 32'hc404985;
      4500: inst = 32'h8220000;
      4501: inst = 32'h10408000;
      4502: inst = 32'hc404986;
      4503: inst = 32'h8220000;
      4504: inst = 32'h10408000;
      4505: inst = 32'hc404987;
      4506: inst = 32'h8220000;
      4507: inst = 32'h10408000;
      4508: inst = 32'hc404988;
      4509: inst = 32'h8220000;
      4510: inst = 32'h10408000;
      4511: inst = 32'hc404989;
      4512: inst = 32'h8220000;
      4513: inst = 32'h10408000;
      4514: inst = 32'hc40498a;
      4515: inst = 32'h8220000;
      4516: inst = 32'h10408000;
      4517: inst = 32'hc40498b;
      4518: inst = 32'h8220000;
      4519: inst = 32'h10408000;
      4520: inst = 32'hc40498c;
      4521: inst = 32'h8220000;
      4522: inst = 32'h10408000;
      4523: inst = 32'hc40498d;
      4524: inst = 32'h8220000;
      4525: inst = 32'h10408000;
      4526: inst = 32'hc40498e;
      4527: inst = 32'h8220000;
      4528: inst = 32'h10408000;
      4529: inst = 32'hc4049a0;
      4530: inst = 32'h8220000;
      4531: inst = 32'h10408000;
      4532: inst = 32'hc4049a1;
      4533: inst = 32'h8220000;
      4534: inst = 32'h10408000;
      4535: inst = 32'hc4049a2;
      4536: inst = 32'h8220000;
      4537: inst = 32'h10408000;
      4538: inst = 32'hc4049a3;
      4539: inst = 32'h8220000;
      4540: inst = 32'h10408000;
      4541: inst = 32'hc4049a4;
      4542: inst = 32'h8220000;
      4543: inst = 32'h10408000;
      4544: inst = 32'hc4049a5;
      4545: inst = 32'h8220000;
      4546: inst = 32'h10408000;
      4547: inst = 32'hc4049a6;
      4548: inst = 32'h8220000;
      4549: inst = 32'h10408000;
      4550: inst = 32'hc4049a7;
      4551: inst = 32'h8220000;
      4552: inst = 32'h10408000;
      4553: inst = 32'hc4049a8;
      4554: inst = 32'h8220000;
      4555: inst = 32'h10408000;
      4556: inst = 32'hc4049a9;
      4557: inst = 32'h8220000;
      4558: inst = 32'h10408000;
      4559: inst = 32'hc4049aa;
      4560: inst = 32'h8220000;
      4561: inst = 32'h10408000;
      4562: inst = 32'hc4049ab;
      4563: inst = 32'h8220000;
      4564: inst = 32'h10408000;
      4565: inst = 32'hc4049ac;
      4566: inst = 32'h8220000;
      4567: inst = 32'h10408000;
      4568: inst = 32'hc4049ad;
      4569: inst = 32'h8220000;
      4570: inst = 32'h10408000;
      4571: inst = 32'hc4049ae;
      4572: inst = 32'h8220000;
      4573: inst = 32'h10408000;
      4574: inst = 32'hc4049af;
      4575: inst = 32'h8220000;
      4576: inst = 32'h10408000;
      4577: inst = 32'hc4049b0;
      4578: inst = 32'h8220000;
      4579: inst = 32'h10408000;
      4580: inst = 32'hc4049b1;
      4581: inst = 32'h8220000;
      4582: inst = 32'h10408000;
      4583: inst = 32'hc4049b2;
      4584: inst = 32'h8220000;
      4585: inst = 32'h10408000;
      4586: inst = 32'hc4049b3;
      4587: inst = 32'h8220000;
      4588: inst = 32'h10408000;
      4589: inst = 32'hc4049b4;
      4590: inst = 32'h8220000;
      4591: inst = 32'h10408000;
      4592: inst = 32'hc4049b5;
      4593: inst = 32'h8220000;
      4594: inst = 32'h10408000;
      4595: inst = 32'hc4049b6;
      4596: inst = 32'h8220000;
      4597: inst = 32'h10408000;
      4598: inst = 32'hc4049b7;
      4599: inst = 32'h8220000;
      4600: inst = 32'h10408000;
      4601: inst = 32'hc4049b8;
      4602: inst = 32'h8220000;
      4603: inst = 32'h10408000;
      4604: inst = 32'hc4049b9;
      4605: inst = 32'h8220000;
      4606: inst = 32'h10408000;
      4607: inst = 32'hc4049ba;
      4608: inst = 32'h8220000;
      4609: inst = 32'h10408000;
      4610: inst = 32'hc4049bb;
      4611: inst = 32'h8220000;
      4612: inst = 32'h10408000;
      4613: inst = 32'hc4049e4;
      4614: inst = 32'h8220000;
      4615: inst = 32'h10408000;
      4616: inst = 32'hc4049e5;
      4617: inst = 32'h8220000;
      4618: inst = 32'h10408000;
      4619: inst = 32'hc4049e6;
      4620: inst = 32'h8220000;
      4621: inst = 32'h10408000;
      4622: inst = 32'hc4049e7;
      4623: inst = 32'h8220000;
      4624: inst = 32'h10408000;
      4625: inst = 32'hc4049e8;
      4626: inst = 32'h8220000;
      4627: inst = 32'h10408000;
      4628: inst = 32'hc4049e9;
      4629: inst = 32'h8220000;
      4630: inst = 32'h10408000;
      4631: inst = 32'hc4049ea;
      4632: inst = 32'h8220000;
      4633: inst = 32'h10408000;
      4634: inst = 32'hc4049eb;
      4635: inst = 32'h8220000;
      4636: inst = 32'h10408000;
      4637: inst = 32'hc4049ec;
      4638: inst = 32'h8220000;
      4639: inst = 32'h10408000;
      4640: inst = 32'hc4049ed;
      4641: inst = 32'h8220000;
      4642: inst = 32'h10408000;
      4643: inst = 32'hc4049ee;
      4644: inst = 32'h8220000;
      4645: inst = 32'h10408000;
      4646: inst = 32'hc404a00;
      4647: inst = 32'h8220000;
      4648: inst = 32'h10408000;
      4649: inst = 32'hc404a01;
      4650: inst = 32'h8220000;
      4651: inst = 32'h10408000;
      4652: inst = 32'hc404a02;
      4653: inst = 32'h8220000;
      4654: inst = 32'h10408000;
      4655: inst = 32'hc404a03;
      4656: inst = 32'h8220000;
      4657: inst = 32'h10408000;
      4658: inst = 32'hc404a04;
      4659: inst = 32'h8220000;
      4660: inst = 32'h10408000;
      4661: inst = 32'hc404a05;
      4662: inst = 32'h8220000;
      4663: inst = 32'h10408000;
      4664: inst = 32'hc404a06;
      4665: inst = 32'h8220000;
      4666: inst = 32'h10408000;
      4667: inst = 32'hc404a07;
      4668: inst = 32'h8220000;
      4669: inst = 32'h10408000;
      4670: inst = 32'hc404a0f;
      4671: inst = 32'h8220000;
      4672: inst = 32'h10408000;
      4673: inst = 32'hc404a10;
      4674: inst = 32'h8220000;
      4675: inst = 32'h10408000;
      4676: inst = 32'hc404a11;
      4677: inst = 32'h8220000;
      4678: inst = 32'h10408000;
      4679: inst = 32'hc404a12;
      4680: inst = 32'h8220000;
      4681: inst = 32'h10408000;
      4682: inst = 32'hc404a13;
      4683: inst = 32'h8220000;
      4684: inst = 32'h10408000;
      4685: inst = 32'hc404a14;
      4686: inst = 32'h8220000;
      4687: inst = 32'h10408000;
      4688: inst = 32'hc404a15;
      4689: inst = 32'h8220000;
      4690: inst = 32'h10408000;
      4691: inst = 32'hc404a16;
      4692: inst = 32'h8220000;
      4693: inst = 32'h10408000;
      4694: inst = 32'hc404a17;
      4695: inst = 32'h8220000;
      4696: inst = 32'h10408000;
      4697: inst = 32'hc404a18;
      4698: inst = 32'h8220000;
      4699: inst = 32'h10408000;
      4700: inst = 32'hc404a19;
      4701: inst = 32'h8220000;
      4702: inst = 32'h10408000;
      4703: inst = 32'hc404a1a;
      4704: inst = 32'h8220000;
      4705: inst = 32'h10408000;
      4706: inst = 32'hc404a1b;
      4707: inst = 32'h8220000;
      4708: inst = 32'h10408000;
      4709: inst = 32'hc404a44;
      4710: inst = 32'h8220000;
      4711: inst = 32'h10408000;
      4712: inst = 32'hc404a45;
      4713: inst = 32'h8220000;
      4714: inst = 32'h10408000;
      4715: inst = 32'hc404a46;
      4716: inst = 32'h8220000;
      4717: inst = 32'h10408000;
      4718: inst = 32'hc404a47;
      4719: inst = 32'h8220000;
      4720: inst = 32'h10408000;
      4721: inst = 32'hc404a48;
      4722: inst = 32'h8220000;
      4723: inst = 32'h10408000;
      4724: inst = 32'hc404a49;
      4725: inst = 32'h8220000;
      4726: inst = 32'h10408000;
      4727: inst = 32'hc404a4a;
      4728: inst = 32'h8220000;
      4729: inst = 32'h10408000;
      4730: inst = 32'hc404a4b;
      4731: inst = 32'h8220000;
      4732: inst = 32'h10408000;
      4733: inst = 32'hc404a4c;
      4734: inst = 32'h8220000;
      4735: inst = 32'h10408000;
      4736: inst = 32'hc404a4d;
      4737: inst = 32'h8220000;
      4738: inst = 32'h10408000;
      4739: inst = 32'hc404a4e;
      4740: inst = 32'h8220000;
      4741: inst = 32'h10408000;
      4742: inst = 32'hc404a60;
      4743: inst = 32'h8220000;
      4744: inst = 32'h10408000;
      4745: inst = 32'hc404a61;
      4746: inst = 32'h8220000;
      4747: inst = 32'h10408000;
      4748: inst = 32'hc404a62;
      4749: inst = 32'h8220000;
      4750: inst = 32'h10408000;
      4751: inst = 32'hc404a63;
      4752: inst = 32'h8220000;
      4753: inst = 32'h10408000;
      4754: inst = 32'hc404a64;
      4755: inst = 32'h8220000;
      4756: inst = 32'h10408000;
      4757: inst = 32'hc404a65;
      4758: inst = 32'h8220000;
      4759: inst = 32'h10408000;
      4760: inst = 32'hc404a66;
      4761: inst = 32'h8220000;
      4762: inst = 32'h10408000;
      4763: inst = 32'hc404a70;
      4764: inst = 32'h8220000;
      4765: inst = 32'h10408000;
      4766: inst = 32'hc404a71;
      4767: inst = 32'h8220000;
      4768: inst = 32'h10408000;
      4769: inst = 32'hc404a72;
      4770: inst = 32'h8220000;
      4771: inst = 32'h10408000;
      4772: inst = 32'hc404a73;
      4773: inst = 32'h8220000;
      4774: inst = 32'h10408000;
      4775: inst = 32'hc404a74;
      4776: inst = 32'h8220000;
      4777: inst = 32'h10408000;
      4778: inst = 32'hc404a75;
      4779: inst = 32'h8220000;
      4780: inst = 32'h10408000;
      4781: inst = 32'hc404a76;
      4782: inst = 32'h8220000;
      4783: inst = 32'h10408000;
      4784: inst = 32'hc404a77;
      4785: inst = 32'h8220000;
      4786: inst = 32'h10408000;
      4787: inst = 32'hc404a78;
      4788: inst = 32'h8220000;
      4789: inst = 32'h10408000;
      4790: inst = 32'hc404a79;
      4791: inst = 32'h8220000;
      4792: inst = 32'h10408000;
      4793: inst = 32'hc404a7a;
      4794: inst = 32'h8220000;
      4795: inst = 32'h10408000;
      4796: inst = 32'hc404a7b;
      4797: inst = 32'h8220000;
      4798: inst = 32'h10408000;
      4799: inst = 32'hc404aa4;
      4800: inst = 32'h8220000;
      4801: inst = 32'h10408000;
      4802: inst = 32'hc404aa5;
      4803: inst = 32'h8220000;
      4804: inst = 32'h10408000;
      4805: inst = 32'hc404aa6;
      4806: inst = 32'h8220000;
      4807: inst = 32'h10408000;
      4808: inst = 32'hc404aa7;
      4809: inst = 32'h8220000;
      4810: inst = 32'h10408000;
      4811: inst = 32'hc404aa8;
      4812: inst = 32'h8220000;
      4813: inst = 32'h10408000;
      4814: inst = 32'hc404aa9;
      4815: inst = 32'h8220000;
      4816: inst = 32'h10408000;
      4817: inst = 32'hc404aaa;
      4818: inst = 32'h8220000;
      4819: inst = 32'h10408000;
      4820: inst = 32'hc404aab;
      4821: inst = 32'h8220000;
      4822: inst = 32'h10408000;
      4823: inst = 32'hc404aac;
      4824: inst = 32'h8220000;
      4825: inst = 32'h10408000;
      4826: inst = 32'hc404aad;
      4827: inst = 32'h8220000;
      4828: inst = 32'h10408000;
      4829: inst = 32'hc404aae;
      4830: inst = 32'h8220000;
      4831: inst = 32'h10408000;
      4832: inst = 32'hc404ac0;
      4833: inst = 32'h8220000;
      4834: inst = 32'h10408000;
      4835: inst = 32'hc404ac1;
      4836: inst = 32'h8220000;
      4837: inst = 32'h10408000;
      4838: inst = 32'hc404ac2;
      4839: inst = 32'h8220000;
      4840: inst = 32'h10408000;
      4841: inst = 32'hc404ac3;
      4842: inst = 32'h8220000;
      4843: inst = 32'h10408000;
      4844: inst = 32'hc404ac4;
      4845: inst = 32'h8220000;
      4846: inst = 32'h10408000;
      4847: inst = 32'hc404ac5;
      4848: inst = 32'h8220000;
      4849: inst = 32'h10408000;
      4850: inst = 32'hc404ac6;
      4851: inst = 32'h8220000;
      4852: inst = 32'h10408000;
      4853: inst = 32'hc404ad0;
      4854: inst = 32'h8220000;
      4855: inst = 32'h10408000;
      4856: inst = 32'hc404ad1;
      4857: inst = 32'h8220000;
      4858: inst = 32'h10408000;
      4859: inst = 32'hc404ad2;
      4860: inst = 32'h8220000;
      4861: inst = 32'h10408000;
      4862: inst = 32'hc404ad3;
      4863: inst = 32'h8220000;
      4864: inst = 32'h10408000;
      4865: inst = 32'hc404ad4;
      4866: inst = 32'h8220000;
      4867: inst = 32'h10408000;
      4868: inst = 32'hc404ad5;
      4869: inst = 32'h8220000;
      4870: inst = 32'h10408000;
      4871: inst = 32'hc404ad6;
      4872: inst = 32'h8220000;
      4873: inst = 32'h10408000;
      4874: inst = 32'hc404ad7;
      4875: inst = 32'h8220000;
      4876: inst = 32'h10408000;
      4877: inst = 32'hc404ad8;
      4878: inst = 32'h8220000;
      4879: inst = 32'h10408000;
      4880: inst = 32'hc404ad9;
      4881: inst = 32'h8220000;
      4882: inst = 32'h10408000;
      4883: inst = 32'hc404ada;
      4884: inst = 32'h8220000;
      4885: inst = 32'h10408000;
      4886: inst = 32'hc404adb;
      4887: inst = 32'h8220000;
      4888: inst = 32'h10408000;
      4889: inst = 32'hc404b04;
      4890: inst = 32'h8220000;
      4891: inst = 32'h10408000;
      4892: inst = 32'hc404b05;
      4893: inst = 32'h8220000;
      4894: inst = 32'h10408000;
      4895: inst = 32'hc404b06;
      4896: inst = 32'h8220000;
      4897: inst = 32'h10408000;
      4898: inst = 32'hc404b07;
      4899: inst = 32'h8220000;
      4900: inst = 32'h10408000;
      4901: inst = 32'hc404b08;
      4902: inst = 32'h8220000;
      4903: inst = 32'h10408000;
      4904: inst = 32'hc404b09;
      4905: inst = 32'h8220000;
      4906: inst = 32'h10408000;
      4907: inst = 32'hc404b0a;
      4908: inst = 32'h8220000;
      4909: inst = 32'h10408000;
      4910: inst = 32'hc404b0b;
      4911: inst = 32'h8220000;
      4912: inst = 32'h10408000;
      4913: inst = 32'hc404b0c;
      4914: inst = 32'h8220000;
      4915: inst = 32'h10408000;
      4916: inst = 32'hc404b0d;
      4917: inst = 32'h8220000;
      4918: inst = 32'h10408000;
      4919: inst = 32'hc404b0e;
      4920: inst = 32'h8220000;
      4921: inst = 32'h10408000;
      4922: inst = 32'hc404b20;
      4923: inst = 32'h8220000;
      4924: inst = 32'h10408000;
      4925: inst = 32'hc404b21;
      4926: inst = 32'h8220000;
      4927: inst = 32'h10408000;
      4928: inst = 32'hc404b22;
      4929: inst = 32'h8220000;
      4930: inst = 32'h10408000;
      4931: inst = 32'hc404b23;
      4932: inst = 32'h8220000;
      4933: inst = 32'h10408000;
      4934: inst = 32'hc404b24;
      4935: inst = 32'h8220000;
      4936: inst = 32'h10408000;
      4937: inst = 32'hc404b25;
      4938: inst = 32'h8220000;
      4939: inst = 32'h10408000;
      4940: inst = 32'hc404b26;
      4941: inst = 32'h8220000;
      4942: inst = 32'h10408000;
      4943: inst = 32'hc404b30;
      4944: inst = 32'h8220000;
      4945: inst = 32'h10408000;
      4946: inst = 32'hc404b31;
      4947: inst = 32'h8220000;
      4948: inst = 32'h10408000;
      4949: inst = 32'hc404b32;
      4950: inst = 32'h8220000;
      4951: inst = 32'h10408000;
      4952: inst = 32'hc404b33;
      4953: inst = 32'h8220000;
      4954: inst = 32'h10408000;
      4955: inst = 32'hc404b34;
      4956: inst = 32'h8220000;
      4957: inst = 32'h10408000;
      4958: inst = 32'hc404b35;
      4959: inst = 32'h8220000;
      4960: inst = 32'h10408000;
      4961: inst = 32'hc404b36;
      4962: inst = 32'h8220000;
      4963: inst = 32'h10408000;
      4964: inst = 32'hc404b37;
      4965: inst = 32'h8220000;
      4966: inst = 32'h10408000;
      4967: inst = 32'hc404b38;
      4968: inst = 32'h8220000;
      4969: inst = 32'h10408000;
      4970: inst = 32'hc404b39;
      4971: inst = 32'h8220000;
      4972: inst = 32'h10408000;
      4973: inst = 32'hc404b3a;
      4974: inst = 32'h8220000;
      4975: inst = 32'h10408000;
      4976: inst = 32'hc404b3b;
      4977: inst = 32'h8220000;
      4978: inst = 32'h10408000;
      4979: inst = 32'hc404b64;
      4980: inst = 32'h8220000;
      4981: inst = 32'h10408000;
      4982: inst = 32'hc404b65;
      4983: inst = 32'h8220000;
      4984: inst = 32'h10408000;
      4985: inst = 32'hc404b66;
      4986: inst = 32'h8220000;
      4987: inst = 32'h10408000;
      4988: inst = 32'hc404b67;
      4989: inst = 32'h8220000;
      4990: inst = 32'h10408000;
      4991: inst = 32'hc404b68;
      4992: inst = 32'h8220000;
      4993: inst = 32'h10408000;
      4994: inst = 32'hc404b69;
      4995: inst = 32'h8220000;
      4996: inst = 32'h10408000;
      4997: inst = 32'hc404b6a;
      4998: inst = 32'h8220000;
      4999: inst = 32'h10408000;
      5000: inst = 32'hc404b6b;
      5001: inst = 32'h8220000;
      5002: inst = 32'h10408000;
      5003: inst = 32'hc404b6c;
      5004: inst = 32'h8220000;
      5005: inst = 32'h10408000;
      5006: inst = 32'hc404b6d;
      5007: inst = 32'h8220000;
      5008: inst = 32'h10408000;
      5009: inst = 32'hc404b6e;
      5010: inst = 32'h8220000;
      5011: inst = 32'h10408000;
      5012: inst = 32'hc404b80;
      5013: inst = 32'h8220000;
      5014: inst = 32'h10408000;
      5015: inst = 32'hc404b81;
      5016: inst = 32'h8220000;
      5017: inst = 32'h10408000;
      5018: inst = 32'hc404b82;
      5019: inst = 32'h8220000;
      5020: inst = 32'h10408000;
      5021: inst = 32'hc404b83;
      5022: inst = 32'h8220000;
      5023: inst = 32'h10408000;
      5024: inst = 32'hc404b84;
      5025: inst = 32'h8220000;
      5026: inst = 32'h10408000;
      5027: inst = 32'hc404b85;
      5028: inst = 32'h8220000;
      5029: inst = 32'h10408000;
      5030: inst = 32'hc404b86;
      5031: inst = 32'h8220000;
      5032: inst = 32'h10408000;
      5033: inst = 32'hc404b90;
      5034: inst = 32'h8220000;
      5035: inst = 32'h10408000;
      5036: inst = 32'hc404b91;
      5037: inst = 32'h8220000;
      5038: inst = 32'h10408000;
      5039: inst = 32'hc404b92;
      5040: inst = 32'h8220000;
      5041: inst = 32'h10408000;
      5042: inst = 32'hc404b93;
      5043: inst = 32'h8220000;
      5044: inst = 32'h10408000;
      5045: inst = 32'hc404b94;
      5046: inst = 32'h8220000;
      5047: inst = 32'h10408000;
      5048: inst = 32'hc404b95;
      5049: inst = 32'h8220000;
      5050: inst = 32'h10408000;
      5051: inst = 32'hc404b96;
      5052: inst = 32'h8220000;
      5053: inst = 32'h10408000;
      5054: inst = 32'hc404b97;
      5055: inst = 32'h8220000;
      5056: inst = 32'h10408000;
      5057: inst = 32'hc404b98;
      5058: inst = 32'h8220000;
      5059: inst = 32'h10408000;
      5060: inst = 32'hc404b99;
      5061: inst = 32'h8220000;
      5062: inst = 32'h10408000;
      5063: inst = 32'hc404b9a;
      5064: inst = 32'h8220000;
      5065: inst = 32'h10408000;
      5066: inst = 32'hc404b9b;
      5067: inst = 32'h8220000;
      5068: inst = 32'h10408000;
      5069: inst = 32'hc404bc4;
      5070: inst = 32'h8220000;
      5071: inst = 32'h10408000;
      5072: inst = 32'hc404bc5;
      5073: inst = 32'h8220000;
      5074: inst = 32'h10408000;
      5075: inst = 32'hc404bc6;
      5076: inst = 32'h8220000;
      5077: inst = 32'h10408000;
      5078: inst = 32'hc404bc7;
      5079: inst = 32'h8220000;
      5080: inst = 32'h10408000;
      5081: inst = 32'hc404bc8;
      5082: inst = 32'h8220000;
      5083: inst = 32'h10408000;
      5084: inst = 32'hc404bc9;
      5085: inst = 32'h8220000;
      5086: inst = 32'h10408000;
      5087: inst = 32'hc404bca;
      5088: inst = 32'h8220000;
      5089: inst = 32'h10408000;
      5090: inst = 32'hc404bcb;
      5091: inst = 32'h8220000;
      5092: inst = 32'h10408000;
      5093: inst = 32'hc404bcc;
      5094: inst = 32'h8220000;
      5095: inst = 32'h10408000;
      5096: inst = 32'hc404bcd;
      5097: inst = 32'h8220000;
      5098: inst = 32'h10408000;
      5099: inst = 32'hc404bce;
      5100: inst = 32'h8220000;
      5101: inst = 32'h10408000;
      5102: inst = 32'hc404be0;
      5103: inst = 32'h8220000;
      5104: inst = 32'h10408000;
      5105: inst = 32'hc404be1;
      5106: inst = 32'h8220000;
      5107: inst = 32'h10408000;
      5108: inst = 32'hc404be2;
      5109: inst = 32'h8220000;
      5110: inst = 32'h10408000;
      5111: inst = 32'hc404be3;
      5112: inst = 32'h8220000;
      5113: inst = 32'h10408000;
      5114: inst = 32'hc404be4;
      5115: inst = 32'h8220000;
      5116: inst = 32'h10408000;
      5117: inst = 32'hc404be5;
      5118: inst = 32'h8220000;
      5119: inst = 32'h10408000;
      5120: inst = 32'hc404be6;
      5121: inst = 32'h8220000;
      5122: inst = 32'h10408000;
      5123: inst = 32'hc404bf0;
      5124: inst = 32'h8220000;
      5125: inst = 32'h10408000;
      5126: inst = 32'hc404bf1;
      5127: inst = 32'h8220000;
      5128: inst = 32'h10408000;
      5129: inst = 32'hc404bf2;
      5130: inst = 32'h8220000;
      5131: inst = 32'h10408000;
      5132: inst = 32'hc404bf3;
      5133: inst = 32'h8220000;
      5134: inst = 32'h10408000;
      5135: inst = 32'hc404bf4;
      5136: inst = 32'h8220000;
      5137: inst = 32'h10408000;
      5138: inst = 32'hc404bf5;
      5139: inst = 32'h8220000;
      5140: inst = 32'h10408000;
      5141: inst = 32'hc404bf6;
      5142: inst = 32'h8220000;
      5143: inst = 32'h10408000;
      5144: inst = 32'hc404bf7;
      5145: inst = 32'h8220000;
      5146: inst = 32'h10408000;
      5147: inst = 32'hc404bf8;
      5148: inst = 32'h8220000;
      5149: inst = 32'h10408000;
      5150: inst = 32'hc404bf9;
      5151: inst = 32'h8220000;
      5152: inst = 32'h10408000;
      5153: inst = 32'hc404c26;
      5154: inst = 32'h8220000;
      5155: inst = 32'h10408000;
      5156: inst = 32'hc404c27;
      5157: inst = 32'h8220000;
      5158: inst = 32'h10408000;
      5159: inst = 32'hc404c28;
      5160: inst = 32'h8220000;
      5161: inst = 32'h10408000;
      5162: inst = 32'hc404c29;
      5163: inst = 32'h8220000;
      5164: inst = 32'h10408000;
      5165: inst = 32'hc404c2a;
      5166: inst = 32'h8220000;
      5167: inst = 32'h10408000;
      5168: inst = 32'hc404c2b;
      5169: inst = 32'h8220000;
      5170: inst = 32'h10408000;
      5171: inst = 32'hc404c2c;
      5172: inst = 32'h8220000;
      5173: inst = 32'h10408000;
      5174: inst = 32'hc404c2d;
      5175: inst = 32'h8220000;
      5176: inst = 32'h10408000;
      5177: inst = 32'hc404c2e;
      5178: inst = 32'h8220000;
      5179: inst = 32'h10408000;
      5180: inst = 32'hc404c40;
      5181: inst = 32'h8220000;
      5182: inst = 32'h10408000;
      5183: inst = 32'hc404c41;
      5184: inst = 32'h8220000;
      5185: inst = 32'h10408000;
      5186: inst = 32'hc404c42;
      5187: inst = 32'h8220000;
      5188: inst = 32'h10408000;
      5189: inst = 32'hc404c43;
      5190: inst = 32'h8220000;
      5191: inst = 32'h10408000;
      5192: inst = 32'hc404c44;
      5193: inst = 32'h8220000;
      5194: inst = 32'h10408000;
      5195: inst = 32'hc404c45;
      5196: inst = 32'h8220000;
      5197: inst = 32'h10408000;
      5198: inst = 32'hc404c46;
      5199: inst = 32'h8220000;
      5200: inst = 32'h10408000;
      5201: inst = 32'hc404c4f;
      5202: inst = 32'h8220000;
      5203: inst = 32'h10408000;
      5204: inst = 32'hc404c50;
      5205: inst = 32'h8220000;
      5206: inst = 32'h10408000;
      5207: inst = 32'hc404c51;
      5208: inst = 32'h8220000;
      5209: inst = 32'h10408000;
      5210: inst = 32'hc404c52;
      5211: inst = 32'h8220000;
      5212: inst = 32'h10408000;
      5213: inst = 32'hc404c53;
      5214: inst = 32'h8220000;
      5215: inst = 32'h10408000;
      5216: inst = 32'hc404c54;
      5217: inst = 32'h8220000;
      5218: inst = 32'h10408000;
      5219: inst = 32'hc404c55;
      5220: inst = 32'h8220000;
      5221: inst = 32'h10408000;
      5222: inst = 32'hc404c56;
      5223: inst = 32'h8220000;
      5224: inst = 32'h10408000;
      5225: inst = 32'hc404c57;
      5226: inst = 32'h8220000;
      5227: inst = 32'h10408000;
      5228: inst = 32'hc404c58;
      5229: inst = 32'h8220000;
      5230: inst = 32'h10408000;
      5231: inst = 32'hc404c59;
      5232: inst = 32'h8220000;
      5233: inst = 32'h10408000;
      5234: inst = 32'hc404c5a;
      5235: inst = 32'h8220000;
      5236: inst = 32'h10408000;
      5237: inst = 32'hc404c5b;
      5238: inst = 32'h8220000;
      5239: inst = 32'h10408000;
      5240: inst = 32'hc404c5c;
      5241: inst = 32'h8220000;
      5242: inst = 32'h10408000;
      5243: inst = 32'hc404c5d;
      5244: inst = 32'h8220000;
      5245: inst = 32'h10408000;
      5246: inst = 32'hc404c5e;
      5247: inst = 32'h8220000;
      5248: inst = 32'h10408000;
      5249: inst = 32'hc404c5f;
      5250: inst = 32'h8220000;
      5251: inst = 32'h10408000;
      5252: inst = 32'hc404c60;
      5253: inst = 32'h8220000;
      5254: inst = 32'h10408000;
      5255: inst = 32'hc404c61;
      5256: inst = 32'h8220000;
      5257: inst = 32'h10408000;
      5258: inst = 32'hc404c62;
      5259: inst = 32'h8220000;
      5260: inst = 32'h10408000;
      5261: inst = 32'hc404c63;
      5262: inst = 32'h8220000;
      5263: inst = 32'h10408000;
      5264: inst = 32'hc404c64;
      5265: inst = 32'h8220000;
      5266: inst = 32'h10408000;
      5267: inst = 32'hc404c65;
      5268: inst = 32'h8220000;
      5269: inst = 32'h10408000;
      5270: inst = 32'hc404c66;
      5271: inst = 32'h8220000;
      5272: inst = 32'h10408000;
      5273: inst = 32'hc404c67;
      5274: inst = 32'h8220000;
      5275: inst = 32'h10408000;
      5276: inst = 32'hc404c68;
      5277: inst = 32'h8220000;
      5278: inst = 32'h10408000;
      5279: inst = 32'hc404c69;
      5280: inst = 32'h8220000;
      5281: inst = 32'h10408000;
      5282: inst = 32'hc404c6a;
      5283: inst = 32'h8220000;
      5284: inst = 32'h10408000;
      5285: inst = 32'hc404c6b;
      5286: inst = 32'h8220000;
      5287: inst = 32'h10408000;
      5288: inst = 32'hc404c6c;
      5289: inst = 32'h8220000;
      5290: inst = 32'h10408000;
      5291: inst = 32'hc404c6d;
      5292: inst = 32'h8220000;
      5293: inst = 32'h10408000;
      5294: inst = 32'hc404c6e;
      5295: inst = 32'h8220000;
      5296: inst = 32'h10408000;
      5297: inst = 32'hc404c6f;
      5298: inst = 32'h8220000;
      5299: inst = 32'h10408000;
      5300: inst = 32'hc404c70;
      5301: inst = 32'h8220000;
      5302: inst = 32'h10408000;
      5303: inst = 32'hc404c71;
      5304: inst = 32'h8220000;
      5305: inst = 32'h10408000;
      5306: inst = 32'hc404c72;
      5307: inst = 32'h8220000;
      5308: inst = 32'h10408000;
      5309: inst = 32'hc404c73;
      5310: inst = 32'h8220000;
      5311: inst = 32'h10408000;
      5312: inst = 32'hc404c74;
      5313: inst = 32'h8220000;
      5314: inst = 32'h10408000;
      5315: inst = 32'hc404c75;
      5316: inst = 32'h8220000;
      5317: inst = 32'h10408000;
      5318: inst = 32'hc404c76;
      5319: inst = 32'h8220000;
      5320: inst = 32'h10408000;
      5321: inst = 32'hc404c77;
      5322: inst = 32'h8220000;
      5323: inst = 32'h10408000;
      5324: inst = 32'hc404c78;
      5325: inst = 32'h8220000;
      5326: inst = 32'h10408000;
      5327: inst = 32'hc404c79;
      5328: inst = 32'h8220000;
      5329: inst = 32'h10408000;
      5330: inst = 32'hc404c7a;
      5331: inst = 32'h8220000;
      5332: inst = 32'h10408000;
      5333: inst = 32'hc404c7b;
      5334: inst = 32'h8220000;
      5335: inst = 32'h10408000;
      5336: inst = 32'hc404c7c;
      5337: inst = 32'h8220000;
      5338: inst = 32'h10408000;
      5339: inst = 32'hc404c7d;
      5340: inst = 32'h8220000;
      5341: inst = 32'h10408000;
      5342: inst = 32'hc404c7e;
      5343: inst = 32'h8220000;
      5344: inst = 32'h10408000;
      5345: inst = 32'hc404c7f;
      5346: inst = 32'h8220000;
      5347: inst = 32'h10408000;
      5348: inst = 32'hc404c80;
      5349: inst = 32'h8220000;
      5350: inst = 32'h10408000;
      5351: inst = 32'hc404c81;
      5352: inst = 32'h8220000;
      5353: inst = 32'h10408000;
      5354: inst = 32'hc404c82;
      5355: inst = 32'h8220000;
      5356: inst = 32'h10408000;
      5357: inst = 32'hc404c83;
      5358: inst = 32'h8220000;
      5359: inst = 32'h10408000;
      5360: inst = 32'hc404c84;
      5361: inst = 32'h8220000;
      5362: inst = 32'h10408000;
      5363: inst = 32'hc404c85;
      5364: inst = 32'h8220000;
      5365: inst = 32'h10408000;
      5366: inst = 32'hc404c86;
      5367: inst = 32'h8220000;
      5368: inst = 32'h10408000;
      5369: inst = 32'hc404c87;
      5370: inst = 32'h8220000;
      5371: inst = 32'h10408000;
      5372: inst = 32'hc404c88;
      5373: inst = 32'h8220000;
      5374: inst = 32'h10408000;
      5375: inst = 32'hc404c89;
      5376: inst = 32'h8220000;
      5377: inst = 32'h10408000;
      5378: inst = 32'hc404c8a;
      5379: inst = 32'h8220000;
      5380: inst = 32'h10408000;
      5381: inst = 32'hc404c8b;
      5382: inst = 32'h8220000;
      5383: inst = 32'h10408000;
      5384: inst = 32'hc404c8c;
      5385: inst = 32'h8220000;
      5386: inst = 32'h10408000;
      5387: inst = 32'hc404c8d;
      5388: inst = 32'h8220000;
      5389: inst = 32'h10408000;
      5390: inst = 32'hc404c8e;
      5391: inst = 32'h8220000;
      5392: inst = 32'h10408000;
      5393: inst = 32'hc404ca0;
      5394: inst = 32'h8220000;
      5395: inst = 32'h10408000;
      5396: inst = 32'hc404ca1;
      5397: inst = 32'h8220000;
      5398: inst = 32'h10408000;
      5399: inst = 32'hc404cb7;
      5400: inst = 32'h8220000;
      5401: inst = 32'h10408000;
      5402: inst = 32'hc404cb8;
      5403: inst = 32'h8220000;
      5404: inst = 32'h10408000;
      5405: inst = 32'hc404cb9;
      5406: inst = 32'h8220000;
      5407: inst = 32'h10408000;
      5408: inst = 32'hc404cba;
      5409: inst = 32'h8220000;
      5410: inst = 32'h10408000;
      5411: inst = 32'hc404cbb;
      5412: inst = 32'h8220000;
      5413: inst = 32'h10408000;
      5414: inst = 32'hc404cbc;
      5415: inst = 32'h8220000;
      5416: inst = 32'h10408000;
      5417: inst = 32'hc404cbd;
      5418: inst = 32'h8220000;
      5419: inst = 32'h10408000;
      5420: inst = 32'hc404cbe;
      5421: inst = 32'h8220000;
      5422: inst = 32'h10408000;
      5423: inst = 32'hc404cbf;
      5424: inst = 32'h8220000;
      5425: inst = 32'h10408000;
      5426: inst = 32'hc404cc0;
      5427: inst = 32'h8220000;
      5428: inst = 32'h10408000;
      5429: inst = 32'hc404cc1;
      5430: inst = 32'h8220000;
      5431: inst = 32'h10408000;
      5432: inst = 32'hc404cc2;
      5433: inst = 32'h8220000;
      5434: inst = 32'h10408000;
      5435: inst = 32'hc404cc3;
      5436: inst = 32'h8220000;
      5437: inst = 32'h10408000;
      5438: inst = 32'hc404cc4;
      5439: inst = 32'h8220000;
      5440: inst = 32'h10408000;
      5441: inst = 32'hc404cc5;
      5442: inst = 32'h8220000;
      5443: inst = 32'h10408000;
      5444: inst = 32'hc404cc6;
      5445: inst = 32'h8220000;
      5446: inst = 32'h10408000;
      5447: inst = 32'hc404cc7;
      5448: inst = 32'h8220000;
      5449: inst = 32'h10408000;
      5450: inst = 32'hc404cc8;
      5451: inst = 32'h8220000;
      5452: inst = 32'h10408000;
      5453: inst = 32'hc404cc9;
      5454: inst = 32'h8220000;
      5455: inst = 32'h10408000;
      5456: inst = 32'hc404cca;
      5457: inst = 32'h8220000;
      5458: inst = 32'h10408000;
      5459: inst = 32'hc404ccb;
      5460: inst = 32'h8220000;
      5461: inst = 32'h10408000;
      5462: inst = 32'hc404ccc;
      5463: inst = 32'h8220000;
      5464: inst = 32'h10408000;
      5465: inst = 32'hc404ccd;
      5466: inst = 32'h8220000;
      5467: inst = 32'h10408000;
      5468: inst = 32'hc404cce;
      5469: inst = 32'h8220000;
      5470: inst = 32'h10408000;
      5471: inst = 32'hc404ccf;
      5472: inst = 32'h8220000;
      5473: inst = 32'h10408000;
      5474: inst = 32'hc404cd0;
      5475: inst = 32'h8220000;
      5476: inst = 32'h10408000;
      5477: inst = 32'hc404cd1;
      5478: inst = 32'h8220000;
      5479: inst = 32'h10408000;
      5480: inst = 32'hc404cd2;
      5481: inst = 32'h8220000;
      5482: inst = 32'h10408000;
      5483: inst = 32'hc404cd3;
      5484: inst = 32'h8220000;
      5485: inst = 32'h10408000;
      5486: inst = 32'hc404cd4;
      5487: inst = 32'h8220000;
      5488: inst = 32'h10408000;
      5489: inst = 32'hc404cd5;
      5490: inst = 32'h8220000;
      5491: inst = 32'h10408000;
      5492: inst = 32'hc404cd6;
      5493: inst = 32'h8220000;
      5494: inst = 32'h10408000;
      5495: inst = 32'hc404cd7;
      5496: inst = 32'h8220000;
      5497: inst = 32'h10408000;
      5498: inst = 32'hc404cd8;
      5499: inst = 32'h8220000;
      5500: inst = 32'h10408000;
      5501: inst = 32'hc404cd9;
      5502: inst = 32'h8220000;
      5503: inst = 32'h10408000;
      5504: inst = 32'hc404cda;
      5505: inst = 32'h8220000;
      5506: inst = 32'h10408000;
      5507: inst = 32'hc404cdb;
      5508: inst = 32'h8220000;
      5509: inst = 32'h10408000;
      5510: inst = 32'hc404cdc;
      5511: inst = 32'h8220000;
      5512: inst = 32'h10408000;
      5513: inst = 32'hc404cdd;
      5514: inst = 32'h8220000;
      5515: inst = 32'h10408000;
      5516: inst = 32'hc404cde;
      5517: inst = 32'h8220000;
      5518: inst = 32'h10408000;
      5519: inst = 32'hc404cdf;
      5520: inst = 32'h8220000;
      5521: inst = 32'h10408000;
      5522: inst = 32'hc404ce0;
      5523: inst = 32'h8220000;
      5524: inst = 32'h10408000;
      5525: inst = 32'hc404ce1;
      5526: inst = 32'h8220000;
      5527: inst = 32'h10408000;
      5528: inst = 32'hc404ce2;
      5529: inst = 32'h8220000;
      5530: inst = 32'h10408000;
      5531: inst = 32'hc404ce3;
      5532: inst = 32'h8220000;
      5533: inst = 32'h10408000;
      5534: inst = 32'hc404ce4;
      5535: inst = 32'h8220000;
      5536: inst = 32'h10408000;
      5537: inst = 32'hc404ce5;
      5538: inst = 32'h8220000;
      5539: inst = 32'h10408000;
      5540: inst = 32'hc404ce6;
      5541: inst = 32'h8220000;
      5542: inst = 32'h10408000;
      5543: inst = 32'hc404ce7;
      5544: inst = 32'h8220000;
      5545: inst = 32'h10408000;
      5546: inst = 32'hc404ce8;
      5547: inst = 32'h8220000;
      5548: inst = 32'h10408000;
      5549: inst = 32'hc404ce9;
      5550: inst = 32'h8220000;
      5551: inst = 32'h10408000;
      5552: inst = 32'hc404cea;
      5553: inst = 32'h8220000;
      5554: inst = 32'h10408000;
      5555: inst = 32'hc404ceb;
      5556: inst = 32'h8220000;
      5557: inst = 32'h10408000;
      5558: inst = 32'hc404cec;
      5559: inst = 32'h8220000;
      5560: inst = 32'h10408000;
      5561: inst = 32'hc404ced;
      5562: inst = 32'h8220000;
      5563: inst = 32'h10408000;
      5564: inst = 32'hc404cee;
      5565: inst = 32'h8220000;
      5566: inst = 32'h10408000;
      5567: inst = 32'hc404d17;
      5568: inst = 32'h8220000;
      5569: inst = 32'h10408000;
      5570: inst = 32'hc404d18;
      5571: inst = 32'h8220000;
      5572: inst = 32'h10408000;
      5573: inst = 32'hc404d19;
      5574: inst = 32'h8220000;
      5575: inst = 32'h10408000;
      5576: inst = 32'hc404d1a;
      5577: inst = 32'h8220000;
      5578: inst = 32'h10408000;
      5579: inst = 32'hc404d1b;
      5580: inst = 32'h8220000;
      5581: inst = 32'h10408000;
      5582: inst = 32'hc404d1c;
      5583: inst = 32'h8220000;
      5584: inst = 32'h10408000;
      5585: inst = 32'hc404d1d;
      5586: inst = 32'h8220000;
      5587: inst = 32'h10408000;
      5588: inst = 32'hc404d1e;
      5589: inst = 32'h8220000;
      5590: inst = 32'h10408000;
      5591: inst = 32'hc404d1f;
      5592: inst = 32'h8220000;
      5593: inst = 32'h10408000;
      5594: inst = 32'hc404d20;
      5595: inst = 32'h8220000;
      5596: inst = 32'h10408000;
      5597: inst = 32'hc404d21;
      5598: inst = 32'h8220000;
      5599: inst = 32'h10408000;
      5600: inst = 32'hc404d22;
      5601: inst = 32'h8220000;
      5602: inst = 32'h10408000;
      5603: inst = 32'hc404d23;
      5604: inst = 32'h8220000;
      5605: inst = 32'h10408000;
      5606: inst = 32'hc404d24;
      5607: inst = 32'h8220000;
      5608: inst = 32'h10408000;
      5609: inst = 32'hc404d25;
      5610: inst = 32'h8220000;
      5611: inst = 32'h10408000;
      5612: inst = 32'hc404d26;
      5613: inst = 32'h8220000;
      5614: inst = 32'h10408000;
      5615: inst = 32'hc404d27;
      5616: inst = 32'h8220000;
      5617: inst = 32'h10408000;
      5618: inst = 32'hc404d28;
      5619: inst = 32'h8220000;
      5620: inst = 32'h10408000;
      5621: inst = 32'hc404d29;
      5622: inst = 32'h8220000;
      5623: inst = 32'h10408000;
      5624: inst = 32'hc404d2a;
      5625: inst = 32'h8220000;
      5626: inst = 32'h10408000;
      5627: inst = 32'hc404d2b;
      5628: inst = 32'h8220000;
      5629: inst = 32'h10408000;
      5630: inst = 32'hc404d2c;
      5631: inst = 32'h8220000;
      5632: inst = 32'h10408000;
      5633: inst = 32'hc404d2d;
      5634: inst = 32'h8220000;
      5635: inst = 32'h10408000;
      5636: inst = 32'hc404d2e;
      5637: inst = 32'h8220000;
      5638: inst = 32'h10408000;
      5639: inst = 32'hc404d2f;
      5640: inst = 32'h8220000;
      5641: inst = 32'h10408000;
      5642: inst = 32'hc404d30;
      5643: inst = 32'h8220000;
      5644: inst = 32'h10408000;
      5645: inst = 32'hc404d31;
      5646: inst = 32'h8220000;
      5647: inst = 32'h10408000;
      5648: inst = 32'hc404d32;
      5649: inst = 32'h8220000;
      5650: inst = 32'h10408000;
      5651: inst = 32'hc404d33;
      5652: inst = 32'h8220000;
      5653: inst = 32'h10408000;
      5654: inst = 32'hc404d34;
      5655: inst = 32'h8220000;
      5656: inst = 32'h10408000;
      5657: inst = 32'hc404d35;
      5658: inst = 32'h8220000;
      5659: inst = 32'h10408000;
      5660: inst = 32'hc404d36;
      5661: inst = 32'h8220000;
      5662: inst = 32'h10408000;
      5663: inst = 32'hc404d37;
      5664: inst = 32'h8220000;
      5665: inst = 32'h10408000;
      5666: inst = 32'hc404d38;
      5667: inst = 32'h8220000;
      5668: inst = 32'h10408000;
      5669: inst = 32'hc404d39;
      5670: inst = 32'h8220000;
      5671: inst = 32'h10408000;
      5672: inst = 32'hc404d3a;
      5673: inst = 32'h8220000;
      5674: inst = 32'h10408000;
      5675: inst = 32'hc404d3b;
      5676: inst = 32'h8220000;
      5677: inst = 32'h10408000;
      5678: inst = 32'hc404d3c;
      5679: inst = 32'h8220000;
      5680: inst = 32'h10408000;
      5681: inst = 32'hc404d3d;
      5682: inst = 32'h8220000;
      5683: inst = 32'h10408000;
      5684: inst = 32'hc404d3e;
      5685: inst = 32'h8220000;
      5686: inst = 32'h10408000;
      5687: inst = 32'hc404d3f;
      5688: inst = 32'h8220000;
      5689: inst = 32'h10408000;
      5690: inst = 32'hc404d40;
      5691: inst = 32'h8220000;
      5692: inst = 32'h10408000;
      5693: inst = 32'hc404d41;
      5694: inst = 32'h8220000;
      5695: inst = 32'h10408000;
      5696: inst = 32'hc404d42;
      5697: inst = 32'h8220000;
      5698: inst = 32'h10408000;
      5699: inst = 32'hc404d43;
      5700: inst = 32'h8220000;
      5701: inst = 32'h10408000;
      5702: inst = 32'hc404d44;
      5703: inst = 32'h8220000;
      5704: inst = 32'h10408000;
      5705: inst = 32'hc404d45;
      5706: inst = 32'h8220000;
      5707: inst = 32'h10408000;
      5708: inst = 32'hc404d46;
      5709: inst = 32'h8220000;
      5710: inst = 32'h10408000;
      5711: inst = 32'hc404d47;
      5712: inst = 32'h8220000;
      5713: inst = 32'h10408000;
      5714: inst = 32'hc404d48;
      5715: inst = 32'h8220000;
      5716: inst = 32'h10408000;
      5717: inst = 32'hc404d49;
      5718: inst = 32'h8220000;
      5719: inst = 32'h10408000;
      5720: inst = 32'hc404d4a;
      5721: inst = 32'h8220000;
      5722: inst = 32'h10408000;
      5723: inst = 32'hc404d4b;
      5724: inst = 32'h8220000;
      5725: inst = 32'h10408000;
      5726: inst = 32'hc404d4c;
      5727: inst = 32'h8220000;
      5728: inst = 32'h10408000;
      5729: inst = 32'hc404d4d;
      5730: inst = 32'h8220000;
      5731: inst = 32'h10408000;
      5732: inst = 32'hc404d4e;
      5733: inst = 32'h8220000;
      5734: inst = 32'h10408000;
      5735: inst = 32'hc404d77;
      5736: inst = 32'h8220000;
      5737: inst = 32'h10408000;
      5738: inst = 32'hc404d78;
      5739: inst = 32'h8220000;
      5740: inst = 32'h10408000;
      5741: inst = 32'hc404d79;
      5742: inst = 32'h8220000;
      5743: inst = 32'h10408000;
      5744: inst = 32'hc404d7a;
      5745: inst = 32'h8220000;
      5746: inst = 32'h10408000;
      5747: inst = 32'hc404d7b;
      5748: inst = 32'h8220000;
      5749: inst = 32'h10408000;
      5750: inst = 32'hc404d7c;
      5751: inst = 32'h8220000;
      5752: inst = 32'h10408000;
      5753: inst = 32'hc404d7d;
      5754: inst = 32'h8220000;
      5755: inst = 32'h10408000;
      5756: inst = 32'hc404d7e;
      5757: inst = 32'h8220000;
      5758: inst = 32'h10408000;
      5759: inst = 32'hc404d7f;
      5760: inst = 32'h8220000;
      5761: inst = 32'h10408000;
      5762: inst = 32'hc404d80;
      5763: inst = 32'h8220000;
      5764: inst = 32'h10408000;
      5765: inst = 32'hc404d81;
      5766: inst = 32'h8220000;
      5767: inst = 32'h10408000;
      5768: inst = 32'hc404d82;
      5769: inst = 32'h8220000;
      5770: inst = 32'h10408000;
      5771: inst = 32'hc404d83;
      5772: inst = 32'h8220000;
      5773: inst = 32'h10408000;
      5774: inst = 32'hc404d84;
      5775: inst = 32'h8220000;
      5776: inst = 32'h10408000;
      5777: inst = 32'hc404d85;
      5778: inst = 32'h8220000;
      5779: inst = 32'h10408000;
      5780: inst = 32'hc404d86;
      5781: inst = 32'h8220000;
      5782: inst = 32'h10408000;
      5783: inst = 32'hc404d87;
      5784: inst = 32'h8220000;
      5785: inst = 32'h10408000;
      5786: inst = 32'hc404d88;
      5787: inst = 32'h8220000;
      5788: inst = 32'h10408000;
      5789: inst = 32'hc404d89;
      5790: inst = 32'h8220000;
      5791: inst = 32'h10408000;
      5792: inst = 32'hc404d8a;
      5793: inst = 32'h8220000;
      5794: inst = 32'h10408000;
      5795: inst = 32'hc404d8b;
      5796: inst = 32'h8220000;
      5797: inst = 32'h10408000;
      5798: inst = 32'hc404d8c;
      5799: inst = 32'h8220000;
      5800: inst = 32'h10408000;
      5801: inst = 32'hc404d8d;
      5802: inst = 32'h8220000;
      5803: inst = 32'h10408000;
      5804: inst = 32'hc404d8e;
      5805: inst = 32'h8220000;
      5806: inst = 32'h10408000;
      5807: inst = 32'hc404d8f;
      5808: inst = 32'h8220000;
      5809: inst = 32'h10408000;
      5810: inst = 32'hc404d90;
      5811: inst = 32'h8220000;
      5812: inst = 32'h10408000;
      5813: inst = 32'hc404d91;
      5814: inst = 32'h8220000;
      5815: inst = 32'h10408000;
      5816: inst = 32'hc404d92;
      5817: inst = 32'h8220000;
      5818: inst = 32'h10408000;
      5819: inst = 32'hc404d93;
      5820: inst = 32'h8220000;
      5821: inst = 32'h10408000;
      5822: inst = 32'hc404d94;
      5823: inst = 32'h8220000;
      5824: inst = 32'h10408000;
      5825: inst = 32'hc404d95;
      5826: inst = 32'h8220000;
      5827: inst = 32'h10408000;
      5828: inst = 32'hc404d96;
      5829: inst = 32'h8220000;
      5830: inst = 32'h10408000;
      5831: inst = 32'hc404d97;
      5832: inst = 32'h8220000;
      5833: inst = 32'h10408000;
      5834: inst = 32'hc404d98;
      5835: inst = 32'h8220000;
      5836: inst = 32'h10408000;
      5837: inst = 32'hc404d99;
      5838: inst = 32'h8220000;
      5839: inst = 32'h10408000;
      5840: inst = 32'hc404d9a;
      5841: inst = 32'h8220000;
      5842: inst = 32'h10408000;
      5843: inst = 32'hc404d9b;
      5844: inst = 32'h8220000;
      5845: inst = 32'h10408000;
      5846: inst = 32'hc404d9c;
      5847: inst = 32'h8220000;
      5848: inst = 32'h10408000;
      5849: inst = 32'hc404d9d;
      5850: inst = 32'h8220000;
      5851: inst = 32'h10408000;
      5852: inst = 32'hc404d9e;
      5853: inst = 32'h8220000;
      5854: inst = 32'h10408000;
      5855: inst = 32'hc404d9f;
      5856: inst = 32'h8220000;
      5857: inst = 32'h10408000;
      5858: inst = 32'hc404da0;
      5859: inst = 32'h8220000;
      5860: inst = 32'h10408000;
      5861: inst = 32'hc404da1;
      5862: inst = 32'h8220000;
      5863: inst = 32'h10408000;
      5864: inst = 32'hc404da2;
      5865: inst = 32'h8220000;
      5866: inst = 32'h10408000;
      5867: inst = 32'hc404da3;
      5868: inst = 32'h8220000;
      5869: inst = 32'h10408000;
      5870: inst = 32'hc404da4;
      5871: inst = 32'h8220000;
      5872: inst = 32'h10408000;
      5873: inst = 32'hc404da5;
      5874: inst = 32'h8220000;
      5875: inst = 32'h10408000;
      5876: inst = 32'hc404da6;
      5877: inst = 32'h8220000;
      5878: inst = 32'h10408000;
      5879: inst = 32'hc404da7;
      5880: inst = 32'h8220000;
      5881: inst = 32'h10408000;
      5882: inst = 32'hc404da8;
      5883: inst = 32'h8220000;
      5884: inst = 32'h10408000;
      5885: inst = 32'hc404da9;
      5886: inst = 32'h8220000;
      5887: inst = 32'h10408000;
      5888: inst = 32'hc404daa;
      5889: inst = 32'h8220000;
      5890: inst = 32'h10408000;
      5891: inst = 32'hc404dab;
      5892: inst = 32'h8220000;
      5893: inst = 32'h10408000;
      5894: inst = 32'hc404dac;
      5895: inst = 32'h8220000;
      5896: inst = 32'h10408000;
      5897: inst = 32'hc404dad;
      5898: inst = 32'h8220000;
      5899: inst = 32'h10408000;
      5900: inst = 32'hc404dae;
      5901: inst = 32'h8220000;
      5902: inst = 32'h10408000;
      5903: inst = 32'hc404dd7;
      5904: inst = 32'h8220000;
      5905: inst = 32'h10408000;
      5906: inst = 32'hc404dd8;
      5907: inst = 32'h8220000;
      5908: inst = 32'h10408000;
      5909: inst = 32'hc404dd9;
      5910: inst = 32'h8220000;
      5911: inst = 32'h10408000;
      5912: inst = 32'hc404dda;
      5913: inst = 32'h8220000;
      5914: inst = 32'h10408000;
      5915: inst = 32'hc404ddb;
      5916: inst = 32'h8220000;
      5917: inst = 32'h10408000;
      5918: inst = 32'hc404ddc;
      5919: inst = 32'h8220000;
      5920: inst = 32'h10408000;
      5921: inst = 32'hc404ddd;
      5922: inst = 32'h8220000;
      5923: inst = 32'h10408000;
      5924: inst = 32'hc404dde;
      5925: inst = 32'h8220000;
      5926: inst = 32'h10408000;
      5927: inst = 32'hc404ddf;
      5928: inst = 32'h8220000;
      5929: inst = 32'h10408000;
      5930: inst = 32'hc404de0;
      5931: inst = 32'h8220000;
      5932: inst = 32'h10408000;
      5933: inst = 32'hc404de1;
      5934: inst = 32'h8220000;
      5935: inst = 32'h10408000;
      5936: inst = 32'hc404de2;
      5937: inst = 32'h8220000;
      5938: inst = 32'h10408000;
      5939: inst = 32'hc404de3;
      5940: inst = 32'h8220000;
      5941: inst = 32'h10408000;
      5942: inst = 32'hc404de4;
      5943: inst = 32'h8220000;
      5944: inst = 32'h10408000;
      5945: inst = 32'hc404de5;
      5946: inst = 32'h8220000;
      5947: inst = 32'h10408000;
      5948: inst = 32'hc404de6;
      5949: inst = 32'h8220000;
      5950: inst = 32'h10408000;
      5951: inst = 32'hc404de7;
      5952: inst = 32'h8220000;
      5953: inst = 32'h10408000;
      5954: inst = 32'hc404de8;
      5955: inst = 32'h8220000;
      5956: inst = 32'h10408000;
      5957: inst = 32'hc404de9;
      5958: inst = 32'h8220000;
      5959: inst = 32'h10408000;
      5960: inst = 32'hc404dea;
      5961: inst = 32'h8220000;
      5962: inst = 32'h10408000;
      5963: inst = 32'hc404deb;
      5964: inst = 32'h8220000;
      5965: inst = 32'h10408000;
      5966: inst = 32'hc404dec;
      5967: inst = 32'h8220000;
      5968: inst = 32'h10408000;
      5969: inst = 32'hc404ded;
      5970: inst = 32'h8220000;
      5971: inst = 32'h10408000;
      5972: inst = 32'hc404dee;
      5973: inst = 32'h8220000;
      5974: inst = 32'h10408000;
      5975: inst = 32'hc404def;
      5976: inst = 32'h8220000;
      5977: inst = 32'h10408000;
      5978: inst = 32'hc404df0;
      5979: inst = 32'h8220000;
      5980: inst = 32'h10408000;
      5981: inst = 32'hc404df1;
      5982: inst = 32'h8220000;
      5983: inst = 32'h10408000;
      5984: inst = 32'hc404df2;
      5985: inst = 32'h8220000;
      5986: inst = 32'h10408000;
      5987: inst = 32'hc404df3;
      5988: inst = 32'h8220000;
      5989: inst = 32'h10408000;
      5990: inst = 32'hc404df4;
      5991: inst = 32'h8220000;
      5992: inst = 32'h10408000;
      5993: inst = 32'hc404df5;
      5994: inst = 32'h8220000;
      5995: inst = 32'h10408000;
      5996: inst = 32'hc404df6;
      5997: inst = 32'h8220000;
      5998: inst = 32'h10408000;
      5999: inst = 32'hc404df7;
      6000: inst = 32'h8220000;
      6001: inst = 32'h10408000;
      6002: inst = 32'hc404df8;
      6003: inst = 32'h8220000;
      6004: inst = 32'h10408000;
      6005: inst = 32'hc404df9;
      6006: inst = 32'h8220000;
      6007: inst = 32'h10408000;
      6008: inst = 32'hc404dfa;
      6009: inst = 32'h8220000;
      6010: inst = 32'h10408000;
      6011: inst = 32'hc404dfb;
      6012: inst = 32'h8220000;
      6013: inst = 32'h10408000;
      6014: inst = 32'hc404dfc;
      6015: inst = 32'h8220000;
      6016: inst = 32'h10408000;
      6017: inst = 32'hc404dfd;
      6018: inst = 32'h8220000;
      6019: inst = 32'h10408000;
      6020: inst = 32'hc404dfe;
      6021: inst = 32'h8220000;
      6022: inst = 32'h10408000;
      6023: inst = 32'hc404dff;
      6024: inst = 32'h8220000;
      6025: inst = 32'h10408000;
      6026: inst = 32'hc404e00;
      6027: inst = 32'h8220000;
      6028: inst = 32'h10408000;
      6029: inst = 32'hc404e01;
      6030: inst = 32'h8220000;
      6031: inst = 32'h10408000;
      6032: inst = 32'hc404e02;
      6033: inst = 32'h8220000;
      6034: inst = 32'h10408000;
      6035: inst = 32'hc404e03;
      6036: inst = 32'h8220000;
      6037: inst = 32'h10408000;
      6038: inst = 32'hc404e04;
      6039: inst = 32'h8220000;
      6040: inst = 32'h10408000;
      6041: inst = 32'hc404e05;
      6042: inst = 32'h8220000;
      6043: inst = 32'h10408000;
      6044: inst = 32'hc404e06;
      6045: inst = 32'h8220000;
      6046: inst = 32'h10408000;
      6047: inst = 32'hc404e07;
      6048: inst = 32'h8220000;
      6049: inst = 32'h10408000;
      6050: inst = 32'hc404e08;
      6051: inst = 32'h8220000;
      6052: inst = 32'h10408000;
      6053: inst = 32'hc404e09;
      6054: inst = 32'h8220000;
      6055: inst = 32'h10408000;
      6056: inst = 32'hc404e0a;
      6057: inst = 32'h8220000;
      6058: inst = 32'h10408000;
      6059: inst = 32'hc404e0b;
      6060: inst = 32'h8220000;
      6061: inst = 32'h10408000;
      6062: inst = 32'hc404e0c;
      6063: inst = 32'h8220000;
      6064: inst = 32'h10408000;
      6065: inst = 32'hc404e0d;
      6066: inst = 32'h8220000;
      6067: inst = 32'h10408000;
      6068: inst = 32'hc404e0e;
      6069: inst = 32'h8220000;
      6070: inst = 32'h10408000;
      6071: inst = 32'hc404e37;
      6072: inst = 32'h8220000;
      6073: inst = 32'h10408000;
      6074: inst = 32'hc404e38;
      6075: inst = 32'h8220000;
      6076: inst = 32'h10408000;
      6077: inst = 32'hc404e39;
      6078: inst = 32'h8220000;
      6079: inst = 32'h10408000;
      6080: inst = 32'hc404e3a;
      6081: inst = 32'h8220000;
      6082: inst = 32'h10408000;
      6083: inst = 32'hc404e3b;
      6084: inst = 32'h8220000;
      6085: inst = 32'h10408000;
      6086: inst = 32'hc404e3c;
      6087: inst = 32'h8220000;
      6088: inst = 32'h10408000;
      6089: inst = 32'hc404e3d;
      6090: inst = 32'h8220000;
      6091: inst = 32'h10408000;
      6092: inst = 32'hc404e3e;
      6093: inst = 32'h8220000;
      6094: inst = 32'h10408000;
      6095: inst = 32'hc404e3f;
      6096: inst = 32'h8220000;
      6097: inst = 32'h10408000;
      6098: inst = 32'hc404e40;
      6099: inst = 32'h8220000;
      6100: inst = 32'h10408000;
      6101: inst = 32'hc404e41;
      6102: inst = 32'h8220000;
      6103: inst = 32'h10408000;
      6104: inst = 32'hc404e42;
      6105: inst = 32'h8220000;
      6106: inst = 32'h10408000;
      6107: inst = 32'hc404e43;
      6108: inst = 32'h8220000;
      6109: inst = 32'h10408000;
      6110: inst = 32'hc404e44;
      6111: inst = 32'h8220000;
      6112: inst = 32'h10408000;
      6113: inst = 32'hc404e45;
      6114: inst = 32'h8220000;
      6115: inst = 32'h10408000;
      6116: inst = 32'hc404e46;
      6117: inst = 32'h8220000;
      6118: inst = 32'h10408000;
      6119: inst = 32'hc404e47;
      6120: inst = 32'h8220000;
      6121: inst = 32'h10408000;
      6122: inst = 32'hc404e48;
      6123: inst = 32'h8220000;
      6124: inst = 32'h10408000;
      6125: inst = 32'hc404e49;
      6126: inst = 32'h8220000;
      6127: inst = 32'h10408000;
      6128: inst = 32'hc404e4a;
      6129: inst = 32'h8220000;
      6130: inst = 32'h10408000;
      6131: inst = 32'hc404e4b;
      6132: inst = 32'h8220000;
      6133: inst = 32'h10408000;
      6134: inst = 32'hc404e4c;
      6135: inst = 32'h8220000;
      6136: inst = 32'h10408000;
      6137: inst = 32'hc404e4d;
      6138: inst = 32'h8220000;
      6139: inst = 32'h10408000;
      6140: inst = 32'hc404e4e;
      6141: inst = 32'h8220000;
      6142: inst = 32'h10408000;
      6143: inst = 32'hc404e4f;
      6144: inst = 32'h8220000;
      6145: inst = 32'h10408000;
      6146: inst = 32'hc404e50;
      6147: inst = 32'h8220000;
      6148: inst = 32'h10408000;
      6149: inst = 32'hc404e51;
      6150: inst = 32'h8220000;
      6151: inst = 32'h10408000;
      6152: inst = 32'hc404e52;
      6153: inst = 32'h8220000;
      6154: inst = 32'h10408000;
      6155: inst = 32'hc404e53;
      6156: inst = 32'h8220000;
      6157: inst = 32'h10408000;
      6158: inst = 32'hc404e54;
      6159: inst = 32'h8220000;
      6160: inst = 32'h10408000;
      6161: inst = 32'hc404e55;
      6162: inst = 32'h8220000;
      6163: inst = 32'h10408000;
      6164: inst = 32'hc404e56;
      6165: inst = 32'h8220000;
      6166: inst = 32'h10408000;
      6167: inst = 32'hc404e57;
      6168: inst = 32'h8220000;
      6169: inst = 32'h10408000;
      6170: inst = 32'hc404e58;
      6171: inst = 32'h8220000;
      6172: inst = 32'h10408000;
      6173: inst = 32'hc404e59;
      6174: inst = 32'h8220000;
      6175: inst = 32'h10408000;
      6176: inst = 32'hc404e5a;
      6177: inst = 32'h8220000;
      6178: inst = 32'h10408000;
      6179: inst = 32'hc404e5b;
      6180: inst = 32'h8220000;
      6181: inst = 32'h10408000;
      6182: inst = 32'hc404e5c;
      6183: inst = 32'h8220000;
      6184: inst = 32'h10408000;
      6185: inst = 32'hc404e5d;
      6186: inst = 32'h8220000;
      6187: inst = 32'h10408000;
      6188: inst = 32'hc404e5e;
      6189: inst = 32'h8220000;
      6190: inst = 32'h10408000;
      6191: inst = 32'hc404e5f;
      6192: inst = 32'h8220000;
      6193: inst = 32'h10408000;
      6194: inst = 32'hc404e60;
      6195: inst = 32'h8220000;
      6196: inst = 32'h10408000;
      6197: inst = 32'hc404e61;
      6198: inst = 32'h8220000;
      6199: inst = 32'h10408000;
      6200: inst = 32'hc404e62;
      6201: inst = 32'h8220000;
      6202: inst = 32'h10408000;
      6203: inst = 32'hc404e63;
      6204: inst = 32'h8220000;
      6205: inst = 32'h10408000;
      6206: inst = 32'hc404e64;
      6207: inst = 32'h8220000;
      6208: inst = 32'h10408000;
      6209: inst = 32'hc404e65;
      6210: inst = 32'h8220000;
      6211: inst = 32'h10408000;
      6212: inst = 32'hc404e66;
      6213: inst = 32'h8220000;
      6214: inst = 32'h10408000;
      6215: inst = 32'hc404e67;
      6216: inst = 32'h8220000;
      6217: inst = 32'h10408000;
      6218: inst = 32'hc404e68;
      6219: inst = 32'h8220000;
      6220: inst = 32'h10408000;
      6221: inst = 32'hc404e69;
      6222: inst = 32'h8220000;
      6223: inst = 32'h10408000;
      6224: inst = 32'hc404e6a;
      6225: inst = 32'h8220000;
      6226: inst = 32'h10408000;
      6227: inst = 32'hc404e6b;
      6228: inst = 32'h8220000;
      6229: inst = 32'h10408000;
      6230: inst = 32'hc404e6c;
      6231: inst = 32'h8220000;
      6232: inst = 32'h10408000;
      6233: inst = 32'hc404e6d;
      6234: inst = 32'h8220000;
      6235: inst = 32'h10408000;
      6236: inst = 32'hc404e6e;
      6237: inst = 32'h8220000;
      6238: inst = 32'h10408000;
      6239: inst = 32'hc404e97;
      6240: inst = 32'h8220000;
      6241: inst = 32'h10408000;
      6242: inst = 32'hc404e98;
      6243: inst = 32'h8220000;
      6244: inst = 32'h10408000;
      6245: inst = 32'hc404e99;
      6246: inst = 32'h8220000;
      6247: inst = 32'h10408000;
      6248: inst = 32'hc404e9a;
      6249: inst = 32'h8220000;
      6250: inst = 32'h10408000;
      6251: inst = 32'hc404e9b;
      6252: inst = 32'h8220000;
      6253: inst = 32'h10408000;
      6254: inst = 32'hc404e9c;
      6255: inst = 32'h8220000;
      6256: inst = 32'h10408000;
      6257: inst = 32'hc404e9d;
      6258: inst = 32'h8220000;
      6259: inst = 32'h10408000;
      6260: inst = 32'hc404e9e;
      6261: inst = 32'h8220000;
      6262: inst = 32'h10408000;
      6263: inst = 32'hc404ea8;
      6264: inst = 32'h8220000;
      6265: inst = 32'h10408000;
      6266: inst = 32'hc404ea9;
      6267: inst = 32'h8220000;
      6268: inst = 32'h10408000;
      6269: inst = 32'hc404eaa;
      6270: inst = 32'h8220000;
      6271: inst = 32'h10408000;
      6272: inst = 32'hc404eab;
      6273: inst = 32'h8220000;
      6274: inst = 32'h10408000;
      6275: inst = 32'hc404eac;
      6276: inst = 32'h8220000;
      6277: inst = 32'h10408000;
      6278: inst = 32'hc404ead;
      6279: inst = 32'h8220000;
      6280: inst = 32'h10408000;
      6281: inst = 32'hc404eae;
      6282: inst = 32'h8220000;
      6283: inst = 32'h10408000;
      6284: inst = 32'hc404eaf;
      6285: inst = 32'h8220000;
      6286: inst = 32'h10408000;
      6287: inst = 32'hc404eb0;
      6288: inst = 32'h8220000;
      6289: inst = 32'h10408000;
      6290: inst = 32'hc404eb1;
      6291: inst = 32'h8220000;
      6292: inst = 32'h10408000;
      6293: inst = 32'hc404eb2;
      6294: inst = 32'h8220000;
      6295: inst = 32'h10408000;
      6296: inst = 32'hc404eb3;
      6297: inst = 32'h8220000;
      6298: inst = 32'h10408000;
      6299: inst = 32'hc404eb4;
      6300: inst = 32'h8220000;
      6301: inst = 32'h10408000;
      6302: inst = 32'hc404eb5;
      6303: inst = 32'h8220000;
      6304: inst = 32'h10408000;
      6305: inst = 32'hc404eb6;
      6306: inst = 32'h8220000;
      6307: inst = 32'h10408000;
      6308: inst = 32'hc404eb7;
      6309: inst = 32'h8220000;
      6310: inst = 32'h10408000;
      6311: inst = 32'hc404ec1;
      6312: inst = 32'h8220000;
      6313: inst = 32'h10408000;
      6314: inst = 32'hc404ec2;
      6315: inst = 32'h8220000;
      6316: inst = 32'h10408000;
      6317: inst = 32'hc404ec3;
      6318: inst = 32'h8220000;
      6319: inst = 32'h10408000;
      6320: inst = 32'hc404ec4;
      6321: inst = 32'h8220000;
      6322: inst = 32'h10408000;
      6323: inst = 32'hc404ec5;
      6324: inst = 32'h8220000;
      6325: inst = 32'h10408000;
      6326: inst = 32'hc404ec6;
      6327: inst = 32'h8220000;
      6328: inst = 32'h10408000;
      6329: inst = 32'hc404ec7;
      6330: inst = 32'h8220000;
      6331: inst = 32'h10408000;
      6332: inst = 32'hc404ec8;
      6333: inst = 32'h8220000;
      6334: inst = 32'h10408000;
      6335: inst = 32'hc404ec9;
      6336: inst = 32'h8220000;
      6337: inst = 32'h10408000;
      6338: inst = 32'hc404eca;
      6339: inst = 32'h8220000;
      6340: inst = 32'h10408000;
      6341: inst = 32'hc404ecb;
      6342: inst = 32'h8220000;
      6343: inst = 32'h10408000;
      6344: inst = 32'hc404ecc;
      6345: inst = 32'h8220000;
      6346: inst = 32'h10408000;
      6347: inst = 32'hc404ecd;
      6348: inst = 32'h8220000;
      6349: inst = 32'h10408000;
      6350: inst = 32'hc404ece;
      6351: inst = 32'h8220000;
      6352: inst = 32'h10408000;
      6353: inst = 32'hc404ef7;
      6354: inst = 32'h8220000;
      6355: inst = 32'h10408000;
      6356: inst = 32'hc404ef8;
      6357: inst = 32'h8220000;
      6358: inst = 32'h10408000;
      6359: inst = 32'hc404ef9;
      6360: inst = 32'h8220000;
      6361: inst = 32'h10408000;
      6362: inst = 32'hc404efa;
      6363: inst = 32'h8220000;
      6364: inst = 32'h10408000;
      6365: inst = 32'hc404efb;
      6366: inst = 32'h8220000;
      6367: inst = 32'h10408000;
      6368: inst = 32'hc404efc;
      6369: inst = 32'h8220000;
      6370: inst = 32'h10408000;
      6371: inst = 32'hc404efd;
      6372: inst = 32'h8220000;
      6373: inst = 32'h10408000;
      6374: inst = 32'hc404efe;
      6375: inst = 32'h8220000;
      6376: inst = 32'h10408000;
      6377: inst = 32'hc404f08;
      6378: inst = 32'h8220000;
      6379: inst = 32'h10408000;
      6380: inst = 32'hc404f09;
      6381: inst = 32'h8220000;
      6382: inst = 32'h10408000;
      6383: inst = 32'hc404f0a;
      6384: inst = 32'h8220000;
      6385: inst = 32'h10408000;
      6386: inst = 32'hc404f0b;
      6387: inst = 32'h8220000;
      6388: inst = 32'h10408000;
      6389: inst = 32'hc404f0c;
      6390: inst = 32'h8220000;
      6391: inst = 32'h10408000;
      6392: inst = 32'hc404f0d;
      6393: inst = 32'h8220000;
      6394: inst = 32'h10408000;
      6395: inst = 32'hc404f0e;
      6396: inst = 32'h8220000;
      6397: inst = 32'h10408000;
      6398: inst = 32'hc404f0f;
      6399: inst = 32'h8220000;
      6400: inst = 32'h10408000;
      6401: inst = 32'hc404f10;
      6402: inst = 32'h8220000;
      6403: inst = 32'h10408000;
      6404: inst = 32'hc404f11;
      6405: inst = 32'h8220000;
      6406: inst = 32'h10408000;
      6407: inst = 32'hc404f12;
      6408: inst = 32'h8220000;
      6409: inst = 32'h10408000;
      6410: inst = 32'hc404f13;
      6411: inst = 32'h8220000;
      6412: inst = 32'h10408000;
      6413: inst = 32'hc404f14;
      6414: inst = 32'h8220000;
      6415: inst = 32'h10408000;
      6416: inst = 32'hc404f15;
      6417: inst = 32'h8220000;
      6418: inst = 32'h10408000;
      6419: inst = 32'hc404f16;
      6420: inst = 32'h8220000;
      6421: inst = 32'h10408000;
      6422: inst = 32'hc404f17;
      6423: inst = 32'h8220000;
      6424: inst = 32'h10408000;
      6425: inst = 32'hc404f21;
      6426: inst = 32'h8220000;
      6427: inst = 32'h10408000;
      6428: inst = 32'hc404f22;
      6429: inst = 32'h8220000;
      6430: inst = 32'h10408000;
      6431: inst = 32'hc404f23;
      6432: inst = 32'h8220000;
      6433: inst = 32'h10408000;
      6434: inst = 32'hc404f24;
      6435: inst = 32'h8220000;
      6436: inst = 32'h10408000;
      6437: inst = 32'hc404f25;
      6438: inst = 32'h8220000;
      6439: inst = 32'h10408000;
      6440: inst = 32'hc404f26;
      6441: inst = 32'h8220000;
      6442: inst = 32'h10408000;
      6443: inst = 32'hc404f27;
      6444: inst = 32'h8220000;
      6445: inst = 32'h10408000;
      6446: inst = 32'hc404f28;
      6447: inst = 32'h8220000;
      6448: inst = 32'h10408000;
      6449: inst = 32'hc404f29;
      6450: inst = 32'h8220000;
      6451: inst = 32'h10408000;
      6452: inst = 32'hc404f2a;
      6453: inst = 32'h8220000;
      6454: inst = 32'h10408000;
      6455: inst = 32'hc404f2b;
      6456: inst = 32'h8220000;
      6457: inst = 32'h10408000;
      6458: inst = 32'hc404f2c;
      6459: inst = 32'h8220000;
      6460: inst = 32'h10408000;
      6461: inst = 32'hc404f2d;
      6462: inst = 32'h8220000;
      6463: inst = 32'h10408000;
      6464: inst = 32'hc404f2e;
      6465: inst = 32'h8220000;
      6466: inst = 32'h10408000;
      6467: inst = 32'hc404f57;
      6468: inst = 32'h8220000;
      6469: inst = 32'h10408000;
      6470: inst = 32'hc404f58;
      6471: inst = 32'h8220000;
      6472: inst = 32'h10408000;
      6473: inst = 32'hc404f59;
      6474: inst = 32'h8220000;
      6475: inst = 32'h10408000;
      6476: inst = 32'hc404f5a;
      6477: inst = 32'h8220000;
      6478: inst = 32'h10408000;
      6479: inst = 32'hc404f5b;
      6480: inst = 32'h8220000;
      6481: inst = 32'h10408000;
      6482: inst = 32'hc404f5c;
      6483: inst = 32'h8220000;
      6484: inst = 32'h10408000;
      6485: inst = 32'hc404f5d;
      6486: inst = 32'h8220000;
      6487: inst = 32'h10408000;
      6488: inst = 32'hc404f5e;
      6489: inst = 32'h8220000;
      6490: inst = 32'h10408000;
      6491: inst = 32'hc404f68;
      6492: inst = 32'h8220000;
      6493: inst = 32'h10408000;
      6494: inst = 32'hc404f69;
      6495: inst = 32'h8220000;
      6496: inst = 32'h10408000;
      6497: inst = 32'hc404f6a;
      6498: inst = 32'h8220000;
      6499: inst = 32'h10408000;
      6500: inst = 32'hc404f6b;
      6501: inst = 32'h8220000;
      6502: inst = 32'h10408000;
      6503: inst = 32'hc404f6c;
      6504: inst = 32'h8220000;
      6505: inst = 32'h10408000;
      6506: inst = 32'hc404f6d;
      6507: inst = 32'h8220000;
      6508: inst = 32'h10408000;
      6509: inst = 32'hc404f6e;
      6510: inst = 32'h8220000;
      6511: inst = 32'h10408000;
      6512: inst = 32'hc404f6f;
      6513: inst = 32'h8220000;
      6514: inst = 32'h10408000;
      6515: inst = 32'hc404f70;
      6516: inst = 32'h8220000;
      6517: inst = 32'h10408000;
      6518: inst = 32'hc404f71;
      6519: inst = 32'h8220000;
      6520: inst = 32'h10408000;
      6521: inst = 32'hc404f72;
      6522: inst = 32'h8220000;
      6523: inst = 32'h10408000;
      6524: inst = 32'hc404f73;
      6525: inst = 32'h8220000;
      6526: inst = 32'h10408000;
      6527: inst = 32'hc404f74;
      6528: inst = 32'h8220000;
      6529: inst = 32'h10408000;
      6530: inst = 32'hc404f75;
      6531: inst = 32'h8220000;
      6532: inst = 32'h10408000;
      6533: inst = 32'hc404f76;
      6534: inst = 32'h8220000;
      6535: inst = 32'h10408000;
      6536: inst = 32'hc404f77;
      6537: inst = 32'h8220000;
      6538: inst = 32'h10408000;
      6539: inst = 32'hc404f81;
      6540: inst = 32'h8220000;
      6541: inst = 32'h10408000;
      6542: inst = 32'hc404f82;
      6543: inst = 32'h8220000;
      6544: inst = 32'h10408000;
      6545: inst = 32'hc404f83;
      6546: inst = 32'h8220000;
      6547: inst = 32'h10408000;
      6548: inst = 32'hc404f84;
      6549: inst = 32'h8220000;
      6550: inst = 32'h10408000;
      6551: inst = 32'hc404f85;
      6552: inst = 32'h8220000;
      6553: inst = 32'h10408000;
      6554: inst = 32'hc404f86;
      6555: inst = 32'h8220000;
      6556: inst = 32'h10408000;
      6557: inst = 32'hc404f87;
      6558: inst = 32'h8220000;
      6559: inst = 32'h10408000;
      6560: inst = 32'hc404f88;
      6561: inst = 32'h8220000;
      6562: inst = 32'h10408000;
      6563: inst = 32'hc404f89;
      6564: inst = 32'h8220000;
      6565: inst = 32'h10408000;
      6566: inst = 32'hc404f8a;
      6567: inst = 32'h8220000;
      6568: inst = 32'h10408000;
      6569: inst = 32'hc404f8b;
      6570: inst = 32'h8220000;
      6571: inst = 32'h10408000;
      6572: inst = 32'hc404f8c;
      6573: inst = 32'h8220000;
      6574: inst = 32'h10408000;
      6575: inst = 32'hc404f8d;
      6576: inst = 32'h8220000;
      6577: inst = 32'h10408000;
      6578: inst = 32'hc404f8e;
      6579: inst = 32'h8220000;
      6580: inst = 32'h10408000;
      6581: inst = 32'hc404fb7;
      6582: inst = 32'h8220000;
      6583: inst = 32'h10408000;
      6584: inst = 32'hc404fb8;
      6585: inst = 32'h8220000;
      6586: inst = 32'h10408000;
      6587: inst = 32'hc404fb9;
      6588: inst = 32'h8220000;
      6589: inst = 32'h10408000;
      6590: inst = 32'hc404fba;
      6591: inst = 32'h8220000;
      6592: inst = 32'h10408000;
      6593: inst = 32'hc404fbb;
      6594: inst = 32'h8220000;
      6595: inst = 32'h10408000;
      6596: inst = 32'hc404fbc;
      6597: inst = 32'h8220000;
      6598: inst = 32'h10408000;
      6599: inst = 32'hc404fbd;
      6600: inst = 32'h8220000;
      6601: inst = 32'h10408000;
      6602: inst = 32'hc404fbe;
      6603: inst = 32'h8220000;
      6604: inst = 32'h10408000;
      6605: inst = 32'hc404fc8;
      6606: inst = 32'h8220000;
      6607: inst = 32'h10408000;
      6608: inst = 32'hc404fc9;
      6609: inst = 32'h8220000;
      6610: inst = 32'h10408000;
      6611: inst = 32'hc404fca;
      6612: inst = 32'h8220000;
      6613: inst = 32'h10408000;
      6614: inst = 32'hc404fcb;
      6615: inst = 32'h8220000;
      6616: inst = 32'h10408000;
      6617: inst = 32'hc404fcc;
      6618: inst = 32'h8220000;
      6619: inst = 32'h10408000;
      6620: inst = 32'hc404fcd;
      6621: inst = 32'h8220000;
      6622: inst = 32'h10408000;
      6623: inst = 32'hc404fce;
      6624: inst = 32'h8220000;
      6625: inst = 32'h10408000;
      6626: inst = 32'hc404fcf;
      6627: inst = 32'h8220000;
      6628: inst = 32'h10408000;
      6629: inst = 32'hc404fd0;
      6630: inst = 32'h8220000;
      6631: inst = 32'h10408000;
      6632: inst = 32'hc404fd1;
      6633: inst = 32'h8220000;
      6634: inst = 32'h10408000;
      6635: inst = 32'hc404fd2;
      6636: inst = 32'h8220000;
      6637: inst = 32'h10408000;
      6638: inst = 32'hc404fd3;
      6639: inst = 32'h8220000;
      6640: inst = 32'h10408000;
      6641: inst = 32'hc404fd4;
      6642: inst = 32'h8220000;
      6643: inst = 32'h10408000;
      6644: inst = 32'hc404fd5;
      6645: inst = 32'h8220000;
      6646: inst = 32'h10408000;
      6647: inst = 32'hc404fd6;
      6648: inst = 32'h8220000;
      6649: inst = 32'h10408000;
      6650: inst = 32'hc404fd7;
      6651: inst = 32'h8220000;
      6652: inst = 32'h10408000;
      6653: inst = 32'hc404fe1;
      6654: inst = 32'h8220000;
      6655: inst = 32'h10408000;
      6656: inst = 32'hc404fe2;
      6657: inst = 32'h8220000;
      6658: inst = 32'h10408000;
      6659: inst = 32'hc404fe3;
      6660: inst = 32'h8220000;
      6661: inst = 32'h10408000;
      6662: inst = 32'hc404fe4;
      6663: inst = 32'h8220000;
      6664: inst = 32'h10408000;
      6665: inst = 32'hc404fe5;
      6666: inst = 32'h8220000;
      6667: inst = 32'h10408000;
      6668: inst = 32'hc404fe6;
      6669: inst = 32'h8220000;
      6670: inst = 32'h10408000;
      6671: inst = 32'hc404fe7;
      6672: inst = 32'h8220000;
      6673: inst = 32'h10408000;
      6674: inst = 32'hc404fe8;
      6675: inst = 32'h8220000;
      6676: inst = 32'h10408000;
      6677: inst = 32'hc404fe9;
      6678: inst = 32'h8220000;
      6679: inst = 32'h10408000;
      6680: inst = 32'hc404fea;
      6681: inst = 32'h8220000;
      6682: inst = 32'h10408000;
      6683: inst = 32'hc404feb;
      6684: inst = 32'h8220000;
      6685: inst = 32'h10408000;
      6686: inst = 32'hc404fec;
      6687: inst = 32'h8220000;
      6688: inst = 32'h10408000;
      6689: inst = 32'hc404fed;
      6690: inst = 32'h8220000;
      6691: inst = 32'h10408000;
      6692: inst = 32'hc404fee;
      6693: inst = 32'h8220000;
      6694: inst = 32'h10408000;
      6695: inst = 32'hc405017;
      6696: inst = 32'h8220000;
      6697: inst = 32'h10408000;
      6698: inst = 32'hc405018;
      6699: inst = 32'h8220000;
      6700: inst = 32'h10408000;
      6701: inst = 32'hc405019;
      6702: inst = 32'h8220000;
      6703: inst = 32'h10408000;
      6704: inst = 32'hc40501a;
      6705: inst = 32'h8220000;
      6706: inst = 32'h10408000;
      6707: inst = 32'hc40501b;
      6708: inst = 32'h8220000;
      6709: inst = 32'h10408000;
      6710: inst = 32'hc40501c;
      6711: inst = 32'h8220000;
      6712: inst = 32'h10408000;
      6713: inst = 32'hc40501d;
      6714: inst = 32'h8220000;
      6715: inst = 32'h10408000;
      6716: inst = 32'hc40501e;
      6717: inst = 32'h8220000;
      6718: inst = 32'h10408000;
      6719: inst = 32'hc405028;
      6720: inst = 32'h8220000;
      6721: inst = 32'h10408000;
      6722: inst = 32'hc405029;
      6723: inst = 32'h8220000;
      6724: inst = 32'h10408000;
      6725: inst = 32'hc40502a;
      6726: inst = 32'h8220000;
      6727: inst = 32'h10408000;
      6728: inst = 32'hc40502b;
      6729: inst = 32'h8220000;
      6730: inst = 32'h10408000;
      6731: inst = 32'hc40502c;
      6732: inst = 32'h8220000;
      6733: inst = 32'h10408000;
      6734: inst = 32'hc40502d;
      6735: inst = 32'h8220000;
      6736: inst = 32'h10408000;
      6737: inst = 32'hc40502e;
      6738: inst = 32'h8220000;
      6739: inst = 32'h10408000;
      6740: inst = 32'hc40502f;
      6741: inst = 32'h8220000;
      6742: inst = 32'h10408000;
      6743: inst = 32'hc405030;
      6744: inst = 32'h8220000;
      6745: inst = 32'h10408000;
      6746: inst = 32'hc405031;
      6747: inst = 32'h8220000;
      6748: inst = 32'h10408000;
      6749: inst = 32'hc405032;
      6750: inst = 32'h8220000;
      6751: inst = 32'h10408000;
      6752: inst = 32'hc405033;
      6753: inst = 32'h8220000;
      6754: inst = 32'h10408000;
      6755: inst = 32'hc405034;
      6756: inst = 32'h8220000;
      6757: inst = 32'h10408000;
      6758: inst = 32'hc405035;
      6759: inst = 32'h8220000;
      6760: inst = 32'h10408000;
      6761: inst = 32'hc405036;
      6762: inst = 32'h8220000;
      6763: inst = 32'h10408000;
      6764: inst = 32'hc405037;
      6765: inst = 32'h8220000;
      6766: inst = 32'h10408000;
      6767: inst = 32'hc405041;
      6768: inst = 32'h8220000;
      6769: inst = 32'h10408000;
      6770: inst = 32'hc405042;
      6771: inst = 32'h8220000;
      6772: inst = 32'h10408000;
      6773: inst = 32'hc405043;
      6774: inst = 32'h8220000;
      6775: inst = 32'h10408000;
      6776: inst = 32'hc405044;
      6777: inst = 32'h8220000;
      6778: inst = 32'h10408000;
      6779: inst = 32'hc405045;
      6780: inst = 32'h8220000;
      6781: inst = 32'h10408000;
      6782: inst = 32'hc405046;
      6783: inst = 32'h8220000;
      6784: inst = 32'h10408000;
      6785: inst = 32'hc405047;
      6786: inst = 32'h8220000;
      6787: inst = 32'h10408000;
      6788: inst = 32'hc405048;
      6789: inst = 32'h8220000;
      6790: inst = 32'h10408000;
      6791: inst = 32'hc405049;
      6792: inst = 32'h8220000;
      6793: inst = 32'h10408000;
      6794: inst = 32'hc40504a;
      6795: inst = 32'h8220000;
      6796: inst = 32'h10408000;
      6797: inst = 32'hc40504b;
      6798: inst = 32'h8220000;
      6799: inst = 32'h10408000;
      6800: inst = 32'hc40504c;
      6801: inst = 32'h8220000;
      6802: inst = 32'h10408000;
      6803: inst = 32'hc40504d;
      6804: inst = 32'h8220000;
      6805: inst = 32'h10408000;
      6806: inst = 32'hc40504e;
      6807: inst = 32'h8220000;
      6808: inst = 32'h10408000;
      6809: inst = 32'hc405077;
      6810: inst = 32'h8220000;
      6811: inst = 32'h10408000;
      6812: inst = 32'hc405078;
      6813: inst = 32'h8220000;
      6814: inst = 32'h10408000;
      6815: inst = 32'hc405079;
      6816: inst = 32'h8220000;
      6817: inst = 32'h10408000;
      6818: inst = 32'hc40507a;
      6819: inst = 32'h8220000;
      6820: inst = 32'h10408000;
      6821: inst = 32'hc40507b;
      6822: inst = 32'h8220000;
      6823: inst = 32'h10408000;
      6824: inst = 32'hc40507c;
      6825: inst = 32'h8220000;
      6826: inst = 32'h10408000;
      6827: inst = 32'hc40507d;
      6828: inst = 32'h8220000;
      6829: inst = 32'h10408000;
      6830: inst = 32'hc40507e;
      6831: inst = 32'h8220000;
      6832: inst = 32'h10408000;
      6833: inst = 32'hc405088;
      6834: inst = 32'h8220000;
      6835: inst = 32'h10408000;
      6836: inst = 32'hc405089;
      6837: inst = 32'h8220000;
      6838: inst = 32'h10408000;
      6839: inst = 32'hc40508a;
      6840: inst = 32'h8220000;
      6841: inst = 32'h10408000;
      6842: inst = 32'hc40508b;
      6843: inst = 32'h8220000;
      6844: inst = 32'h10408000;
      6845: inst = 32'hc40508c;
      6846: inst = 32'h8220000;
      6847: inst = 32'h10408000;
      6848: inst = 32'hc40508d;
      6849: inst = 32'h8220000;
      6850: inst = 32'h10408000;
      6851: inst = 32'hc40508e;
      6852: inst = 32'h8220000;
      6853: inst = 32'h10408000;
      6854: inst = 32'hc40508f;
      6855: inst = 32'h8220000;
      6856: inst = 32'h10408000;
      6857: inst = 32'hc405090;
      6858: inst = 32'h8220000;
      6859: inst = 32'h10408000;
      6860: inst = 32'hc405091;
      6861: inst = 32'h8220000;
      6862: inst = 32'h10408000;
      6863: inst = 32'hc405092;
      6864: inst = 32'h8220000;
      6865: inst = 32'h10408000;
      6866: inst = 32'hc405093;
      6867: inst = 32'h8220000;
      6868: inst = 32'h10408000;
      6869: inst = 32'hc405094;
      6870: inst = 32'h8220000;
      6871: inst = 32'h10408000;
      6872: inst = 32'hc405095;
      6873: inst = 32'h8220000;
      6874: inst = 32'h10408000;
      6875: inst = 32'hc405096;
      6876: inst = 32'h8220000;
      6877: inst = 32'h10408000;
      6878: inst = 32'hc405097;
      6879: inst = 32'h8220000;
      6880: inst = 32'h10408000;
      6881: inst = 32'hc4050a1;
      6882: inst = 32'h8220000;
      6883: inst = 32'h10408000;
      6884: inst = 32'hc4050a2;
      6885: inst = 32'h8220000;
      6886: inst = 32'h10408000;
      6887: inst = 32'hc4050a3;
      6888: inst = 32'h8220000;
      6889: inst = 32'h10408000;
      6890: inst = 32'hc4050a4;
      6891: inst = 32'h8220000;
      6892: inst = 32'h10408000;
      6893: inst = 32'hc4050a5;
      6894: inst = 32'h8220000;
      6895: inst = 32'h10408000;
      6896: inst = 32'hc4050a6;
      6897: inst = 32'h8220000;
      6898: inst = 32'h10408000;
      6899: inst = 32'hc4050a7;
      6900: inst = 32'h8220000;
      6901: inst = 32'h10408000;
      6902: inst = 32'hc4050a8;
      6903: inst = 32'h8220000;
      6904: inst = 32'h10408000;
      6905: inst = 32'hc4050a9;
      6906: inst = 32'h8220000;
      6907: inst = 32'h10408000;
      6908: inst = 32'hc4050aa;
      6909: inst = 32'h8220000;
      6910: inst = 32'h10408000;
      6911: inst = 32'hc4050ab;
      6912: inst = 32'h8220000;
      6913: inst = 32'h10408000;
      6914: inst = 32'hc4050ac;
      6915: inst = 32'h8220000;
      6916: inst = 32'h10408000;
      6917: inst = 32'hc4050ad;
      6918: inst = 32'h8220000;
      6919: inst = 32'h10408000;
      6920: inst = 32'hc4050ae;
      6921: inst = 32'h8220000;
      6922: inst = 32'h10408000;
      6923: inst = 32'hc4050d7;
      6924: inst = 32'h8220000;
      6925: inst = 32'h10408000;
      6926: inst = 32'hc4050d8;
      6927: inst = 32'h8220000;
      6928: inst = 32'h10408000;
      6929: inst = 32'hc4050d9;
      6930: inst = 32'h8220000;
      6931: inst = 32'h10408000;
      6932: inst = 32'hc4050da;
      6933: inst = 32'h8220000;
      6934: inst = 32'h10408000;
      6935: inst = 32'hc4050db;
      6936: inst = 32'h8220000;
      6937: inst = 32'h10408000;
      6938: inst = 32'hc4050dc;
      6939: inst = 32'h8220000;
      6940: inst = 32'h10408000;
      6941: inst = 32'hc4050dd;
      6942: inst = 32'h8220000;
      6943: inst = 32'h10408000;
      6944: inst = 32'hc4050de;
      6945: inst = 32'h8220000;
      6946: inst = 32'h10408000;
      6947: inst = 32'hc4050e8;
      6948: inst = 32'h8220000;
      6949: inst = 32'h10408000;
      6950: inst = 32'hc4050e9;
      6951: inst = 32'h8220000;
      6952: inst = 32'h10408000;
      6953: inst = 32'hc4050ea;
      6954: inst = 32'h8220000;
      6955: inst = 32'h10408000;
      6956: inst = 32'hc4050eb;
      6957: inst = 32'h8220000;
      6958: inst = 32'h10408000;
      6959: inst = 32'hc4050ec;
      6960: inst = 32'h8220000;
      6961: inst = 32'h10408000;
      6962: inst = 32'hc4050ed;
      6963: inst = 32'h8220000;
      6964: inst = 32'h10408000;
      6965: inst = 32'hc4050ee;
      6966: inst = 32'h8220000;
      6967: inst = 32'h10408000;
      6968: inst = 32'hc4050ef;
      6969: inst = 32'h8220000;
      6970: inst = 32'h10408000;
      6971: inst = 32'hc4050f0;
      6972: inst = 32'h8220000;
      6973: inst = 32'h10408000;
      6974: inst = 32'hc4050f1;
      6975: inst = 32'h8220000;
      6976: inst = 32'h10408000;
      6977: inst = 32'hc4050f2;
      6978: inst = 32'h8220000;
      6979: inst = 32'h10408000;
      6980: inst = 32'hc4050f3;
      6981: inst = 32'h8220000;
      6982: inst = 32'h10408000;
      6983: inst = 32'hc4050f4;
      6984: inst = 32'h8220000;
      6985: inst = 32'h10408000;
      6986: inst = 32'hc4050f5;
      6987: inst = 32'h8220000;
      6988: inst = 32'h10408000;
      6989: inst = 32'hc4050f6;
      6990: inst = 32'h8220000;
      6991: inst = 32'h10408000;
      6992: inst = 32'hc4050f7;
      6993: inst = 32'h8220000;
      6994: inst = 32'h10408000;
      6995: inst = 32'hc405101;
      6996: inst = 32'h8220000;
      6997: inst = 32'h10408000;
      6998: inst = 32'hc405102;
      6999: inst = 32'h8220000;
      7000: inst = 32'h10408000;
      7001: inst = 32'hc405103;
      7002: inst = 32'h8220000;
      7003: inst = 32'h10408000;
      7004: inst = 32'hc405104;
      7005: inst = 32'h8220000;
      7006: inst = 32'h10408000;
      7007: inst = 32'hc405105;
      7008: inst = 32'h8220000;
      7009: inst = 32'h10408000;
      7010: inst = 32'hc405106;
      7011: inst = 32'h8220000;
      7012: inst = 32'h10408000;
      7013: inst = 32'hc405107;
      7014: inst = 32'h8220000;
      7015: inst = 32'h10408000;
      7016: inst = 32'hc405108;
      7017: inst = 32'h8220000;
      7018: inst = 32'h10408000;
      7019: inst = 32'hc405109;
      7020: inst = 32'h8220000;
      7021: inst = 32'h10408000;
      7022: inst = 32'hc40510a;
      7023: inst = 32'h8220000;
      7024: inst = 32'h10408000;
      7025: inst = 32'hc40510b;
      7026: inst = 32'h8220000;
      7027: inst = 32'h10408000;
      7028: inst = 32'hc40510c;
      7029: inst = 32'h8220000;
      7030: inst = 32'h10408000;
      7031: inst = 32'hc40510d;
      7032: inst = 32'h8220000;
      7033: inst = 32'h10408000;
      7034: inst = 32'hc40510e;
      7035: inst = 32'h8220000;
      7036: inst = 32'h10408000;
      7037: inst = 32'hc405137;
      7038: inst = 32'h8220000;
      7039: inst = 32'h10408000;
      7040: inst = 32'hc405138;
      7041: inst = 32'h8220000;
      7042: inst = 32'h10408000;
      7043: inst = 32'hc405139;
      7044: inst = 32'h8220000;
      7045: inst = 32'h10408000;
      7046: inst = 32'hc40513a;
      7047: inst = 32'h8220000;
      7048: inst = 32'h10408000;
      7049: inst = 32'hc40513b;
      7050: inst = 32'h8220000;
      7051: inst = 32'h10408000;
      7052: inst = 32'hc40513c;
      7053: inst = 32'h8220000;
      7054: inst = 32'h10408000;
      7055: inst = 32'hc40513d;
      7056: inst = 32'h8220000;
      7057: inst = 32'h10408000;
      7058: inst = 32'hc40513e;
      7059: inst = 32'h8220000;
      7060: inst = 32'h10408000;
      7061: inst = 32'hc405148;
      7062: inst = 32'h8220000;
      7063: inst = 32'h10408000;
      7064: inst = 32'hc405149;
      7065: inst = 32'h8220000;
      7066: inst = 32'h10408000;
      7067: inst = 32'hc40514a;
      7068: inst = 32'h8220000;
      7069: inst = 32'h10408000;
      7070: inst = 32'hc40514b;
      7071: inst = 32'h8220000;
      7072: inst = 32'h10408000;
      7073: inst = 32'hc40514c;
      7074: inst = 32'h8220000;
      7075: inst = 32'h10408000;
      7076: inst = 32'hc40514d;
      7077: inst = 32'h8220000;
      7078: inst = 32'h10408000;
      7079: inst = 32'hc40514e;
      7080: inst = 32'h8220000;
      7081: inst = 32'h10408000;
      7082: inst = 32'hc40514f;
      7083: inst = 32'h8220000;
      7084: inst = 32'h10408000;
      7085: inst = 32'hc405150;
      7086: inst = 32'h8220000;
      7087: inst = 32'h10408000;
      7088: inst = 32'hc405151;
      7089: inst = 32'h8220000;
      7090: inst = 32'h10408000;
      7091: inst = 32'hc405152;
      7092: inst = 32'h8220000;
      7093: inst = 32'h10408000;
      7094: inst = 32'hc405153;
      7095: inst = 32'h8220000;
      7096: inst = 32'h10408000;
      7097: inst = 32'hc405154;
      7098: inst = 32'h8220000;
      7099: inst = 32'h10408000;
      7100: inst = 32'hc405155;
      7101: inst = 32'h8220000;
      7102: inst = 32'h10408000;
      7103: inst = 32'hc405156;
      7104: inst = 32'h8220000;
      7105: inst = 32'h10408000;
      7106: inst = 32'hc405157;
      7107: inst = 32'h8220000;
      7108: inst = 32'h10408000;
      7109: inst = 32'hc405161;
      7110: inst = 32'h8220000;
      7111: inst = 32'h10408000;
      7112: inst = 32'hc405162;
      7113: inst = 32'h8220000;
      7114: inst = 32'h10408000;
      7115: inst = 32'hc405163;
      7116: inst = 32'h8220000;
      7117: inst = 32'h10408000;
      7118: inst = 32'hc405164;
      7119: inst = 32'h8220000;
      7120: inst = 32'h10408000;
      7121: inst = 32'hc405165;
      7122: inst = 32'h8220000;
      7123: inst = 32'h10408000;
      7124: inst = 32'hc405166;
      7125: inst = 32'h8220000;
      7126: inst = 32'h10408000;
      7127: inst = 32'hc405167;
      7128: inst = 32'h8220000;
      7129: inst = 32'h10408000;
      7130: inst = 32'hc405168;
      7131: inst = 32'h8220000;
      7132: inst = 32'h10408000;
      7133: inst = 32'hc405169;
      7134: inst = 32'h8220000;
      7135: inst = 32'h10408000;
      7136: inst = 32'hc40516a;
      7137: inst = 32'h8220000;
      7138: inst = 32'h10408000;
      7139: inst = 32'hc40516b;
      7140: inst = 32'h8220000;
      7141: inst = 32'h10408000;
      7142: inst = 32'hc40516c;
      7143: inst = 32'h8220000;
      7144: inst = 32'h10408000;
      7145: inst = 32'hc40516d;
      7146: inst = 32'h8220000;
      7147: inst = 32'h10408000;
      7148: inst = 32'hc40516e;
      7149: inst = 32'h8220000;
      7150: inst = 32'h10408000;
      7151: inst = 32'hc405197;
      7152: inst = 32'h8220000;
      7153: inst = 32'h10408000;
      7154: inst = 32'hc405198;
      7155: inst = 32'h8220000;
      7156: inst = 32'h10408000;
      7157: inst = 32'hc405199;
      7158: inst = 32'h8220000;
      7159: inst = 32'h10408000;
      7160: inst = 32'hc40519a;
      7161: inst = 32'h8220000;
      7162: inst = 32'h10408000;
      7163: inst = 32'hc40519b;
      7164: inst = 32'h8220000;
      7165: inst = 32'h10408000;
      7166: inst = 32'hc40519c;
      7167: inst = 32'h8220000;
      7168: inst = 32'h10408000;
      7169: inst = 32'hc40519d;
      7170: inst = 32'h8220000;
      7171: inst = 32'h10408000;
      7172: inst = 32'hc4051aa;
      7173: inst = 32'h8220000;
      7174: inst = 32'h10408000;
      7175: inst = 32'hc4051ab;
      7176: inst = 32'h8220000;
      7177: inst = 32'h10408000;
      7178: inst = 32'hc4051ac;
      7179: inst = 32'h8220000;
      7180: inst = 32'h10408000;
      7181: inst = 32'hc4051ad;
      7182: inst = 32'h8220000;
      7183: inst = 32'h10408000;
      7184: inst = 32'hc4051ae;
      7185: inst = 32'h8220000;
      7186: inst = 32'h10408000;
      7187: inst = 32'hc4051af;
      7188: inst = 32'h8220000;
      7189: inst = 32'h10408000;
      7190: inst = 32'hc4051b0;
      7191: inst = 32'h8220000;
      7192: inst = 32'h10408000;
      7193: inst = 32'hc4051b1;
      7194: inst = 32'h8220000;
      7195: inst = 32'h10408000;
      7196: inst = 32'hc4051b2;
      7197: inst = 32'h8220000;
      7198: inst = 32'h10408000;
      7199: inst = 32'hc4051b3;
      7200: inst = 32'h8220000;
      7201: inst = 32'h10408000;
      7202: inst = 32'hc4051b4;
      7203: inst = 32'h8220000;
      7204: inst = 32'h10408000;
      7205: inst = 32'hc4051b5;
      7206: inst = 32'h8220000;
      7207: inst = 32'h10408000;
      7208: inst = 32'hc4051c2;
      7209: inst = 32'h8220000;
      7210: inst = 32'h10408000;
      7211: inst = 32'hc4051c3;
      7212: inst = 32'h8220000;
      7213: inst = 32'h10408000;
      7214: inst = 32'hc4051c4;
      7215: inst = 32'h8220000;
      7216: inst = 32'h10408000;
      7217: inst = 32'hc4051c5;
      7218: inst = 32'h8220000;
      7219: inst = 32'h10408000;
      7220: inst = 32'hc4051c6;
      7221: inst = 32'h8220000;
      7222: inst = 32'h10408000;
      7223: inst = 32'hc4051c7;
      7224: inst = 32'h8220000;
      7225: inst = 32'h10408000;
      7226: inst = 32'hc4051c8;
      7227: inst = 32'h8220000;
      7228: inst = 32'h10408000;
      7229: inst = 32'hc4051c9;
      7230: inst = 32'h8220000;
      7231: inst = 32'h10408000;
      7232: inst = 32'hc4051ca;
      7233: inst = 32'h8220000;
      7234: inst = 32'h10408000;
      7235: inst = 32'hc4051cb;
      7236: inst = 32'h8220000;
      7237: inst = 32'h10408000;
      7238: inst = 32'hc4051cc;
      7239: inst = 32'h8220000;
      7240: inst = 32'h10408000;
      7241: inst = 32'hc4051cd;
      7242: inst = 32'h8220000;
      7243: inst = 32'h10408000;
      7244: inst = 32'hc4051ce;
      7245: inst = 32'h8220000;
      7246: inst = 32'h10408000;
      7247: inst = 32'hc4051f7;
      7248: inst = 32'h8220000;
      7249: inst = 32'h10408000;
      7250: inst = 32'hc4051f8;
      7251: inst = 32'h8220000;
      7252: inst = 32'h10408000;
      7253: inst = 32'hc4051f9;
      7254: inst = 32'h8220000;
      7255: inst = 32'h10408000;
      7256: inst = 32'hc4051fa;
      7257: inst = 32'h8220000;
      7258: inst = 32'h10408000;
      7259: inst = 32'hc4051fb;
      7260: inst = 32'h8220000;
      7261: inst = 32'h10408000;
      7262: inst = 32'hc4051fc;
      7263: inst = 32'h8220000;
      7264: inst = 32'h10408000;
      7265: inst = 32'hc40520a;
      7266: inst = 32'h8220000;
      7267: inst = 32'h10408000;
      7268: inst = 32'hc40520b;
      7269: inst = 32'h8220000;
      7270: inst = 32'h10408000;
      7271: inst = 32'hc40520c;
      7272: inst = 32'h8220000;
      7273: inst = 32'h10408000;
      7274: inst = 32'hc40520d;
      7275: inst = 32'h8220000;
      7276: inst = 32'h10408000;
      7277: inst = 32'hc40520e;
      7278: inst = 32'h8220000;
      7279: inst = 32'h10408000;
      7280: inst = 32'hc40520f;
      7281: inst = 32'h8220000;
      7282: inst = 32'h10408000;
      7283: inst = 32'hc405210;
      7284: inst = 32'h8220000;
      7285: inst = 32'h10408000;
      7286: inst = 32'hc405211;
      7287: inst = 32'h8220000;
      7288: inst = 32'h10408000;
      7289: inst = 32'hc405212;
      7290: inst = 32'h8220000;
      7291: inst = 32'h10408000;
      7292: inst = 32'hc405213;
      7293: inst = 32'h8220000;
      7294: inst = 32'h10408000;
      7295: inst = 32'hc405214;
      7296: inst = 32'h8220000;
      7297: inst = 32'h10408000;
      7298: inst = 32'hc405215;
      7299: inst = 32'h8220000;
      7300: inst = 32'h10408000;
      7301: inst = 32'hc405223;
      7302: inst = 32'h8220000;
      7303: inst = 32'h10408000;
      7304: inst = 32'hc405224;
      7305: inst = 32'h8220000;
      7306: inst = 32'h10408000;
      7307: inst = 32'hc405225;
      7308: inst = 32'h8220000;
      7309: inst = 32'h10408000;
      7310: inst = 32'hc405226;
      7311: inst = 32'h8220000;
      7312: inst = 32'h10408000;
      7313: inst = 32'hc405227;
      7314: inst = 32'h8220000;
      7315: inst = 32'h10408000;
      7316: inst = 32'hc405228;
      7317: inst = 32'h8220000;
      7318: inst = 32'h10408000;
      7319: inst = 32'hc405229;
      7320: inst = 32'h8220000;
      7321: inst = 32'h10408000;
      7322: inst = 32'hc40522a;
      7323: inst = 32'h8220000;
      7324: inst = 32'h10408000;
      7325: inst = 32'hc40522b;
      7326: inst = 32'h8220000;
      7327: inst = 32'h10408000;
      7328: inst = 32'hc40522c;
      7329: inst = 32'h8220000;
      7330: inst = 32'h10408000;
      7331: inst = 32'hc40522d;
      7332: inst = 32'h8220000;
      7333: inst = 32'h10408000;
      7334: inst = 32'hc40522e;
      7335: inst = 32'h8220000;
      7336: inst = 32'h10408000;
      7337: inst = 32'hc405257;
      7338: inst = 32'h8220000;
      7339: inst = 32'h10408000;
      7340: inst = 32'hc405258;
      7341: inst = 32'h8220000;
      7342: inst = 32'h10408000;
      7343: inst = 32'hc405259;
      7344: inst = 32'h8220000;
      7345: inst = 32'h10408000;
      7346: inst = 32'hc40525a;
      7347: inst = 32'h8220000;
      7348: inst = 32'h10408000;
      7349: inst = 32'hc40525b;
      7350: inst = 32'h8220000;
      7351: inst = 32'h10408000;
      7352: inst = 32'hc40526a;
      7353: inst = 32'h8220000;
      7354: inst = 32'h10408000;
      7355: inst = 32'hc40526b;
      7356: inst = 32'h8220000;
      7357: inst = 32'h10408000;
      7358: inst = 32'hc40526c;
      7359: inst = 32'h8220000;
      7360: inst = 32'h10408000;
      7361: inst = 32'hc40526d;
      7362: inst = 32'h8220000;
      7363: inst = 32'h10408000;
      7364: inst = 32'hc40526e;
      7365: inst = 32'h8220000;
      7366: inst = 32'h10408000;
      7367: inst = 32'hc40526f;
      7368: inst = 32'h8220000;
      7369: inst = 32'h10408000;
      7370: inst = 32'hc405270;
      7371: inst = 32'h8220000;
      7372: inst = 32'h10408000;
      7373: inst = 32'hc405271;
      7374: inst = 32'h8220000;
      7375: inst = 32'h10408000;
      7376: inst = 32'hc405272;
      7377: inst = 32'h8220000;
      7378: inst = 32'h10408000;
      7379: inst = 32'hc405273;
      7380: inst = 32'h8220000;
      7381: inst = 32'h10408000;
      7382: inst = 32'hc405274;
      7383: inst = 32'h8220000;
      7384: inst = 32'h10408000;
      7385: inst = 32'hc405275;
      7386: inst = 32'h8220000;
      7387: inst = 32'h10408000;
      7388: inst = 32'hc405284;
      7389: inst = 32'h8220000;
      7390: inst = 32'h10408000;
      7391: inst = 32'hc405285;
      7392: inst = 32'h8220000;
      7393: inst = 32'h10408000;
      7394: inst = 32'hc405286;
      7395: inst = 32'h8220000;
      7396: inst = 32'h10408000;
      7397: inst = 32'hc405287;
      7398: inst = 32'h8220000;
      7399: inst = 32'h10408000;
      7400: inst = 32'hc405288;
      7401: inst = 32'h8220000;
      7402: inst = 32'h10408000;
      7403: inst = 32'hc405289;
      7404: inst = 32'h8220000;
      7405: inst = 32'h10408000;
      7406: inst = 32'hc40528a;
      7407: inst = 32'h8220000;
      7408: inst = 32'h10408000;
      7409: inst = 32'hc40528b;
      7410: inst = 32'h8220000;
      7411: inst = 32'h10408000;
      7412: inst = 32'hc40528c;
      7413: inst = 32'h8220000;
      7414: inst = 32'h10408000;
      7415: inst = 32'hc40528d;
      7416: inst = 32'h8220000;
      7417: inst = 32'h10408000;
      7418: inst = 32'hc40528e;
      7419: inst = 32'h8220000;
      7420: inst = 32'h10408000;
      7421: inst = 32'hc4052b7;
      7422: inst = 32'h8220000;
      7423: inst = 32'h10408000;
      7424: inst = 32'hc4052b8;
      7425: inst = 32'h8220000;
      7426: inst = 32'h10408000;
      7427: inst = 32'hc4052b9;
      7428: inst = 32'h8220000;
      7429: inst = 32'h10408000;
      7430: inst = 32'hc4052ba;
      7431: inst = 32'h8220000;
      7432: inst = 32'h10408000;
      7433: inst = 32'hc4052bb;
      7434: inst = 32'h8220000;
      7435: inst = 32'h10408000;
      7436: inst = 32'hc4052ca;
      7437: inst = 32'h8220000;
      7438: inst = 32'h10408000;
      7439: inst = 32'hc4052cb;
      7440: inst = 32'h8220000;
      7441: inst = 32'h10408000;
      7442: inst = 32'hc4052cc;
      7443: inst = 32'h8220000;
      7444: inst = 32'h10408000;
      7445: inst = 32'hc4052cd;
      7446: inst = 32'h8220000;
      7447: inst = 32'h10408000;
      7448: inst = 32'hc4052ce;
      7449: inst = 32'h8220000;
      7450: inst = 32'h10408000;
      7451: inst = 32'hc4052cf;
      7452: inst = 32'h8220000;
      7453: inst = 32'h10408000;
      7454: inst = 32'hc4052d0;
      7455: inst = 32'h8220000;
      7456: inst = 32'h10408000;
      7457: inst = 32'hc4052d1;
      7458: inst = 32'h8220000;
      7459: inst = 32'h10408000;
      7460: inst = 32'hc4052d2;
      7461: inst = 32'h8220000;
      7462: inst = 32'h10408000;
      7463: inst = 32'hc4052d3;
      7464: inst = 32'h8220000;
      7465: inst = 32'h10408000;
      7466: inst = 32'hc4052d4;
      7467: inst = 32'h8220000;
      7468: inst = 32'h10408000;
      7469: inst = 32'hc4052d5;
      7470: inst = 32'h8220000;
      7471: inst = 32'h10408000;
      7472: inst = 32'hc4052e4;
      7473: inst = 32'h8220000;
      7474: inst = 32'h10408000;
      7475: inst = 32'hc4052e5;
      7476: inst = 32'h8220000;
      7477: inst = 32'h10408000;
      7478: inst = 32'hc4052e6;
      7479: inst = 32'h8220000;
      7480: inst = 32'h10408000;
      7481: inst = 32'hc4052e7;
      7482: inst = 32'h8220000;
      7483: inst = 32'h10408000;
      7484: inst = 32'hc4052e8;
      7485: inst = 32'h8220000;
      7486: inst = 32'h10408000;
      7487: inst = 32'hc4052e9;
      7488: inst = 32'h8220000;
      7489: inst = 32'h10408000;
      7490: inst = 32'hc4052ea;
      7491: inst = 32'h8220000;
      7492: inst = 32'h10408000;
      7493: inst = 32'hc4052eb;
      7494: inst = 32'h8220000;
      7495: inst = 32'h10408000;
      7496: inst = 32'hc4052ec;
      7497: inst = 32'h8220000;
      7498: inst = 32'h10408000;
      7499: inst = 32'hc4052ed;
      7500: inst = 32'h8220000;
      7501: inst = 32'h10408000;
      7502: inst = 32'hc4052ee;
      7503: inst = 32'h8220000;
      7504: inst = 32'hc2094b2;
      7505: inst = 32'h10408000;
      7506: inst = 32'hc403feb;
      7507: inst = 32'h8220000;
      7508: inst = 32'h10408000;
      7509: inst = 32'hc40404b;
      7510: inst = 32'h8220000;
      7511: inst = 32'h10408000;
      7512: inst = 32'hc4040ab;
      7513: inst = 32'h8220000;
      7514: inst = 32'h10408000;
      7515: inst = 32'hc40410b;
      7516: inst = 32'h8220000;
      7517: inst = 32'h10408000;
      7518: inst = 32'hc40416b;
      7519: inst = 32'h8220000;
      7520: inst = 32'h10408000;
      7521: inst = 32'hc4041cb;
      7522: inst = 32'h8220000;
      7523: inst = 32'h10408000;
      7524: inst = 32'hc40422b;
      7525: inst = 32'h8220000;
      7526: inst = 32'h10408000;
      7527: inst = 32'hc40428b;
      7528: inst = 32'h8220000;
      7529: inst = 32'hc20b596;
      7530: inst = 32'h10408000;
      7531: inst = 32'hc4041da;
      7532: inst = 32'h8220000;
      7533: inst = 32'h10408000;
      7534: inst = 32'hc4041db;
      7535: inst = 32'h8220000;
      7536: inst = 32'h10408000;
      7537: inst = 32'hc4041dc;
      7538: inst = 32'h8220000;
      7539: inst = 32'h10408000;
      7540: inst = 32'hc4041dd;
      7541: inst = 32'h8220000;
      7542: inst = 32'h10408000;
      7543: inst = 32'hc4041de;
      7544: inst = 32'h8220000;
      7545: inst = 32'h10408000;
      7546: inst = 32'hc4041df;
      7547: inst = 32'h8220000;
      7548: inst = 32'h10408000;
      7549: inst = 32'hc4041e0;
      7550: inst = 32'h8220000;
      7551: inst = 32'h10408000;
      7552: inst = 32'hc4041e1;
      7553: inst = 32'h8220000;
      7554: inst = 32'h10408000;
      7555: inst = 32'hc4041e2;
      7556: inst = 32'h8220000;
      7557: inst = 32'h10408000;
      7558: inst = 32'hc4041e3;
      7559: inst = 32'h8220000;
      7560: inst = 32'h10408000;
      7561: inst = 32'hc4041e4;
      7562: inst = 32'h8220000;
      7563: inst = 32'h10408000;
      7564: inst = 32'hc4041e5;
      7565: inst = 32'h8220000;
      7566: inst = 32'h10408000;
      7567: inst = 32'hc4041e6;
      7568: inst = 32'h8220000;
      7569: inst = 32'h10408000;
      7570: inst = 32'hc4041e7;
      7571: inst = 32'h8220000;
      7572: inst = 32'h10408000;
      7573: inst = 32'hc4041e8;
      7574: inst = 32'h8220000;
      7575: inst = 32'h10408000;
      7576: inst = 32'hc4041e9;
      7577: inst = 32'h8220000;
      7578: inst = 32'h10408000;
      7579: inst = 32'hc4041ea;
      7580: inst = 32'h8220000;
      7581: inst = 32'h10408000;
      7582: inst = 32'hc4041eb;
      7583: inst = 32'h8220000;
      7584: inst = 32'h10408000;
      7585: inst = 32'hc4041ec;
      7586: inst = 32'h8220000;
      7587: inst = 32'h10408000;
      7588: inst = 32'hc4041ed;
      7589: inst = 32'h8220000;
      7590: inst = 32'h10408000;
      7591: inst = 32'hc4041ee;
      7592: inst = 32'h8220000;
      7593: inst = 32'h10408000;
      7594: inst = 32'hc4041ef;
      7595: inst = 32'h8220000;
      7596: inst = 32'h10408000;
      7597: inst = 32'hc4041f0;
      7598: inst = 32'h8220000;
      7599: inst = 32'h10408000;
      7600: inst = 32'hc4041f1;
      7601: inst = 32'h8220000;
      7602: inst = 32'h10408000;
      7603: inst = 32'hc4041f2;
      7604: inst = 32'h8220000;
      7605: inst = 32'h10408000;
      7606: inst = 32'hc4041f3;
      7607: inst = 32'h8220000;
      7608: inst = 32'h10408000;
      7609: inst = 32'hc4041f4;
      7610: inst = 32'h8220000;
      7611: inst = 32'h10408000;
      7612: inst = 32'hc4041f5;
      7613: inst = 32'h8220000;
      7614: inst = 32'h10408000;
      7615: inst = 32'hc4041f6;
      7616: inst = 32'h8220000;
      7617: inst = 32'h10408000;
      7618: inst = 32'hc4041f7;
      7619: inst = 32'h8220000;
      7620: inst = 32'h10408000;
      7621: inst = 32'hc4041f8;
      7622: inst = 32'h8220000;
      7623: inst = 32'h10408000;
      7624: inst = 32'hc4041f9;
      7625: inst = 32'h8220000;
      7626: inst = 32'h10408000;
      7627: inst = 32'hc4041fa;
      7628: inst = 32'h8220000;
      7629: inst = 32'h10408000;
      7630: inst = 32'hc4041fb;
      7631: inst = 32'h8220000;
      7632: inst = 32'h10408000;
      7633: inst = 32'hc4041fc;
      7634: inst = 32'h8220000;
      7635: inst = 32'h10408000;
      7636: inst = 32'hc4041fd;
      7637: inst = 32'h8220000;
      7638: inst = 32'h10408000;
      7639: inst = 32'hc4041fe;
      7640: inst = 32'h8220000;
      7641: inst = 32'h10408000;
      7642: inst = 32'hc4041ff;
      7643: inst = 32'h8220000;
      7644: inst = 32'h10408000;
      7645: inst = 32'hc404200;
      7646: inst = 32'h8220000;
      7647: inst = 32'h10408000;
      7648: inst = 32'hc404201;
      7649: inst = 32'h8220000;
      7650: inst = 32'h10408000;
      7651: inst = 32'hc404202;
      7652: inst = 32'h8220000;
      7653: inst = 32'h10408000;
      7654: inst = 32'hc404203;
      7655: inst = 32'h8220000;
      7656: inst = 32'h10408000;
      7657: inst = 32'hc404204;
      7658: inst = 32'h8220000;
      7659: inst = 32'h10408000;
      7660: inst = 32'hc404205;
      7661: inst = 32'h8220000;
      7662: inst = 32'h10408000;
      7663: inst = 32'hc404bfa;
      7664: inst = 32'h8220000;
      7665: inst = 32'h10408000;
      7666: inst = 32'hc404bfb;
      7667: inst = 32'h8220000;
      7668: inst = 32'h10408000;
      7669: inst = 32'hc404bfc;
      7670: inst = 32'h8220000;
      7671: inst = 32'h10408000;
      7672: inst = 32'hc404bfd;
      7673: inst = 32'h8220000;
      7674: inst = 32'h10408000;
      7675: inst = 32'hc404bfe;
      7676: inst = 32'h8220000;
      7677: inst = 32'h10408000;
      7678: inst = 32'hc404bff;
      7679: inst = 32'h8220000;
      7680: inst = 32'h10408000;
      7681: inst = 32'hc404c00;
      7682: inst = 32'h8220000;
      7683: inst = 32'h10408000;
      7684: inst = 32'hc404c01;
      7685: inst = 32'h8220000;
      7686: inst = 32'h10408000;
      7687: inst = 32'hc404c02;
      7688: inst = 32'h8220000;
      7689: inst = 32'h10408000;
      7690: inst = 32'hc404c03;
      7691: inst = 32'h8220000;
      7692: inst = 32'h10408000;
      7693: inst = 32'hc404c04;
      7694: inst = 32'h8220000;
      7695: inst = 32'h10408000;
      7696: inst = 32'hc404c05;
      7697: inst = 32'h8220000;
      7698: inst = 32'h10408000;
      7699: inst = 32'hc404c06;
      7700: inst = 32'h8220000;
      7701: inst = 32'h10408000;
      7702: inst = 32'hc404c07;
      7703: inst = 32'h8220000;
      7704: inst = 32'h10408000;
      7705: inst = 32'hc404c08;
      7706: inst = 32'h8220000;
      7707: inst = 32'h10408000;
      7708: inst = 32'hc404c09;
      7709: inst = 32'h8220000;
      7710: inst = 32'h10408000;
      7711: inst = 32'hc404c0a;
      7712: inst = 32'h8220000;
      7713: inst = 32'h10408000;
      7714: inst = 32'hc404c0b;
      7715: inst = 32'h8220000;
      7716: inst = 32'h10408000;
      7717: inst = 32'hc404c0c;
      7718: inst = 32'h8220000;
      7719: inst = 32'h10408000;
      7720: inst = 32'hc404c0d;
      7721: inst = 32'h8220000;
      7722: inst = 32'h10408000;
      7723: inst = 32'hc404c0e;
      7724: inst = 32'h8220000;
      7725: inst = 32'h10408000;
      7726: inst = 32'hc404c0f;
      7727: inst = 32'h8220000;
      7728: inst = 32'h10408000;
      7729: inst = 32'hc404c10;
      7730: inst = 32'h8220000;
      7731: inst = 32'h10408000;
      7732: inst = 32'hc404c11;
      7733: inst = 32'h8220000;
      7734: inst = 32'h10408000;
      7735: inst = 32'hc404c12;
      7736: inst = 32'h8220000;
      7737: inst = 32'h10408000;
      7738: inst = 32'hc404c13;
      7739: inst = 32'h8220000;
      7740: inst = 32'h10408000;
      7741: inst = 32'hc404c14;
      7742: inst = 32'h8220000;
      7743: inst = 32'h10408000;
      7744: inst = 32'hc404c15;
      7745: inst = 32'h8220000;
      7746: inst = 32'h10408000;
      7747: inst = 32'hc404c16;
      7748: inst = 32'h8220000;
      7749: inst = 32'h10408000;
      7750: inst = 32'hc404c17;
      7751: inst = 32'h8220000;
      7752: inst = 32'h10408000;
      7753: inst = 32'hc404c18;
      7754: inst = 32'h8220000;
      7755: inst = 32'h10408000;
      7756: inst = 32'hc404c19;
      7757: inst = 32'h8220000;
      7758: inst = 32'h10408000;
      7759: inst = 32'hc404c1a;
      7760: inst = 32'h8220000;
      7761: inst = 32'h10408000;
      7762: inst = 32'hc404c1b;
      7763: inst = 32'h8220000;
      7764: inst = 32'h10408000;
      7765: inst = 32'hc404c1c;
      7766: inst = 32'h8220000;
      7767: inst = 32'h10408000;
      7768: inst = 32'hc404c1d;
      7769: inst = 32'h8220000;
      7770: inst = 32'h10408000;
      7771: inst = 32'hc404c1e;
      7772: inst = 32'h8220000;
      7773: inst = 32'h10408000;
      7774: inst = 32'hc404c1f;
      7775: inst = 32'h8220000;
      7776: inst = 32'h10408000;
      7777: inst = 32'hc404c20;
      7778: inst = 32'h8220000;
      7779: inst = 32'h10408000;
      7780: inst = 32'hc404c21;
      7781: inst = 32'h8220000;
      7782: inst = 32'h10408000;
      7783: inst = 32'hc404c22;
      7784: inst = 32'h8220000;
      7785: inst = 32'h10408000;
      7786: inst = 32'hc404c23;
      7787: inst = 32'h8220000;
      7788: inst = 32'h10408000;
      7789: inst = 32'hc404c24;
      7790: inst = 32'h8220000;
      7791: inst = 32'h10408000;
      7792: inst = 32'hc404c25;
      7793: inst = 32'h8220000;
      7794: inst = 32'hc20ffff;
      7795: inst = 32'h10408000;
      7796: inst = 32'hc40423c;
      7797: inst = 32'h8220000;
      7798: inst = 32'h10408000;
      7799: inst = 32'hc40423d;
      7800: inst = 32'h8220000;
      7801: inst = 32'h10408000;
      7802: inst = 32'hc40423e;
      7803: inst = 32'h8220000;
      7804: inst = 32'h10408000;
      7805: inst = 32'hc40423f;
      7806: inst = 32'h8220000;
      7807: inst = 32'h10408000;
      7808: inst = 32'hc404240;
      7809: inst = 32'h8220000;
      7810: inst = 32'h10408000;
      7811: inst = 32'hc404241;
      7812: inst = 32'h8220000;
      7813: inst = 32'h10408000;
      7814: inst = 32'hc404242;
      7815: inst = 32'h8220000;
      7816: inst = 32'h10408000;
      7817: inst = 32'hc404243;
      7818: inst = 32'h8220000;
      7819: inst = 32'h10408000;
      7820: inst = 32'hc404244;
      7821: inst = 32'h8220000;
      7822: inst = 32'h10408000;
      7823: inst = 32'hc404245;
      7824: inst = 32'h8220000;
      7825: inst = 32'h10408000;
      7826: inst = 32'hc404246;
      7827: inst = 32'h8220000;
      7828: inst = 32'h10408000;
      7829: inst = 32'hc404247;
      7830: inst = 32'h8220000;
      7831: inst = 32'h10408000;
      7832: inst = 32'hc404248;
      7833: inst = 32'h8220000;
      7834: inst = 32'h10408000;
      7835: inst = 32'hc404249;
      7836: inst = 32'h8220000;
      7837: inst = 32'h10408000;
      7838: inst = 32'hc40424a;
      7839: inst = 32'h8220000;
      7840: inst = 32'h10408000;
      7841: inst = 32'hc40424b;
      7842: inst = 32'h8220000;
      7843: inst = 32'h10408000;
      7844: inst = 32'hc40424c;
      7845: inst = 32'h8220000;
      7846: inst = 32'h10408000;
      7847: inst = 32'hc40424d;
      7848: inst = 32'h8220000;
      7849: inst = 32'h10408000;
      7850: inst = 32'hc40424e;
      7851: inst = 32'h8220000;
      7852: inst = 32'h10408000;
      7853: inst = 32'hc40424f;
      7854: inst = 32'h8220000;
      7855: inst = 32'h10408000;
      7856: inst = 32'hc404250;
      7857: inst = 32'h8220000;
      7858: inst = 32'h10408000;
      7859: inst = 32'hc404251;
      7860: inst = 32'h8220000;
      7861: inst = 32'h10408000;
      7862: inst = 32'hc404252;
      7863: inst = 32'h8220000;
      7864: inst = 32'h10408000;
      7865: inst = 32'hc404253;
      7866: inst = 32'h8220000;
      7867: inst = 32'h10408000;
      7868: inst = 32'hc404254;
      7869: inst = 32'h8220000;
      7870: inst = 32'h10408000;
      7871: inst = 32'hc404255;
      7872: inst = 32'h8220000;
      7873: inst = 32'h10408000;
      7874: inst = 32'hc404256;
      7875: inst = 32'h8220000;
      7876: inst = 32'h10408000;
      7877: inst = 32'hc404257;
      7878: inst = 32'h8220000;
      7879: inst = 32'h10408000;
      7880: inst = 32'hc404258;
      7881: inst = 32'h8220000;
      7882: inst = 32'h10408000;
      7883: inst = 32'hc404259;
      7884: inst = 32'h8220000;
      7885: inst = 32'h10408000;
      7886: inst = 32'hc40425a;
      7887: inst = 32'h8220000;
      7888: inst = 32'h10408000;
      7889: inst = 32'hc40425b;
      7890: inst = 32'h8220000;
      7891: inst = 32'h10408000;
      7892: inst = 32'hc40425c;
      7893: inst = 32'h8220000;
      7894: inst = 32'h10408000;
      7895: inst = 32'hc40425d;
      7896: inst = 32'h8220000;
      7897: inst = 32'h10408000;
      7898: inst = 32'hc40425e;
      7899: inst = 32'h8220000;
      7900: inst = 32'h10408000;
      7901: inst = 32'hc40425f;
      7902: inst = 32'h8220000;
      7903: inst = 32'h10408000;
      7904: inst = 32'hc404260;
      7905: inst = 32'h8220000;
      7906: inst = 32'h10408000;
      7907: inst = 32'hc404261;
      7908: inst = 32'h8220000;
      7909: inst = 32'h10408000;
      7910: inst = 32'hc404262;
      7911: inst = 32'h8220000;
      7912: inst = 32'h10408000;
      7913: inst = 32'hc404263;
      7914: inst = 32'h8220000;
      7915: inst = 32'h10408000;
      7916: inst = 32'hc40429c;
      7917: inst = 32'h8220000;
      7918: inst = 32'h10408000;
      7919: inst = 32'hc40429d;
      7920: inst = 32'h8220000;
      7921: inst = 32'h10408000;
      7922: inst = 32'hc40429e;
      7923: inst = 32'h8220000;
      7924: inst = 32'h10408000;
      7925: inst = 32'hc40429f;
      7926: inst = 32'h8220000;
      7927: inst = 32'h10408000;
      7928: inst = 32'hc4042a0;
      7929: inst = 32'h8220000;
      7930: inst = 32'h10408000;
      7931: inst = 32'hc4042a1;
      7932: inst = 32'h8220000;
      7933: inst = 32'h10408000;
      7934: inst = 32'hc4042a2;
      7935: inst = 32'h8220000;
      7936: inst = 32'h10408000;
      7937: inst = 32'hc4042a3;
      7938: inst = 32'h8220000;
      7939: inst = 32'h10408000;
      7940: inst = 32'hc4042a4;
      7941: inst = 32'h8220000;
      7942: inst = 32'h10408000;
      7943: inst = 32'hc4042a5;
      7944: inst = 32'h8220000;
      7945: inst = 32'h10408000;
      7946: inst = 32'hc4042a6;
      7947: inst = 32'h8220000;
      7948: inst = 32'h10408000;
      7949: inst = 32'hc4042a7;
      7950: inst = 32'h8220000;
      7951: inst = 32'h10408000;
      7952: inst = 32'hc4042a8;
      7953: inst = 32'h8220000;
      7954: inst = 32'h10408000;
      7955: inst = 32'hc4042a9;
      7956: inst = 32'h8220000;
      7957: inst = 32'h10408000;
      7958: inst = 32'hc4042aa;
      7959: inst = 32'h8220000;
      7960: inst = 32'h10408000;
      7961: inst = 32'hc4042ab;
      7962: inst = 32'h8220000;
      7963: inst = 32'h10408000;
      7964: inst = 32'hc4042ac;
      7965: inst = 32'h8220000;
      7966: inst = 32'h10408000;
      7967: inst = 32'hc4042ad;
      7968: inst = 32'h8220000;
      7969: inst = 32'h10408000;
      7970: inst = 32'hc4042ae;
      7971: inst = 32'h8220000;
      7972: inst = 32'h10408000;
      7973: inst = 32'hc4042af;
      7974: inst = 32'h8220000;
      7975: inst = 32'h10408000;
      7976: inst = 32'hc4042b0;
      7977: inst = 32'h8220000;
      7978: inst = 32'h10408000;
      7979: inst = 32'hc4042b1;
      7980: inst = 32'h8220000;
      7981: inst = 32'h10408000;
      7982: inst = 32'hc4042b2;
      7983: inst = 32'h8220000;
      7984: inst = 32'h10408000;
      7985: inst = 32'hc4042b3;
      7986: inst = 32'h8220000;
      7987: inst = 32'h10408000;
      7988: inst = 32'hc4042b4;
      7989: inst = 32'h8220000;
      7990: inst = 32'h10408000;
      7991: inst = 32'hc4042b5;
      7992: inst = 32'h8220000;
      7993: inst = 32'h10408000;
      7994: inst = 32'hc4042b6;
      7995: inst = 32'h8220000;
      7996: inst = 32'h10408000;
      7997: inst = 32'hc4042b7;
      7998: inst = 32'h8220000;
      7999: inst = 32'h10408000;
      8000: inst = 32'hc4042b8;
      8001: inst = 32'h8220000;
      8002: inst = 32'h10408000;
      8003: inst = 32'hc4042b9;
      8004: inst = 32'h8220000;
      8005: inst = 32'h10408000;
      8006: inst = 32'hc4042ba;
      8007: inst = 32'h8220000;
      8008: inst = 32'h10408000;
      8009: inst = 32'hc4042bb;
      8010: inst = 32'h8220000;
      8011: inst = 32'h10408000;
      8012: inst = 32'hc4042bc;
      8013: inst = 32'h8220000;
      8014: inst = 32'h10408000;
      8015: inst = 32'hc4042bd;
      8016: inst = 32'h8220000;
      8017: inst = 32'h10408000;
      8018: inst = 32'hc4042be;
      8019: inst = 32'h8220000;
      8020: inst = 32'h10408000;
      8021: inst = 32'hc4042bf;
      8022: inst = 32'h8220000;
      8023: inst = 32'h10408000;
      8024: inst = 32'hc4042c0;
      8025: inst = 32'h8220000;
      8026: inst = 32'h10408000;
      8027: inst = 32'hc4042c1;
      8028: inst = 32'h8220000;
      8029: inst = 32'h10408000;
      8030: inst = 32'hc4042c2;
      8031: inst = 32'h8220000;
      8032: inst = 32'h10408000;
      8033: inst = 32'hc4042c3;
      8034: inst = 32'h8220000;
      8035: inst = 32'h10408000;
      8036: inst = 32'hc4042fc;
      8037: inst = 32'h8220000;
      8038: inst = 32'h10408000;
      8039: inst = 32'hc4042fd;
      8040: inst = 32'h8220000;
      8041: inst = 32'h10408000;
      8042: inst = 32'hc4042fe;
      8043: inst = 32'h8220000;
      8044: inst = 32'h10408000;
      8045: inst = 32'hc4042ff;
      8046: inst = 32'h8220000;
      8047: inst = 32'h10408000;
      8048: inst = 32'hc404300;
      8049: inst = 32'h8220000;
      8050: inst = 32'h10408000;
      8051: inst = 32'hc404301;
      8052: inst = 32'h8220000;
      8053: inst = 32'h10408000;
      8054: inst = 32'hc404302;
      8055: inst = 32'h8220000;
      8056: inst = 32'h10408000;
      8057: inst = 32'hc404303;
      8058: inst = 32'h8220000;
      8059: inst = 32'h10408000;
      8060: inst = 32'hc404304;
      8061: inst = 32'h8220000;
      8062: inst = 32'h10408000;
      8063: inst = 32'hc404305;
      8064: inst = 32'h8220000;
      8065: inst = 32'h10408000;
      8066: inst = 32'hc404306;
      8067: inst = 32'h8220000;
      8068: inst = 32'h10408000;
      8069: inst = 32'hc404307;
      8070: inst = 32'h8220000;
      8071: inst = 32'h10408000;
      8072: inst = 32'hc404308;
      8073: inst = 32'h8220000;
      8074: inst = 32'h10408000;
      8075: inst = 32'hc404309;
      8076: inst = 32'h8220000;
      8077: inst = 32'h10408000;
      8078: inst = 32'hc40430a;
      8079: inst = 32'h8220000;
      8080: inst = 32'h10408000;
      8081: inst = 32'hc40430b;
      8082: inst = 32'h8220000;
      8083: inst = 32'h10408000;
      8084: inst = 32'hc40430c;
      8085: inst = 32'h8220000;
      8086: inst = 32'h10408000;
      8087: inst = 32'hc40430d;
      8088: inst = 32'h8220000;
      8089: inst = 32'h10408000;
      8090: inst = 32'hc40430e;
      8091: inst = 32'h8220000;
      8092: inst = 32'h10408000;
      8093: inst = 32'hc40430f;
      8094: inst = 32'h8220000;
      8095: inst = 32'h10408000;
      8096: inst = 32'hc404310;
      8097: inst = 32'h8220000;
      8098: inst = 32'h10408000;
      8099: inst = 32'hc404311;
      8100: inst = 32'h8220000;
      8101: inst = 32'h10408000;
      8102: inst = 32'hc404312;
      8103: inst = 32'h8220000;
      8104: inst = 32'h10408000;
      8105: inst = 32'hc404313;
      8106: inst = 32'h8220000;
      8107: inst = 32'h10408000;
      8108: inst = 32'hc404314;
      8109: inst = 32'h8220000;
      8110: inst = 32'h10408000;
      8111: inst = 32'hc404315;
      8112: inst = 32'h8220000;
      8113: inst = 32'h10408000;
      8114: inst = 32'hc404316;
      8115: inst = 32'h8220000;
      8116: inst = 32'h10408000;
      8117: inst = 32'hc404317;
      8118: inst = 32'h8220000;
      8119: inst = 32'h10408000;
      8120: inst = 32'hc404318;
      8121: inst = 32'h8220000;
      8122: inst = 32'h10408000;
      8123: inst = 32'hc404319;
      8124: inst = 32'h8220000;
      8125: inst = 32'h10408000;
      8126: inst = 32'hc40431a;
      8127: inst = 32'h8220000;
      8128: inst = 32'h10408000;
      8129: inst = 32'hc40431b;
      8130: inst = 32'h8220000;
      8131: inst = 32'h10408000;
      8132: inst = 32'hc40431c;
      8133: inst = 32'h8220000;
      8134: inst = 32'h10408000;
      8135: inst = 32'hc40431d;
      8136: inst = 32'h8220000;
      8137: inst = 32'h10408000;
      8138: inst = 32'hc40431e;
      8139: inst = 32'h8220000;
      8140: inst = 32'h10408000;
      8141: inst = 32'hc40431f;
      8142: inst = 32'h8220000;
      8143: inst = 32'h10408000;
      8144: inst = 32'hc404320;
      8145: inst = 32'h8220000;
      8146: inst = 32'h10408000;
      8147: inst = 32'hc404321;
      8148: inst = 32'h8220000;
      8149: inst = 32'h10408000;
      8150: inst = 32'hc404322;
      8151: inst = 32'h8220000;
      8152: inst = 32'h10408000;
      8153: inst = 32'hc404323;
      8154: inst = 32'h8220000;
      8155: inst = 32'h10408000;
      8156: inst = 32'hc40435c;
      8157: inst = 32'h8220000;
      8158: inst = 32'h10408000;
      8159: inst = 32'hc40435d;
      8160: inst = 32'h8220000;
      8161: inst = 32'h10408000;
      8162: inst = 32'hc40435e;
      8163: inst = 32'h8220000;
      8164: inst = 32'h10408000;
      8165: inst = 32'hc40435f;
      8166: inst = 32'h8220000;
      8167: inst = 32'h10408000;
      8168: inst = 32'hc404360;
      8169: inst = 32'h8220000;
      8170: inst = 32'h10408000;
      8171: inst = 32'hc404361;
      8172: inst = 32'h8220000;
      8173: inst = 32'h10408000;
      8174: inst = 32'hc404362;
      8175: inst = 32'h8220000;
      8176: inst = 32'h10408000;
      8177: inst = 32'hc404363;
      8178: inst = 32'h8220000;
      8179: inst = 32'h10408000;
      8180: inst = 32'hc404364;
      8181: inst = 32'h8220000;
      8182: inst = 32'h10408000;
      8183: inst = 32'hc404365;
      8184: inst = 32'h8220000;
      8185: inst = 32'h10408000;
      8186: inst = 32'hc404366;
      8187: inst = 32'h8220000;
      8188: inst = 32'h10408000;
      8189: inst = 32'hc404367;
      8190: inst = 32'h8220000;
      8191: inst = 32'h10408000;
      8192: inst = 32'hc404368;
      8193: inst = 32'h8220000;
      8194: inst = 32'h10408000;
      8195: inst = 32'hc404369;
      8196: inst = 32'h8220000;
      8197: inst = 32'h10408000;
      8198: inst = 32'hc40436a;
      8199: inst = 32'h8220000;
      8200: inst = 32'h10408000;
      8201: inst = 32'hc40436b;
      8202: inst = 32'h8220000;
      8203: inst = 32'h10408000;
      8204: inst = 32'hc40436c;
      8205: inst = 32'h8220000;
      8206: inst = 32'h10408000;
      8207: inst = 32'hc40436d;
      8208: inst = 32'h8220000;
      8209: inst = 32'h10408000;
      8210: inst = 32'hc40436e;
      8211: inst = 32'h8220000;
      8212: inst = 32'h10408000;
      8213: inst = 32'hc40436f;
      8214: inst = 32'h8220000;
      8215: inst = 32'h10408000;
      8216: inst = 32'hc404370;
      8217: inst = 32'h8220000;
      8218: inst = 32'h10408000;
      8219: inst = 32'hc404371;
      8220: inst = 32'h8220000;
      8221: inst = 32'h10408000;
      8222: inst = 32'hc404372;
      8223: inst = 32'h8220000;
      8224: inst = 32'h10408000;
      8225: inst = 32'hc404373;
      8226: inst = 32'h8220000;
      8227: inst = 32'h10408000;
      8228: inst = 32'hc404374;
      8229: inst = 32'h8220000;
      8230: inst = 32'h10408000;
      8231: inst = 32'hc404375;
      8232: inst = 32'h8220000;
      8233: inst = 32'h10408000;
      8234: inst = 32'hc404376;
      8235: inst = 32'h8220000;
      8236: inst = 32'h10408000;
      8237: inst = 32'hc404377;
      8238: inst = 32'h8220000;
      8239: inst = 32'h10408000;
      8240: inst = 32'hc404378;
      8241: inst = 32'h8220000;
      8242: inst = 32'h10408000;
      8243: inst = 32'hc404379;
      8244: inst = 32'h8220000;
      8245: inst = 32'h10408000;
      8246: inst = 32'hc40437a;
      8247: inst = 32'h8220000;
      8248: inst = 32'h10408000;
      8249: inst = 32'hc40437b;
      8250: inst = 32'h8220000;
      8251: inst = 32'h10408000;
      8252: inst = 32'hc40437c;
      8253: inst = 32'h8220000;
      8254: inst = 32'h10408000;
      8255: inst = 32'hc40437d;
      8256: inst = 32'h8220000;
      8257: inst = 32'h10408000;
      8258: inst = 32'hc40437e;
      8259: inst = 32'h8220000;
      8260: inst = 32'h10408000;
      8261: inst = 32'hc40437f;
      8262: inst = 32'h8220000;
      8263: inst = 32'h10408000;
      8264: inst = 32'hc404380;
      8265: inst = 32'h8220000;
      8266: inst = 32'h10408000;
      8267: inst = 32'hc404381;
      8268: inst = 32'h8220000;
      8269: inst = 32'h10408000;
      8270: inst = 32'hc404382;
      8271: inst = 32'h8220000;
      8272: inst = 32'h10408000;
      8273: inst = 32'hc404383;
      8274: inst = 32'h8220000;
      8275: inst = 32'h10408000;
      8276: inst = 32'hc4043bc;
      8277: inst = 32'h8220000;
      8278: inst = 32'h10408000;
      8279: inst = 32'hc4043bd;
      8280: inst = 32'h8220000;
      8281: inst = 32'h10408000;
      8282: inst = 32'hc4043be;
      8283: inst = 32'h8220000;
      8284: inst = 32'h10408000;
      8285: inst = 32'hc4043bf;
      8286: inst = 32'h8220000;
      8287: inst = 32'h10408000;
      8288: inst = 32'hc4043c0;
      8289: inst = 32'h8220000;
      8290: inst = 32'h10408000;
      8291: inst = 32'hc4043c1;
      8292: inst = 32'h8220000;
      8293: inst = 32'h10408000;
      8294: inst = 32'hc4043c2;
      8295: inst = 32'h8220000;
      8296: inst = 32'h10408000;
      8297: inst = 32'hc4043c3;
      8298: inst = 32'h8220000;
      8299: inst = 32'h10408000;
      8300: inst = 32'hc4043c4;
      8301: inst = 32'h8220000;
      8302: inst = 32'h10408000;
      8303: inst = 32'hc4043c5;
      8304: inst = 32'h8220000;
      8305: inst = 32'h10408000;
      8306: inst = 32'hc4043c6;
      8307: inst = 32'h8220000;
      8308: inst = 32'h10408000;
      8309: inst = 32'hc4043c7;
      8310: inst = 32'h8220000;
      8311: inst = 32'h10408000;
      8312: inst = 32'hc4043c8;
      8313: inst = 32'h8220000;
      8314: inst = 32'h10408000;
      8315: inst = 32'hc4043c9;
      8316: inst = 32'h8220000;
      8317: inst = 32'h10408000;
      8318: inst = 32'hc4043ca;
      8319: inst = 32'h8220000;
      8320: inst = 32'h10408000;
      8321: inst = 32'hc4043cb;
      8322: inst = 32'h8220000;
      8323: inst = 32'h10408000;
      8324: inst = 32'hc4043cc;
      8325: inst = 32'h8220000;
      8326: inst = 32'h10408000;
      8327: inst = 32'hc4043cd;
      8328: inst = 32'h8220000;
      8329: inst = 32'h10408000;
      8330: inst = 32'hc4043ce;
      8331: inst = 32'h8220000;
      8332: inst = 32'h10408000;
      8333: inst = 32'hc4043cf;
      8334: inst = 32'h8220000;
      8335: inst = 32'h10408000;
      8336: inst = 32'hc4043d0;
      8337: inst = 32'h8220000;
      8338: inst = 32'h10408000;
      8339: inst = 32'hc4043d1;
      8340: inst = 32'h8220000;
      8341: inst = 32'h10408000;
      8342: inst = 32'hc4043d2;
      8343: inst = 32'h8220000;
      8344: inst = 32'h10408000;
      8345: inst = 32'hc4043d3;
      8346: inst = 32'h8220000;
      8347: inst = 32'h10408000;
      8348: inst = 32'hc4043d4;
      8349: inst = 32'h8220000;
      8350: inst = 32'h10408000;
      8351: inst = 32'hc4043d5;
      8352: inst = 32'h8220000;
      8353: inst = 32'h10408000;
      8354: inst = 32'hc4043d6;
      8355: inst = 32'h8220000;
      8356: inst = 32'h10408000;
      8357: inst = 32'hc4043d7;
      8358: inst = 32'h8220000;
      8359: inst = 32'h10408000;
      8360: inst = 32'hc4043d8;
      8361: inst = 32'h8220000;
      8362: inst = 32'h10408000;
      8363: inst = 32'hc4043d9;
      8364: inst = 32'h8220000;
      8365: inst = 32'h10408000;
      8366: inst = 32'hc4043da;
      8367: inst = 32'h8220000;
      8368: inst = 32'h10408000;
      8369: inst = 32'hc4043db;
      8370: inst = 32'h8220000;
      8371: inst = 32'h10408000;
      8372: inst = 32'hc4043dc;
      8373: inst = 32'h8220000;
      8374: inst = 32'h10408000;
      8375: inst = 32'hc4043dd;
      8376: inst = 32'h8220000;
      8377: inst = 32'h10408000;
      8378: inst = 32'hc4043de;
      8379: inst = 32'h8220000;
      8380: inst = 32'h10408000;
      8381: inst = 32'hc4043df;
      8382: inst = 32'h8220000;
      8383: inst = 32'h10408000;
      8384: inst = 32'hc4043e0;
      8385: inst = 32'h8220000;
      8386: inst = 32'h10408000;
      8387: inst = 32'hc4043e1;
      8388: inst = 32'h8220000;
      8389: inst = 32'h10408000;
      8390: inst = 32'hc4043e2;
      8391: inst = 32'h8220000;
      8392: inst = 32'h10408000;
      8393: inst = 32'hc4043e3;
      8394: inst = 32'h8220000;
      8395: inst = 32'h10408000;
      8396: inst = 32'hc40441c;
      8397: inst = 32'h8220000;
      8398: inst = 32'h10408000;
      8399: inst = 32'hc40441d;
      8400: inst = 32'h8220000;
      8401: inst = 32'h10408000;
      8402: inst = 32'hc40441e;
      8403: inst = 32'h8220000;
      8404: inst = 32'h10408000;
      8405: inst = 32'hc40441f;
      8406: inst = 32'h8220000;
      8407: inst = 32'h10408000;
      8408: inst = 32'hc404420;
      8409: inst = 32'h8220000;
      8410: inst = 32'h10408000;
      8411: inst = 32'hc404421;
      8412: inst = 32'h8220000;
      8413: inst = 32'h10408000;
      8414: inst = 32'hc404422;
      8415: inst = 32'h8220000;
      8416: inst = 32'h10408000;
      8417: inst = 32'hc404423;
      8418: inst = 32'h8220000;
      8419: inst = 32'h10408000;
      8420: inst = 32'hc404424;
      8421: inst = 32'h8220000;
      8422: inst = 32'h10408000;
      8423: inst = 32'hc404425;
      8424: inst = 32'h8220000;
      8425: inst = 32'h10408000;
      8426: inst = 32'hc404426;
      8427: inst = 32'h8220000;
      8428: inst = 32'h10408000;
      8429: inst = 32'hc404427;
      8430: inst = 32'h8220000;
      8431: inst = 32'h10408000;
      8432: inst = 32'hc404428;
      8433: inst = 32'h8220000;
      8434: inst = 32'h10408000;
      8435: inst = 32'hc404429;
      8436: inst = 32'h8220000;
      8437: inst = 32'h10408000;
      8438: inst = 32'hc40442a;
      8439: inst = 32'h8220000;
      8440: inst = 32'h10408000;
      8441: inst = 32'hc40442b;
      8442: inst = 32'h8220000;
      8443: inst = 32'h10408000;
      8444: inst = 32'hc40442c;
      8445: inst = 32'h8220000;
      8446: inst = 32'h10408000;
      8447: inst = 32'hc40442d;
      8448: inst = 32'h8220000;
      8449: inst = 32'h10408000;
      8450: inst = 32'hc40442e;
      8451: inst = 32'h8220000;
      8452: inst = 32'h10408000;
      8453: inst = 32'hc40442f;
      8454: inst = 32'h8220000;
      8455: inst = 32'h10408000;
      8456: inst = 32'hc404430;
      8457: inst = 32'h8220000;
      8458: inst = 32'h10408000;
      8459: inst = 32'hc404431;
      8460: inst = 32'h8220000;
      8461: inst = 32'h10408000;
      8462: inst = 32'hc404432;
      8463: inst = 32'h8220000;
      8464: inst = 32'h10408000;
      8465: inst = 32'hc404433;
      8466: inst = 32'h8220000;
      8467: inst = 32'h10408000;
      8468: inst = 32'hc404434;
      8469: inst = 32'h8220000;
      8470: inst = 32'h10408000;
      8471: inst = 32'hc404435;
      8472: inst = 32'h8220000;
      8473: inst = 32'h10408000;
      8474: inst = 32'hc404436;
      8475: inst = 32'h8220000;
      8476: inst = 32'h10408000;
      8477: inst = 32'hc404437;
      8478: inst = 32'h8220000;
      8479: inst = 32'h10408000;
      8480: inst = 32'hc404438;
      8481: inst = 32'h8220000;
      8482: inst = 32'h10408000;
      8483: inst = 32'hc404439;
      8484: inst = 32'h8220000;
      8485: inst = 32'h10408000;
      8486: inst = 32'hc40443a;
      8487: inst = 32'h8220000;
      8488: inst = 32'h10408000;
      8489: inst = 32'hc40443b;
      8490: inst = 32'h8220000;
      8491: inst = 32'h10408000;
      8492: inst = 32'hc40443c;
      8493: inst = 32'h8220000;
      8494: inst = 32'h10408000;
      8495: inst = 32'hc40443d;
      8496: inst = 32'h8220000;
      8497: inst = 32'h10408000;
      8498: inst = 32'hc40443e;
      8499: inst = 32'h8220000;
      8500: inst = 32'h10408000;
      8501: inst = 32'hc40443f;
      8502: inst = 32'h8220000;
      8503: inst = 32'h10408000;
      8504: inst = 32'hc404440;
      8505: inst = 32'h8220000;
      8506: inst = 32'h10408000;
      8507: inst = 32'hc404441;
      8508: inst = 32'h8220000;
      8509: inst = 32'h10408000;
      8510: inst = 32'hc404442;
      8511: inst = 32'h8220000;
      8512: inst = 32'h10408000;
      8513: inst = 32'hc404443;
      8514: inst = 32'h8220000;
      8515: inst = 32'h10408000;
      8516: inst = 32'hc40447c;
      8517: inst = 32'h8220000;
      8518: inst = 32'h10408000;
      8519: inst = 32'hc40447d;
      8520: inst = 32'h8220000;
      8521: inst = 32'h10408000;
      8522: inst = 32'hc40447e;
      8523: inst = 32'h8220000;
      8524: inst = 32'h10408000;
      8525: inst = 32'hc40447f;
      8526: inst = 32'h8220000;
      8527: inst = 32'h10408000;
      8528: inst = 32'hc404480;
      8529: inst = 32'h8220000;
      8530: inst = 32'h10408000;
      8531: inst = 32'hc404481;
      8532: inst = 32'h8220000;
      8533: inst = 32'h10408000;
      8534: inst = 32'hc404482;
      8535: inst = 32'h8220000;
      8536: inst = 32'h10408000;
      8537: inst = 32'hc404483;
      8538: inst = 32'h8220000;
      8539: inst = 32'h10408000;
      8540: inst = 32'hc404484;
      8541: inst = 32'h8220000;
      8542: inst = 32'h10408000;
      8543: inst = 32'hc404485;
      8544: inst = 32'h8220000;
      8545: inst = 32'h10408000;
      8546: inst = 32'hc404486;
      8547: inst = 32'h8220000;
      8548: inst = 32'h10408000;
      8549: inst = 32'hc404487;
      8550: inst = 32'h8220000;
      8551: inst = 32'h10408000;
      8552: inst = 32'hc404488;
      8553: inst = 32'h8220000;
      8554: inst = 32'h10408000;
      8555: inst = 32'hc404489;
      8556: inst = 32'h8220000;
      8557: inst = 32'h10408000;
      8558: inst = 32'hc40448a;
      8559: inst = 32'h8220000;
      8560: inst = 32'h10408000;
      8561: inst = 32'hc40448b;
      8562: inst = 32'h8220000;
      8563: inst = 32'h10408000;
      8564: inst = 32'hc40448c;
      8565: inst = 32'h8220000;
      8566: inst = 32'h10408000;
      8567: inst = 32'hc40448d;
      8568: inst = 32'h8220000;
      8569: inst = 32'h10408000;
      8570: inst = 32'hc40448e;
      8571: inst = 32'h8220000;
      8572: inst = 32'h10408000;
      8573: inst = 32'hc40448f;
      8574: inst = 32'h8220000;
      8575: inst = 32'h10408000;
      8576: inst = 32'hc404490;
      8577: inst = 32'h8220000;
      8578: inst = 32'h10408000;
      8579: inst = 32'hc404491;
      8580: inst = 32'h8220000;
      8581: inst = 32'h10408000;
      8582: inst = 32'hc404492;
      8583: inst = 32'h8220000;
      8584: inst = 32'h10408000;
      8585: inst = 32'hc404493;
      8586: inst = 32'h8220000;
      8587: inst = 32'h10408000;
      8588: inst = 32'hc404494;
      8589: inst = 32'h8220000;
      8590: inst = 32'h10408000;
      8591: inst = 32'hc404495;
      8592: inst = 32'h8220000;
      8593: inst = 32'h10408000;
      8594: inst = 32'hc404496;
      8595: inst = 32'h8220000;
      8596: inst = 32'h10408000;
      8597: inst = 32'hc404497;
      8598: inst = 32'h8220000;
      8599: inst = 32'h10408000;
      8600: inst = 32'hc404498;
      8601: inst = 32'h8220000;
      8602: inst = 32'h10408000;
      8603: inst = 32'hc404499;
      8604: inst = 32'h8220000;
      8605: inst = 32'h10408000;
      8606: inst = 32'hc40449a;
      8607: inst = 32'h8220000;
      8608: inst = 32'h10408000;
      8609: inst = 32'hc40449b;
      8610: inst = 32'h8220000;
      8611: inst = 32'h10408000;
      8612: inst = 32'hc40449c;
      8613: inst = 32'h8220000;
      8614: inst = 32'h10408000;
      8615: inst = 32'hc40449d;
      8616: inst = 32'h8220000;
      8617: inst = 32'h10408000;
      8618: inst = 32'hc40449e;
      8619: inst = 32'h8220000;
      8620: inst = 32'h10408000;
      8621: inst = 32'hc40449f;
      8622: inst = 32'h8220000;
      8623: inst = 32'h10408000;
      8624: inst = 32'hc4044a0;
      8625: inst = 32'h8220000;
      8626: inst = 32'h10408000;
      8627: inst = 32'hc4044a1;
      8628: inst = 32'h8220000;
      8629: inst = 32'h10408000;
      8630: inst = 32'hc4044a2;
      8631: inst = 32'h8220000;
      8632: inst = 32'h10408000;
      8633: inst = 32'hc4044a3;
      8634: inst = 32'h8220000;
      8635: inst = 32'h10408000;
      8636: inst = 32'hc4044dc;
      8637: inst = 32'h8220000;
      8638: inst = 32'h10408000;
      8639: inst = 32'hc4044dd;
      8640: inst = 32'h8220000;
      8641: inst = 32'h10408000;
      8642: inst = 32'hc4044de;
      8643: inst = 32'h8220000;
      8644: inst = 32'h10408000;
      8645: inst = 32'hc4044df;
      8646: inst = 32'h8220000;
      8647: inst = 32'h10408000;
      8648: inst = 32'hc4044e0;
      8649: inst = 32'h8220000;
      8650: inst = 32'h10408000;
      8651: inst = 32'hc4044e1;
      8652: inst = 32'h8220000;
      8653: inst = 32'h10408000;
      8654: inst = 32'hc4044e2;
      8655: inst = 32'h8220000;
      8656: inst = 32'h10408000;
      8657: inst = 32'hc4044e3;
      8658: inst = 32'h8220000;
      8659: inst = 32'h10408000;
      8660: inst = 32'hc4044e4;
      8661: inst = 32'h8220000;
      8662: inst = 32'h10408000;
      8663: inst = 32'hc4044e5;
      8664: inst = 32'h8220000;
      8665: inst = 32'h10408000;
      8666: inst = 32'hc4044e6;
      8667: inst = 32'h8220000;
      8668: inst = 32'h10408000;
      8669: inst = 32'hc4044e7;
      8670: inst = 32'h8220000;
      8671: inst = 32'h10408000;
      8672: inst = 32'hc4044e8;
      8673: inst = 32'h8220000;
      8674: inst = 32'h10408000;
      8675: inst = 32'hc4044e9;
      8676: inst = 32'h8220000;
      8677: inst = 32'h10408000;
      8678: inst = 32'hc4044ea;
      8679: inst = 32'h8220000;
      8680: inst = 32'h10408000;
      8681: inst = 32'hc4044eb;
      8682: inst = 32'h8220000;
      8683: inst = 32'h10408000;
      8684: inst = 32'hc4044ec;
      8685: inst = 32'h8220000;
      8686: inst = 32'h10408000;
      8687: inst = 32'hc4044ed;
      8688: inst = 32'h8220000;
      8689: inst = 32'h10408000;
      8690: inst = 32'hc4044ee;
      8691: inst = 32'h8220000;
      8692: inst = 32'h10408000;
      8693: inst = 32'hc4044ef;
      8694: inst = 32'h8220000;
      8695: inst = 32'h10408000;
      8696: inst = 32'hc4044f0;
      8697: inst = 32'h8220000;
      8698: inst = 32'h10408000;
      8699: inst = 32'hc4044f1;
      8700: inst = 32'h8220000;
      8701: inst = 32'h10408000;
      8702: inst = 32'hc4044f2;
      8703: inst = 32'h8220000;
      8704: inst = 32'h10408000;
      8705: inst = 32'hc4044f3;
      8706: inst = 32'h8220000;
      8707: inst = 32'h10408000;
      8708: inst = 32'hc4044f4;
      8709: inst = 32'h8220000;
      8710: inst = 32'h10408000;
      8711: inst = 32'hc4044f5;
      8712: inst = 32'h8220000;
      8713: inst = 32'h10408000;
      8714: inst = 32'hc4044f6;
      8715: inst = 32'h8220000;
      8716: inst = 32'h10408000;
      8717: inst = 32'hc4044f7;
      8718: inst = 32'h8220000;
      8719: inst = 32'h10408000;
      8720: inst = 32'hc4044f8;
      8721: inst = 32'h8220000;
      8722: inst = 32'h10408000;
      8723: inst = 32'hc4044f9;
      8724: inst = 32'h8220000;
      8725: inst = 32'h10408000;
      8726: inst = 32'hc4044fa;
      8727: inst = 32'h8220000;
      8728: inst = 32'h10408000;
      8729: inst = 32'hc4044fb;
      8730: inst = 32'h8220000;
      8731: inst = 32'h10408000;
      8732: inst = 32'hc4044fc;
      8733: inst = 32'h8220000;
      8734: inst = 32'h10408000;
      8735: inst = 32'hc4044fd;
      8736: inst = 32'h8220000;
      8737: inst = 32'h10408000;
      8738: inst = 32'hc4044fe;
      8739: inst = 32'h8220000;
      8740: inst = 32'h10408000;
      8741: inst = 32'hc4044ff;
      8742: inst = 32'h8220000;
      8743: inst = 32'h10408000;
      8744: inst = 32'hc404500;
      8745: inst = 32'h8220000;
      8746: inst = 32'h10408000;
      8747: inst = 32'hc404501;
      8748: inst = 32'h8220000;
      8749: inst = 32'h10408000;
      8750: inst = 32'hc404502;
      8751: inst = 32'h8220000;
      8752: inst = 32'h10408000;
      8753: inst = 32'hc404503;
      8754: inst = 32'h8220000;
      8755: inst = 32'h10408000;
      8756: inst = 32'hc40453c;
      8757: inst = 32'h8220000;
      8758: inst = 32'h10408000;
      8759: inst = 32'hc40453d;
      8760: inst = 32'h8220000;
      8761: inst = 32'h10408000;
      8762: inst = 32'hc40453e;
      8763: inst = 32'h8220000;
      8764: inst = 32'h10408000;
      8765: inst = 32'hc40453f;
      8766: inst = 32'h8220000;
      8767: inst = 32'h10408000;
      8768: inst = 32'hc404540;
      8769: inst = 32'h8220000;
      8770: inst = 32'h10408000;
      8771: inst = 32'hc404541;
      8772: inst = 32'h8220000;
      8773: inst = 32'h10408000;
      8774: inst = 32'hc404542;
      8775: inst = 32'h8220000;
      8776: inst = 32'h10408000;
      8777: inst = 32'hc404543;
      8778: inst = 32'h8220000;
      8779: inst = 32'h10408000;
      8780: inst = 32'hc404544;
      8781: inst = 32'h8220000;
      8782: inst = 32'h10408000;
      8783: inst = 32'hc404545;
      8784: inst = 32'h8220000;
      8785: inst = 32'h10408000;
      8786: inst = 32'hc404546;
      8787: inst = 32'h8220000;
      8788: inst = 32'h10408000;
      8789: inst = 32'hc404547;
      8790: inst = 32'h8220000;
      8791: inst = 32'h10408000;
      8792: inst = 32'hc404548;
      8793: inst = 32'h8220000;
      8794: inst = 32'h10408000;
      8795: inst = 32'hc404549;
      8796: inst = 32'h8220000;
      8797: inst = 32'h10408000;
      8798: inst = 32'hc40454a;
      8799: inst = 32'h8220000;
      8800: inst = 32'h10408000;
      8801: inst = 32'hc40454b;
      8802: inst = 32'h8220000;
      8803: inst = 32'h10408000;
      8804: inst = 32'hc40454c;
      8805: inst = 32'h8220000;
      8806: inst = 32'h10408000;
      8807: inst = 32'hc40454d;
      8808: inst = 32'h8220000;
      8809: inst = 32'h10408000;
      8810: inst = 32'hc40454e;
      8811: inst = 32'h8220000;
      8812: inst = 32'h10408000;
      8813: inst = 32'hc40454f;
      8814: inst = 32'h8220000;
      8815: inst = 32'h10408000;
      8816: inst = 32'hc404550;
      8817: inst = 32'h8220000;
      8818: inst = 32'h10408000;
      8819: inst = 32'hc404551;
      8820: inst = 32'h8220000;
      8821: inst = 32'h10408000;
      8822: inst = 32'hc404552;
      8823: inst = 32'h8220000;
      8824: inst = 32'h10408000;
      8825: inst = 32'hc404553;
      8826: inst = 32'h8220000;
      8827: inst = 32'h10408000;
      8828: inst = 32'hc404554;
      8829: inst = 32'h8220000;
      8830: inst = 32'h10408000;
      8831: inst = 32'hc404555;
      8832: inst = 32'h8220000;
      8833: inst = 32'h10408000;
      8834: inst = 32'hc404556;
      8835: inst = 32'h8220000;
      8836: inst = 32'h10408000;
      8837: inst = 32'hc404557;
      8838: inst = 32'h8220000;
      8839: inst = 32'h10408000;
      8840: inst = 32'hc404558;
      8841: inst = 32'h8220000;
      8842: inst = 32'h10408000;
      8843: inst = 32'hc404559;
      8844: inst = 32'h8220000;
      8845: inst = 32'h10408000;
      8846: inst = 32'hc40455a;
      8847: inst = 32'h8220000;
      8848: inst = 32'h10408000;
      8849: inst = 32'hc40455b;
      8850: inst = 32'h8220000;
      8851: inst = 32'h10408000;
      8852: inst = 32'hc40455c;
      8853: inst = 32'h8220000;
      8854: inst = 32'h10408000;
      8855: inst = 32'hc40455d;
      8856: inst = 32'h8220000;
      8857: inst = 32'h10408000;
      8858: inst = 32'hc40455e;
      8859: inst = 32'h8220000;
      8860: inst = 32'h10408000;
      8861: inst = 32'hc40455f;
      8862: inst = 32'h8220000;
      8863: inst = 32'h10408000;
      8864: inst = 32'hc404560;
      8865: inst = 32'h8220000;
      8866: inst = 32'h10408000;
      8867: inst = 32'hc404561;
      8868: inst = 32'h8220000;
      8869: inst = 32'h10408000;
      8870: inst = 32'hc404562;
      8871: inst = 32'h8220000;
      8872: inst = 32'h10408000;
      8873: inst = 32'hc404563;
      8874: inst = 32'h8220000;
      8875: inst = 32'h10408000;
      8876: inst = 32'hc40459c;
      8877: inst = 32'h8220000;
      8878: inst = 32'h10408000;
      8879: inst = 32'hc40459d;
      8880: inst = 32'h8220000;
      8881: inst = 32'h10408000;
      8882: inst = 32'hc40459e;
      8883: inst = 32'h8220000;
      8884: inst = 32'h10408000;
      8885: inst = 32'hc40459f;
      8886: inst = 32'h8220000;
      8887: inst = 32'h10408000;
      8888: inst = 32'hc4045a0;
      8889: inst = 32'h8220000;
      8890: inst = 32'h10408000;
      8891: inst = 32'hc4045a1;
      8892: inst = 32'h8220000;
      8893: inst = 32'h10408000;
      8894: inst = 32'hc4045a2;
      8895: inst = 32'h8220000;
      8896: inst = 32'h10408000;
      8897: inst = 32'hc4045a3;
      8898: inst = 32'h8220000;
      8899: inst = 32'h10408000;
      8900: inst = 32'hc4045a4;
      8901: inst = 32'h8220000;
      8902: inst = 32'h10408000;
      8903: inst = 32'hc4045a5;
      8904: inst = 32'h8220000;
      8905: inst = 32'h10408000;
      8906: inst = 32'hc4045a6;
      8907: inst = 32'h8220000;
      8908: inst = 32'h10408000;
      8909: inst = 32'hc4045a7;
      8910: inst = 32'h8220000;
      8911: inst = 32'h10408000;
      8912: inst = 32'hc4045a8;
      8913: inst = 32'h8220000;
      8914: inst = 32'h10408000;
      8915: inst = 32'hc4045a9;
      8916: inst = 32'h8220000;
      8917: inst = 32'h10408000;
      8918: inst = 32'hc4045aa;
      8919: inst = 32'h8220000;
      8920: inst = 32'h10408000;
      8921: inst = 32'hc4045ab;
      8922: inst = 32'h8220000;
      8923: inst = 32'h10408000;
      8924: inst = 32'hc4045ac;
      8925: inst = 32'h8220000;
      8926: inst = 32'h10408000;
      8927: inst = 32'hc4045ad;
      8928: inst = 32'h8220000;
      8929: inst = 32'h10408000;
      8930: inst = 32'hc4045ae;
      8931: inst = 32'h8220000;
      8932: inst = 32'h10408000;
      8933: inst = 32'hc4045af;
      8934: inst = 32'h8220000;
      8935: inst = 32'h10408000;
      8936: inst = 32'hc4045b0;
      8937: inst = 32'h8220000;
      8938: inst = 32'h10408000;
      8939: inst = 32'hc4045b1;
      8940: inst = 32'h8220000;
      8941: inst = 32'h10408000;
      8942: inst = 32'hc4045b2;
      8943: inst = 32'h8220000;
      8944: inst = 32'h10408000;
      8945: inst = 32'hc4045b3;
      8946: inst = 32'h8220000;
      8947: inst = 32'h10408000;
      8948: inst = 32'hc4045b4;
      8949: inst = 32'h8220000;
      8950: inst = 32'h10408000;
      8951: inst = 32'hc4045b5;
      8952: inst = 32'h8220000;
      8953: inst = 32'h10408000;
      8954: inst = 32'hc4045b6;
      8955: inst = 32'h8220000;
      8956: inst = 32'h10408000;
      8957: inst = 32'hc4045b7;
      8958: inst = 32'h8220000;
      8959: inst = 32'h10408000;
      8960: inst = 32'hc4045b8;
      8961: inst = 32'h8220000;
      8962: inst = 32'h10408000;
      8963: inst = 32'hc4045b9;
      8964: inst = 32'h8220000;
      8965: inst = 32'h10408000;
      8966: inst = 32'hc4045ba;
      8967: inst = 32'h8220000;
      8968: inst = 32'h10408000;
      8969: inst = 32'hc4045bb;
      8970: inst = 32'h8220000;
      8971: inst = 32'h10408000;
      8972: inst = 32'hc4045bc;
      8973: inst = 32'h8220000;
      8974: inst = 32'h10408000;
      8975: inst = 32'hc4045bd;
      8976: inst = 32'h8220000;
      8977: inst = 32'h10408000;
      8978: inst = 32'hc4045be;
      8979: inst = 32'h8220000;
      8980: inst = 32'h10408000;
      8981: inst = 32'hc4045bf;
      8982: inst = 32'h8220000;
      8983: inst = 32'h10408000;
      8984: inst = 32'hc4045c0;
      8985: inst = 32'h8220000;
      8986: inst = 32'h10408000;
      8987: inst = 32'hc4045c1;
      8988: inst = 32'h8220000;
      8989: inst = 32'h10408000;
      8990: inst = 32'hc4045c2;
      8991: inst = 32'h8220000;
      8992: inst = 32'h10408000;
      8993: inst = 32'hc4045c3;
      8994: inst = 32'h8220000;
      8995: inst = 32'h10408000;
      8996: inst = 32'hc4045fc;
      8997: inst = 32'h8220000;
      8998: inst = 32'h10408000;
      8999: inst = 32'hc4045fd;
      9000: inst = 32'h8220000;
      9001: inst = 32'h10408000;
      9002: inst = 32'hc4045fe;
      9003: inst = 32'h8220000;
      9004: inst = 32'h10408000;
      9005: inst = 32'hc4045ff;
      9006: inst = 32'h8220000;
      9007: inst = 32'h10408000;
      9008: inst = 32'hc404600;
      9009: inst = 32'h8220000;
      9010: inst = 32'h10408000;
      9011: inst = 32'hc404601;
      9012: inst = 32'h8220000;
      9013: inst = 32'h10408000;
      9014: inst = 32'hc404602;
      9015: inst = 32'h8220000;
      9016: inst = 32'h10408000;
      9017: inst = 32'hc404603;
      9018: inst = 32'h8220000;
      9019: inst = 32'h10408000;
      9020: inst = 32'hc404604;
      9021: inst = 32'h8220000;
      9022: inst = 32'h10408000;
      9023: inst = 32'hc404605;
      9024: inst = 32'h8220000;
      9025: inst = 32'h10408000;
      9026: inst = 32'hc404606;
      9027: inst = 32'h8220000;
      9028: inst = 32'h10408000;
      9029: inst = 32'hc404607;
      9030: inst = 32'h8220000;
      9031: inst = 32'h10408000;
      9032: inst = 32'hc404608;
      9033: inst = 32'h8220000;
      9034: inst = 32'h10408000;
      9035: inst = 32'hc404609;
      9036: inst = 32'h8220000;
      9037: inst = 32'h10408000;
      9038: inst = 32'hc40460a;
      9039: inst = 32'h8220000;
      9040: inst = 32'h10408000;
      9041: inst = 32'hc40460b;
      9042: inst = 32'h8220000;
      9043: inst = 32'h10408000;
      9044: inst = 32'hc40460c;
      9045: inst = 32'h8220000;
      9046: inst = 32'h10408000;
      9047: inst = 32'hc40460d;
      9048: inst = 32'h8220000;
      9049: inst = 32'h10408000;
      9050: inst = 32'hc40460e;
      9051: inst = 32'h8220000;
      9052: inst = 32'h10408000;
      9053: inst = 32'hc40460f;
      9054: inst = 32'h8220000;
      9055: inst = 32'h10408000;
      9056: inst = 32'hc404610;
      9057: inst = 32'h8220000;
      9058: inst = 32'h10408000;
      9059: inst = 32'hc404611;
      9060: inst = 32'h8220000;
      9061: inst = 32'h10408000;
      9062: inst = 32'hc404612;
      9063: inst = 32'h8220000;
      9064: inst = 32'h10408000;
      9065: inst = 32'hc404613;
      9066: inst = 32'h8220000;
      9067: inst = 32'h10408000;
      9068: inst = 32'hc404614;
      9069: inst = 32'h8220000;
      9070: inst = 32'h10408000;
      9071: inst = 32'hc404615;
      9072: inst = 32'h8220000;
      9073: inst = 32'h10408000;
      9074: inst = 32'hc404616;
      9075: inst = 32'h8220000;
      9076: inst = 32'h10408000;
      9077: inst = 32'hc404617;
      9078: inst = 32'h8220000;
      9079: inst = 32'h10408000;
      9080: inst = 32'hc404618;
      9081: inst = 32'h8220000;
      9082: inst = 32'h10408000;
      9083: inst = 32'hc404619;
      9084: inst = 32'h8220000;
      9085: inst = 32'h10408000;
      9086: inst = 32'hc40461a;
      9087: inst = 32'h8220000;
      9088: inst = 32'h10408000;
      9089: inst = 32'hc40461b;
      9090: inst = 32'h8220000;
      9091: inst = 32'h10408000;
      9092: inst = 32'hc40461c;
      9093: inst = 32'h8220000;
      9094: inst = 32'h10408000;
      9095: inst = 32'hc40461d;
      9096: inst = 32'h8220000;
      9097: inst = 32'h10408000;
      9098: inst = 32'hc40461e;
      9099: inst = 32'h8220000;
      9100: inst = 32'h10408000;
      9101: inst = 32'hc40461f;
      9102: inst = 32'h8220000;
      9103: inst = 32'h10408000;
      9104: inst = 32'hc404620;
      9105: inst = 32'h8220000;
      9106: inst = 32'h10408000;
      9107: inst = 32'hc404621;
      9108: inst = 32'h8220000;
      9109: inst = 32'h10408000;
      9110: inst = 32'hc404622;
      9111: inst = 32'h8220000;
      9112: inst = 32'h10408000;
      9113: inst = 32'hc404623;
      9114: inst = 32'h8220000;
      9115: inst = 32'h10408000;
      9116: inst = 32'hc40465c;
      9117: inst = 32'h8220000;
      9118: inst = 32'h10408000;
      9119: inst = 32'hc40465d;
      9120: inst = 32'h8220000;
      9121: inst = 32'h10408000;
      9122: inst = 32'hc40465e;
      9123: inst = 32'h8220000;
      9124: inst = 32'h10408000;
      9125: inst = 32'hc40465f;
      9126: inst = 32'h8220000;
      9127: inst = 32'h10408000;
      9128: inst = 32'hc404660;
      9129: inst = 32'h8220000;
      9130: inst = 32'h10408000;
      9131: inst = 32'hc404661;
      9132: inst = 32'h8220000;
      9133: inst = 32'h10408000;
      9134: inst = 32'hc404662;
      9135: inst = 32'h8220000;
      9136: inst = 32'h10408000;
      9137: inst = 32'hc404663;
      9138: inst = 32'h8220000;
      9139: inst = 32'h10408000;
      9140: inst = 32'hc404664;
      9141: inst = 32'h8220000;
      9142: inst = 32'h10408000;
      9143: inst = 32'hc404665;
      9144: inst = 32'h8220000;
      9145: inst = 32'h10408000;
      9146: inst = 32'hc404666;
      9147: inst = 32'h8220000;
      9148: inst = 32'h10408000;
      9149: inst = 32'hc404667;
      9150: inst = 32'h8220000;
      9151: inst = 32'h10408000;
      9152: inst = 32'hc404668;
      9153: inst = 32'h8220000;
      9154: inst = 32'h10408000;
      9155: inst = 32'hc404669;
      9156: inst = 32'h8220000;
      9157: inst = 32'h10408000;
      9158: inst = 32'hc40466a;
      9159: inst = 32'h8220000;
      9160: inst = 32'h10408000;
      9161: inst = 32'hc40466b;
      9162: inst = 32'h8220000;
      9163: inst = 32'h10408000;
      9164: inst = 32'hc40466c;
      9165: inst = 32'h8220000;
      9166: inst = 32'h10408000;
      9167: inst = 32'hc40466d;
      9168: inst = 32'h8220000;
      9169: inst = 32'h10408000;
      9170: inst = 32'hc40466e;
      9171: inst = 32'h8220000;
      9172: inst = 32'h10408000;
      9173: inst = 32'hc40466f;
      9174: inst = 32'h8220000;
      9175: inst = 32'h10408000;
      9176: inst = 32'hc404670;
      9177: inst = 32'h8220000;
      9178: inst = 32'h10408000;
      9179: inst = 32'hc404671;
      9180: inst = 32'h8220000;
      9181: inst = 32'h10408000;
      9182: inst = 32'hc404672;
      9183: inst = 32'h8220000;
      9184: inst = 32'h10408000;
      9185: inst = 32'hc404673;
      9186: inst = 32'h8220000;
      9187: inst = 32'h10408000;
      9188: inst = 32'hc404674;
      9189: inst = 32'h8220000;
      9190: inst = 32'h10408000;
      9191: inst = 32'hc404675;
      9192: inst = 32'h8220000;
      9193: inst = 32'h10408000;
      9194: inst = 32'hc404676;
      9195: inst = 32'h8220000;
      9196: inst = 32'h10408000;
      9197: inst = 32'hc404677;
      9198: inst = 32'h8220000;
      9199: inst = 32'h10408000;
      9200: inst = 32'hc404678;
      9201: inst = 32'h8220000;
      9202: inst = 32'h10408000;
      9203: inst = 32'hc404679;
      9204: inst = 32'h8220000;
      9205: inst = 32'h10408000;
      9206: inst = 32'hc40467a;
      9207: inst = 32'h8220000;
      9208: inst = 32'h10408000;
      9209: inst = 32'hc40467b;
      9210: inst = 32'h8220000;
      9211: inst = 32'h10408000;
      9212: inst = 32'hc40467c;
      9213: inst = 32'h8220000;
      9214: inst = 32'h10408000;
      9215: inst = 32'hc40467d;
      9216: inst = 32'h8220000;
      9217: inst = 32'h10408000;
      9218: inst = 32'hc40467e;
      9219: inst = 32'h8220000;
      9220: inst = 32'h10408000;
      9221: inst = 32'hc40467f;
      9222: inst = 32'h8220000;
      9223: inst = 32'h10408000;
      9224: inst = 32'hc404680;
      9225: inst = 32'h8220000;
      9226: inst = 32'h10408000;
      9227: inst = 32'hc404681;
      9228: inst = 32'h8220000;
      9229: inst = 32'h10408000;
      9230: inst = 32'hc404682;
      9231: inst = 32'h8220000;
      9232: inst = 32'h10408000;
      9233: inst = 32'hc404683;
      9234: inst = 32'h8220000;
      9235: inst = 32'h10408000;
      9236: inst = 32'hc4046bc;
      9237: inst = 32'h8220000;
      9238: inst = 32'h10408000;
      9239: inst = 32'hc4046bd;
      9240: inst = 32'h8220000;
      9241: inst = 32'h10408000;
      9242: inst = 32'hc4046be;
      9243: inst = 32'h8220000;
      9244: inst = 32'h10408000;
      9245: inst = 32'hc4046bf;
      9246: inst = 32'h8220000;
      9247: inst = 32'h10408000;
      9248: inst = 32'hc4046c0;
      9249: inst = 32'h8220000;
      9250: inst = 32'h10408000;
      9251: inst = 32'hc4046c1;
      9252: inst = 32'h8220000;
      9253: inst = 32'h10408000;
      9254: inst = 32'hc4046c2;
      9255: inst = 32'h8220000;
      9256: inst = 32'h10408000;
      9257: inst = 32'hc4046c3;
      9258: inst = 32'h8220000;
      9259: inst = 32'h10408000;
      9260: inst = 32'hc4046c4;
      9261: inst = 32'h8220000;
      9262: inst = 32'h10408000;
      9263: inst = 32'hc4046c5;
      9264: inst = 32'h8220000;
      9265: inst = 32'h10408000;
      9266: inst = 32'hc4046c6;
      9267: inst = 32'h8220000;
      9268: inst = 32'h10408000;
      9269: inst = 32'hc4046c7;
      9270: inst = 32'h8220000;
      9271: inst = 32'h10408000;
      9272: inst = 32'hc4046c8;
      9273: inst = 32'h8220000;
      9274: inst = 32'h10408000;
      9275: inst = 32'hc4046c9;
      9276: inst = 32'h8220000;
      9277: inst = 32'h10408000;
      9278: inst = 32'hc4046ca;
      9279: inst = 32'h8220000;
      9280: inst = 32'h10408000;
      9281: inst = 32'hc4046cb;
      9282: inst = 32'h8220000;
      9283: inst = 32'h10408000;
      9284: inst = 32'hc4046cc;
      9285: inst = 32'h8220000;
      9286: inst = 32'h10408000;
      9287: inst = 32'hc4046cd;
      9288: inst = 32'h8220000;
      9289: inst = 32'h10408000;
      9290: inst = 32'hc4046ce;
      9291: inst = 32'h8220000;
      9292: inst = 32'h10408000;
      9293: inst = 32'hc4046cf;
      9294: inst = 32'h8220000;
      9295: inst = 32'h10408000;
      9296: inst = 32'hc4046d0;
      9297: inst = 32'h8220000;
      9298: inst = 32'h10408000;
      9299: inst = 32'hc4046d1;
      9300: inst = 32'h8220000;
      9301: inst = 32'h10408000;
      9302: inst = 32'hc4046d2;
      9303: inst = 32'h8220000;
      9304: inst = 32'h10408000;
      9305: inst = 32'hc4046d3;
      9306: inst = 32'h8220000;
      9307: inst = 32'h10408000;
      9308: inst = 32'hc4046d4;
      9309: inst = 32'h8220000;
      9310: inst = 32'h10408000;
      9311: inst = 32'hc4046d5;
      9312: inst = 32'h8220000;
      9313: inst = 32'h10408000;
      9314: inst = 32'hc4046d6;
      9315: inst = 32'h8220000;
      9316: inst = 32'h10408000;
      9317: inst = 32'hc4046d7;
      9318: inst = 32'h8220000;
      9319: inst = 32'h10408000;
      9320: inst = 32'hc4046d8;
      9321: inst = 32'h8220000;
      9322: inst = 32'h10408000;
      9323: inst = 32'hc4046d9;
      9324: inst = 32'h8220000;
      9325: inst = 32'h10408000;
      9326: inst = 32'hc4046da;
      9327: inst = 32'h8220000;
      9328: inst = 32'h10408000;
      9329: inst = 32'hc4046db;
      9330: inst = 32'h8220000;
      9331: inst = 32'h10408000;
      9332: inst = 32'hc4046dc;
      9333: inst = 32'h8220000;
      9334: inst = 32'h10408000;
      9335: inst = 32'hc4046dd;
      9336: inst = 32'h8220000;
      9337: inst = 32'h10408000;
      9338: inst = 32'hc4046de;
      9339: inst = 32'h8220000;
      9340: inst = 32'h10408000;
      9341: inst = 32'hc4046df;
      9342: inst = 32'h8220000;
      9343: inst = 32'h10408000;
      9344: inst = 32'hc4046e0;
      9345: inst = 32'h8220000;
      9346: inst = 32'h10408000;
      9347: inst = 32'hc4046e1;
      9348: inst = 32'h8220000;
      9349: inst = 32'h10408000;
      9350: inst = 32'hc4046e2;
      9351: inst = 32'h8220000;
      9352: inst = 32'h10408000;
      9353: inst = 32'hc4046e3;
      9354: inst = 32'h8220000;
      9355: inst = 32'h10408000;
      9356: inst = 32'hc40471c;
      9357: inst = 32'h8220000;
      9358: inst = 32'h10408000;
      9359: inst = 32'hc40471d;
      9360: inst = 32'h8220000;
      9361: inst = 32'h10408000;
      9362: inst = 32'hc40471e;
      9363: inst = 32'h8220000;
      9364: inst = 32'h10408000;
      9365: inst = 32'hc40471f;
      9366: inst = 32'h8220000;
      9367: inst = 32'h10408000;
      9368: inst = 32'hc404720;
      9369: inst = 32'h8220000;
      9370: inst = 32'h10408000;
      9371: inst = 32'hc404721;
      9372: inst = 32'h8220000;
      9373: inst = 32'h10408000;
      9374: inst = 32'hc404722;
      9375: inst = 32'h8220000;
      9376: inst = 32'h10408000;
      9377: inst = 32'hc404723;
      9378: inst = 32'h8220000;
      9379: inst = 32'h10408000;
      9380: inst = 32'hc404724;
      9381: inst = 32'h8220000;
      9382: inst = 32'h10408000;
      9383: inst = 32'hc404725;
      9384: inst = 32'h8220000;
      9385: inst = 32'h10408000;
      9386: inst = 32'hc404726;
      9387: inst = 32'h8220000;
      9388: inst = 32'h10408000;
      9389: inst = 32'hc404727;
      9390: inst = 32'h8220000;
      9391: inst = 32'h10408000;
      9392: inst = 32'hc404728;
      9393: inst = 32'h8220000;
      9394: inst = 32'h10408000;
      9395: inst = 32'hc404729;
      9396: inst = 32'h8220000;
      9397: inst = 32'h10408000;
      9398: inst = 32'hc40472a;
      9399: inst = 32'h8220000;
      9400: inst = 32'h10408000;
      9401: inst = 32'hc40472b;
      9402: inst = 32'h8220000;
      9403: inst = 32'h10408000;
      9404: inst = 32'hc40472c;
      9405: inst = 32'h8220000;
      9406: inst = 32'h10408000;
      9407: inst = 32'hc40472d;
      9408: inst = 32'h8220000;
      9409: inst = 32'h10408000;
      9410: inst = 32'hc40472e;
      9411: inst = 32'h8220000;
      9412: inst = 32'h10408000;
      9413: inst = 32'hc40472f;
      9414: inst = 32'h8220000;
      9415: inst = 32'h10408000;
      9416: inst = 32'hc404730;
      9417: inst = 32'h8220000;
      9418: inst = 32'h10408000;
      9419: inst = 32'hc404731;
      9420: inst = 32'h8220000;
      9421: inst = 32'h10408000;
      9422: inst = 32'hc404732;
      9423: inst = 32'h8220000;
      9424: inst = 32'h10408000;
      9425: inst = 32'hc404733;
      9426: inst = 32'h8220000;
      9427: inst = 32'h10408000;
      9428: inst = 32'hc404734;
      9429: inst = 32'h8220000;
      9430: inst = 32'h10408000;
      9431: inst = 32'hc404735;
      9432: inst = 32'h8220000;
      9433: inst = 32'h10408000;
      9434: inst = 32'hc404736;
      9435: inst = 32'h8220000;
      9436: inst = 32'h10408000;
      9437: inst = 32'hc404737;
      9438: inst = 32'h8220000;
      9439: inst = 32'h10408000;
      9440: inst = 32'hc404738;
      9441: inst = 32'h8220000;
      9442: inst = 32'h10408000;
      9443: inst = 32'hc404739;
      9444: inst = 32'h8220000;
      9445: inst = 32'h10408000;
      9446: inst = 32'hc40473a;
      9447: inst = 32'h8220000;
      9448: inst = 32'h10408000;
      9449: inst = 32'hc40473b;
      9450: inst = 32'h8220000;
      9451: inst = 32'h10408000;
      9452: inst = 32'hc40473c;
      9453: inst = 32'h8220000;
      9454: inst = 32'h10408000;
      9455: inst = 32'hc40473d;
      9456: inst = 32'h8220000;
      9457: inst = 32'h10408000;
      9458: inst = 32'hc40473e;
      9459: inst = 32'h8220000;
      9460: inst = 32'h10408000;
      9461: inst = 32'hc40473f;
      9462: inst = 32'h8220000;
      9463: inst = 32'h10408000;
      9464: inst = 32'hc404740;
      9465: inst = 32'h8220000;
      9466: inst = 32'h10408000;
      9467: inst = 32'hc404741;
      9468: inst = 32'h8220000;
      9469: inst = 32'h10408000;
      9470: inst = 32'hc404742;
      9471: inst = 32'h8220000;
      9472: inst = 32'h10408000;
      9473: inst = 32'hc404743;
      9474: inst = 32'h8220000;
      9475: inst = 32'h10408000;
      9476: inst = 32'hc40477c;
      9477: inst = 32'h8220000;
      9478: inst = 32'h10408000;
      9479: inst = 32'hc40477d;
      9480: inst = 32'h8220000;
      9481: inst = 32'h10408000;
      9482: inst = 32'hc40477e;
      9483: inst = 32'h8220000;
      9484: inst = 32'h10408000;
      9485: inst = 32'hc40477f;
      9486: inst = 32'h8220000;
      9487: inst = 32'h10408000;
      9488: inst = 32'hc404780;
      9489: inst = 32'h8220000;
      9490: inst = 32'h10408000;
      9491: inst = 32'hc404781;
      9492: inst = 32'h8220000;
      9493: inst = 32'h10408000;
      9494: inst = 32'hc404782;
      9495: inst = 32'h8220000;
      9496: inst = 32'h10408000;
      9497: inst = 32'hc404783;
      9498: inst = 32'h8220000;
      9499: inst = 32'h10408000;
      9500: inst = 32'hc404784;
      9501: inst = 32'h8220000;
      9502: inst = 32'h10408000;
      9503: inst = 32'hc404785;
      9504: inst = 32'h8220000;
      9505: inst = 32'h10408000;
      9506: inst = 32'hc404786;
      9507: inst = 32'h8220000;
      9508: inst = 32'h10408000;
      9509: inst = 32'hc404787;
      9510: inst = 32'h8220000;
      9511: inst = 32'h10408000;
      9512: inst = 32'hc404788;
      9513: inst = 32'h8220000;
      9514: inst = 32'h10408000;
      9515: inst = 32'hc404789;
      9516: inst = 32'h8220000;
      9517: inst = 32'h10408000;
      9518: inst = 32'hc40478a;
      9519: inst = 32'h8220000;
      9520: inst = 32'h10408000;
      9521: inst = 32'hc40478b;
      9522: inst = 32'h8220000;
      9523: inst = 32'h10408000;
      9524: inst = 32'hc40478c;
      9525: inst = 32'h8220000;
      9526: inst = 32'h10408000;
      9527: inst = 32'hc40478d;
      9528: inst = 32'h8220000;
      9529: inst = 32'h10408000;
      9530: inst = 32'hc40478e;
      9531: inst = 32'h8220000;
      9532: inst = 32'h10408000;
      9533: inst = 32'hc40478f;
      9534: inst = 32'h8220000;
      9535: inst = 32'h10408000;
      9536: inst = 32'hc404790;
      9537: inst = 32'h8220000;
      9538: inst = 32'h10408000;
      9539: inst = 32'hc404791;
      9540: inst = 32'h8220000;
      9541: inst = 32'h10408000;
      9542: inst = 32'hc404792;
      9543: inst = 32'h8220000;
      9544: inst = 32'h10408000;
      9545: inst = 32'hc404793;
      9546: inst = 32'h8220000;
      9547: inst = 32'h10408000;
      9548: inst = 32'hc404794;
      9549: inst = 32'h8220000;
      9550: inst = 32'h10408000;
      9551: inst = 32'hc404795;
      9552: inst = 32'h8220000;
      9553: inst = 32'h10408000;
      9554: inst = 32'hc404796;
      9555: inst = 32'h8220000;
      9556: inst = 32'h10408000;
      9557: inst = 32'hc404797;
      9558: inst = 32'h8220000;
      9559: inst = 32'h10408000;
      9560: inst = 32'hc404798;
      9561: inst = 32'h8220000;
      9562: inst = 32'h10408000;
      9563: inst = 32'hc404799;
      9564: inst = 32'h8220000;
      9565: inst = 32'h10408000;
      9566: inst = 32'hc40479a;
      9567: inst = 32'h8220000;
      9568: inst = 32'h10408000;
      9569: inst = 32'hc40479b;
      9570: inst = 32'h8220000;
      9571: inst = 32'h10408000;
      9572: inst = 32'hc40479c;
      9573: inst = 32'h8220000;
      9574: inst = 32'h10408000;
      9575: inst = 32'hc40479d;
      9576: inst = 32'h8220000;
      9577: inst = 32'h10408000;
      9578: inst = 32'hc40479e;
      9579: inst = 32'h8220000;
      9580: inst = 32'h10408000;
      9581: inst = 32'hc40479f;
      9582: inst = 32'h8220000;
      9583: inst = 32'h10408000;
      9584: inst = 32'hc4047a0;
      9585: inst = 32'h8220000;
      9586: inst = 32'h10408000;
      9587: inst = 32'hc4047a1;
      9588: inst = 32'h8220000;
      9589: inst = 32'h10408000;
      9590: inst = 32'hc4047a2;
      9591: inst = 32'h8220000;
      9592: inst = 32'h10408000;
      9593: inst = 32'hc4047a3;
      9594: inst = 32'h8220000;
      9595: inst = 32'h10408000;
      9596: inst = 32'hc4047dc;
      9597: inst = 32'h8220000;
      9598: inst = 32'h10408000;
      9599: inst = 32'hc4047dd;
      9600: inst = 32'h8220000;
      9601: inst = 32'h10408000;
      9602: inst = 32'hc4047de;
      9603: inst = 32'h8220000;
      9604: inst = 32'h10408000;
      9605: inst = 32'hc4047df;
      9606: inst = 32'h8220000;
      9607: inst = 32'h10408000;
      9608: inst = 32'hc4047e0;
      9609: inst = 32'h8220000;
      9610: inst = 32'h10408000;
      9611: inst = 32'hc4047e1;
      9612: inst = 32'h8220000;
      9613: inst = 32'h10408000;
      9614: inst = 32'hc4047e2;
      9615: inst = 32'h8220000;
      9616: inst = 32'h10408000;
      9617: inst = 32'hc4047e3;
      9618: inst = 32'h8220000;
      9619: inst = 32'h10408000;
      9620: inst = 32'hc4047e4;
      9621: inst = 32'h8220000;
      9622: inst = 32'h10408000;
      9623: inst = 32'hc4047e5;
      9624: inst = 32'h8220000;
      9625: inst = 32'h10408000;
      9626: inst = 32'hc4047e6;
      9627: inst = 32'h8220000;
      9628: inst = 32'h10408000;
      9629: inst = 32'hc4047e7;
      9630: inst = 32'h8220000;
      9631: inst = 32'h10408000;
      9632: inst = 32'hc4047e8;
      9633: inst = 32'h8220000;
      9634: inst = 32'h10408000;
      9635: inst = 32'hc4047e9;
      9636: inst = 32'h8220000;
      9637: inst = 32'h10408000;
      9638: inst = 32'hc4047ea;
      9639: inst = 32'h8220000;
      9640: inst = 32'h10408000;
      9641: inst = 32'hc4047eb;
      9642: inst = 32'h8220000;
      9643: inst = 32'h10408000;
      9644: inst = 32'hc4047ec;
      9645: inst = 32'h8220000;
      9646: inst = 32'h10408000;
      9647: inst = 32'hc4047ed;
      9648: inst = 32'h8220000;
      9649: inst = 32'h10408000;
      9650: inst = 32'hc4047ee;
      9651: inst = 32'h8220000;
      9652: inst = 32'h10408000;
      9653: inst = 32'hc4047ef;
      9654: inst = 32'h8220000;
      9655: inst = 32'h10408000;
      9656: inst = 32'hc4047f0;
      9657: inst = 32'h8220000;
      9658: inst = 32'h10408000;
      9659: inst = 32'hc4047f1;
      9660: inst = 32'h8220000;
      9661: inst = 32'h10408000;
      9662: inst = 32'hc4047f2;
      9663: inst = 32'h8220000;
      9664: inst = 32'h10408000;
      9665: inst = 32'hc4047f3;
      9666: inst = 32'h8220000;
      9667: inst = 32'h10408000;
      9668: inst = 32'hc4047f4;
      9669: inst = 32'h8220000;
      9670: inst = 32'h10408000;
      9671: inst = 32'hc4047f5;
      9672: inst = 32'h8220000;
      9673: inst = 32'h10408000;
      9674: inst = 32'hc4047f6;
      9675: inst = 32'h8220000;
      9676: inst = 32'h10408000;
      9677: inst = 32'hc4047f7;
      9678: inst = 32'h8220000;
      9679: inst = 32'h10408000;
      9680: inst = 32'hc4047f8;
      9681: inst = 32'h8220000;
      9682: inst = 32'h10408000;
      9683: inst = 32'hc4047f9;
      9684: inst = 32'h8220000;
      9685: inst = 32'h10408000;
      9686: inst = 32'hc4047fa;
      9687: inst = 32'h8220000;
      9688: inst = 32'h10408000;
      9689: inst = 32'hc4047fb;
      9690: inst = 32'h8220000;
      9691: inst = 32'h10408000;
      9692: inst = 32'hc4047fc;
      9693: inst = 32'h8220000;
      9694: inst = 32'h10408000;
      9695: inst = 32'hc4047fd;
      9696: inst = 32'h8220000;
      9697: inst = 32'h10408000;
      9698: inst = 32'hc4047fe;
      9699: inst = 32'h8220000;
      9700: inst = 32'h10408000;
      9701: inst = 32'hc4047ff;
      9702: inst = 32'h8220000;
      9703: inst = 32'h10408000;
      9704: inst = 32'hc404800;
      9705: inst = 32'h8220000;
      9706: inst = 32'h10408000;
      9707: inst = 32'hc404801;
      9708: inst = 32'h8220000;
      9709: inst = 32'h10408000;
      9710: inst = 32'hc404802;
      9711: inst = 32'h8220000;
      9712: inst = 32'h10408000;
      9713: inst = 32'hc404803;
      9714: inst = 32'h8220000;
      9715: inst = 32'h10408000;
      9716: inst = 32'hc40483c;
      9717: inst = 32'h8220000;
      9718: inst = 32'h10408000;
      9719: inst = 32'hc40483d;
      9720: inst = 32'h8220000;
      9721: inst = 32'h10408000;
      9722: inst = 32'hc40483e;
      9723: inst = 32'h8220000;
      9724: inst = 32'h10408000;
      9725: inst = 32'hc40483f;
      9726: inst = 32'h8220000;
      9727: inst = 32'h10408000;
      9728: inst = 32'hc404840;
      9729: inst = 32'h8220000;
      9730: inst = 32'h10408000;
      9731: inst = 32'hc404841;
      9732: inst = 32'h8220000;
      9733: inst = 32'h10408000;
      9734: inst = 32'hc404842;
      9735: inst = 32'h8220000;
      9736: inst = 32'h10408000;
      9737: inst = 32'hc404843;
      9738: inst = 32'h8220000;
      9739: inst = 32'h10408000;
      9740: inst = 32'hc404844;
      9741: inst = 32'h8220000;
      9742: inst = 32'h10408000;
      9743: inst = 32'hc404845;
      9744: inst = 32'h8220000;
      9745: inst = 32'h10408000;
      9746: inst = 32'hc404846;
      9747: inst = 32'h8220000;
      9748: inst = 32'h10408000;
      9749: inst = 32'hc404847;
      9750: inst = 32'h8220000;
      9751: inst = 32'h10408000;
      9752: inst = 32'hc404848;
      9753: inst = 32'h8220000;
      9754: inst = 32'h10408000;
      9755: inst = 32'hc404849;
      9756: inst = 32'h8220000;
      9757: inst = 32'h10408000;
      9758: inst = 32'hc40484a;
      9759: inst = 32'h8220000;
      9760: inst = 32'h10408000;
      9761: inst = 32'hc40484b;
      9762: inst = 32'h8220000;
      9763: inst = 32'h10408000;
      9764: inst = 32'hc40484c;
      9765: inst = 32'h8220000;
      9766: inst = 32'h10408000;
      9767: inst = 32'hc40484d;
      9768: inst = 32'h8220000;
      9769: inst = 32'h10408000;
      9770: inst = 32'hc40484e;
      9771: inst = 32'h8220000;
      9772: inst = 32'h10408000;
      9773: inst = 32'hc40484f;
      9774: inst = 32'h8220000;
      9775: inst = 32'h10408000;
      9776: inst = 32'hc404850;
      9777: inst = 32'h8220000;
      9778: inst = 32'h10408000;
      9779: inst = 32'hc404851;
      9780: inst = 32'h8220000;
      9781: inst = 32'h10408000;
      9782: inst = 32'hc404852;
      9783: inst = 32'h8220000;
      9784: inst = 32'h10408000;
      9785: inst = 32'hc404853;
      9786: inst = 32'h8220000;
      9787: inst = 32'h10408000;
      9788: inst = 32'hc404854;
      9789: inst = 32'h8220000;
      9790: inst = 32'h10408000;
      9791: inst = 32'hc404855;
      9792: inst = 32'h8220000;
      9793: inst = 32'h10408000;
      9794: inst = 32'hc404856;
      9795: inst = 32'h8220000;
      9796: inst = 32'h10408000;
      9797: inst = 32'hc404857;
      9798: inst = 32'h8220000;
      9799: inst = 32'h10408000;
      9800: inst = 32'hc404858;
      9801: inst = 32'h8220000;
      9802: inst = 32'h10408000;
      9803: inst = 32'hc404859;
      9804: inst = 32'h8220000;
      9805: inst = 32'h10408000;
      9806: inst = 32'hc40485a;
      9807: inst = 32'h8220000;
      9808: inst = 32'h10408000;
      9809: inst = 32'hc40485b;
      9810: inst = 32'h8220000;
      9811: inst = 32'h10408000;
      9812: inst = 32'hc40485c;
      9813: inst = 32'h8220000;
      9814: inst = 32'h10408000;
      9815: inst = 32'hc40485d;
      9816: inst = 32'h8220000;
      9817: inst = 32'h10408000;
      9818: inst = 32'hc40485e;
      9819: inst = 32'h8220000;
      9820: inst = 32'h10408000;
      9821: inst = 32'hc40485f;
      9822: inst = 32'h8220000;
      9823: inst = 32'h10408000;
      9824: inst = 32'hc404860;
      9825: inst = 32'h8220000;
      9826: inst = 32'h10408000;
      9827: inst = 32'hc404861;
      9828: inst = 32'h8220000;
      9829: inst = 32'h10408000;
      9830: inst = 32'hc404862;
      9831: inst = 32'h8220000;
      9832: inst = 32'h10408000;
      9833: inst = 32'hc404863;
      9834: inst = 32'h8220000;
      9835: inst = 32'h10408000;
      9836: inst = 32'hc40489c;
      9837: inst = 32'h8220000;
      9838: inst = 32'h10408000;
      9839: inst = 32'hc40489d;
      9840: inst = 32'h8220000;
      9841: inst = 32'h10408000;
      9842: inst = 32'hc40489e;
      9843: inst = 32'h8220000;
      9844: inst = 32'h10408000;
      9845: inst = 32'hc40489f;
      9846: inst = 32'h8220000;
      9847: inst = 32'h10408000;
      9848: inst = 32'hc4048a0;
      9849: inst = 32'h8220000;
      9850: inst = 32'h10408000;
      9851: inst = 32'hc4048a1;
      9852: inst = 32'h8220000;
      9853: inst = 32'h10408000;
      9854: inst = 32'hc4048a2;
      9855: inst = 32'h8220000;
      9856: inst = 32'h10408000;
      9857: inst = 32'hc4048a3;
      9858: inst = 32'h8220000;
      9859: inst = 32'h10408000;
      9860: inst = 32'hc4048a4;
      9861: inst = 32'h8220000;
      9862: inst = 32'h10408000;
      9863: inst = 32'hc4048a5;
      9864: inst = 32'h8220000;
      9865: inst = 32'h10408000;
      9866: inst = 32'hc4048a6;
      9867: inst = 32'h8220000;
      9868: inst = 32'h10408000;
      9869: inst = 32'hc4048a7;
      9870: inst = 32'h8220000;
      9871: inst = 32'h10408000;
      9872: inst = 32'hc4048a8;
      9873: inst = 32'h8220000;
      9874: inst = 32'h10408000;
      9875: inst = 32'hc4048a9;
      9876: inst = 32'h8220000;
      9877: inst = 32'h10408000;
      9878: inst = 32'hc4048aa;
      9879: inst = 32'h8220000;
      9880: inst = 32'h10408000;
      9881: inst = 32'hc4048ab;
      9882: inst = 32'h8220000;
      9883: inst = 32'h10408000;
      9884: inst = 32'hc4048ac;
      9885: inst = 32'h8220000;
      9886: inst = 32'h10408000;
      9887: inst = 32'hc4048ad;
      9888: inst = 32'h8220000;
      9889: inst = 32'h10408000;
      9890: inst = 32'hc4048ae;
      9891: inst = 32'h8220000;
      9892: inst = 32'h10408000;
      9893: inst = 32'hc4048af;
      9894: inst = 32'h8220000;
      9895: inst = 32'h10408000;
      9896: inst = 32'hc4048b0;
      9897: inst = 32'h8220000;
      9898: inst = 32'h10408000;
      9899: inst = 32'hc4048b1;
      9900: inst = 32'h8220000;
      9901: inst = 32'h10408000;
      9902: inst = 32'hc4048b2;
      9903: inst = 32'h8220000;
      9904: inst = 32'h10408000;
      9905: inst = 32'hc4048b3;
      9906: inst = 32'h8220000;
      9907: inst = 32'h10408000;
      9908: inst = 32'hc4048b4;
      9909: inst = 32'h8220000;
      9910: inst = 32'h10408000;
      9911: inst = 32'hc4048b5;
      9912: inst = 32'h8220000;
      9913: inst = 32'h10408000;
      9914: inst = 32'hc4048b6;
      9915: inst = 32'h8220000;
      9916: inst = 32'h10408000;
      9917: inst = 32'hc4048b7;
      9918: inst = 32'h8220000;
      9919: inst = 32'h10408000;
      9920: inst = 32'hc4048b8;
      9921: inst = 32'h8220000;
      9922: inst = 32'h10408000;
      9923: inst = 32'hc4048b9;
      9924: inst = 32'h8220000;
      9925: inst = 32'h10408000;
      9926: inst = 32'hc4048ba;
      9927: inst = 32'h8220000;
      9928: inst = 32'h10408000;
      9929: inst = 32'hc4048bb;
      9930: inst = 32'h8220000;
      9931: inst = 32'h10408000;
      9932: inst = 32'hc4048bc;
      9933: inst = 32'h8220000;
      9934: inst = 32'h10408000;
      9935: inst = 32'hc4048bd;
      9936: inst = 32'h8220000;
      9937: inst = 32'h10408000;
      9938: inst = 32'hc4048be;
      9939: inst = 32'h8220000;
      9940: inst = 32'h10408000;
      9941: inst = 32'hc4048bf;
      9942: inst = 32'h8220000;
      9943: inst = 32'h10408000;
      9944: inst = 32'hc4048c0;
      9945: inst = 32'h8220000;
      9946: inst = 32'h10408000;
      9947: inst = 32'hc4048c1;
      9948: inst = 32'h8220000;
      9949: inst = 32'h10408000;
      9950: inst = 32'hc4048c2;
      9951: inst = 32'h8220000;
      9952: inst = 32'h10408000;
      9953: inst = 32'hc4048c3;
      9954: inst = 32'h8220000;
      9955: inst = 32'h10408000;
      9956: inst = 32'hc4048fc;
      9957: inst = 32'h8220000;
      9958: inst = 32'h10408000;
      9959: inst = 32'hc4048fd;
      9960: inst = 32'h8220000;
      9961: inst = 32'h10408000;
      9962: inst = 32'hc4048fe;
      9963: inst = 32'h8220000;
      9964: inst = 32'h10408000;
      9965: inst = 32'hc4048ff;
      9966: inst = 32'h8220000;
      9967: inst = 32'h10408000;
      9968: inst = 32'hc404900;
      9969: inst = 32'h8220000;
      9970: inst = 32'h10408000;
      9971: inst = 32'hc404901;
      9972: inst = 32'h8220000;
      9973: inst = 32'h10408000;
      9974: inst = 32'hc404902;
      9975: inst = 32'h8220000;
      9976: inst = 32'h10408000;
      9977: inst = 32'hc404903;
      9978: inst = 32'h8220000;
      9979: inst = 32'h10408000;
      9980: inst = 32'hc404904;
      9981: inst = 32'h8220000;
      9982: inst = 32'h10408000;
      9983: inst = 32'hc404905;
      9984: inst = 32'h8220000;
      9985: inst = 32'h10408000;
      9986: inst = 32'hc404906;
      9987: inst = 32'h8220000;
      9988: inst = 32'h10408000;
      9989: inst = 32'hc404907;
      9990: inst = 32'h8220000;
      9991: inst = 32'h10408000;
      9992: inst = 32'hc404908;
      9993: inst = 32'h8220000;
      9994: inst = 32'h10408000;
      9995: inst = 32'hc404909;
      9996: inst = 32'h8220000;
      9997: inst = 32'h10408000;
      9998: inst = 32'hc40490a;
      9999: inst = 32'h8220000;
      10000: inst = 32'h10408000;
      10001: inst = 32'hc40490b;
      10002: inst = 32'h8220000;
      10003: inst = 32'h10408000;
      10004: inst = 32'hc40490c;
      10005: inst = 32'h8220000;
      10006: inst = 32'h10408000;
      10007: inst = 32'hc40490d;
      10008: inst = 32'h8220000;
      10009: inst = 32'h10408000;
      10010: inst = 32'hc40490e;
      10011: inst = 32'h8220000;
      10012: inst = 32'h10408000;
      10013: inst = 32'hc40490f;
      10014: inst = 32'h8220000;
      10015: inst = 32'h10408000;
      10016: inst = 32'hc404910;
      10017: inst = 32'h8220000;
      10018: inst = 32'h10408000;
      10019: inst = 32'hc404911;
      10020: inst = 32'h8220000;
      10021: inst = 32'h10408000;
      10022: inst = 32'hc404912;
      10023: inst = 32'h8220000;
      10024: inst = 32'h10408000;
      10025: inst = 32'hc404913;
      10026: inst = 32'h8220000;
      10027: inst = 32'h10408000;
      10028: inst = 32'hc404914;
      10029: inst = 32'h8220000;
      10030: inst = 32'h10408000;
      10031: inst = 32'hc404915;
      10032: inst = 32'h8220000;
      10033: inst = 32'h10408000;
      10034: inst = 32'hc404916;
      10035: inst = 32'h8220000;
      10036: inst = 32'h10408000;
      10037: inst = 32'hc404917;
      10038: inst = 32'h8220000;
      10039: inst = 32'h10408000;
      10040: inst = 32'hc404918;
      10041: inst = 32'h8220000;
      10042: inst = 32'h10408000;
      10043: inst = 32'hc404919;
      10044: inst = 32'h8220000;
      10045: inst = 32'h10408000;
      10046: inst = 32'hc40491a;
      10047: inst = 32'h8220000;
      10048: inst = 32'h10408000;
      10049: inst = 32'hc40491b;
      10050: inst = 32'h8220000;
      10051: inst = 32'h10408000;
      10052: inst = 32'hc40491c;
      10053: inst = 32'h8220000;
      10054: inst = 32'h10408000;
      10055: inst = 32'hc40491d;
      10056: inst = 32'h8220000;
      10057: inst = 32'h10408000;
      10058: inst = 32'hc40491e;
      10059: inst = 32'h8220000;
      10060: inst = 32'h10408000;
      10061: inst = 32'hc40491f;
      10062: inst = 32'h8220000;
      10063: inst = 32'h10408000;
      10064: inst = 32'hc404920;
      10065: inst = 32'h8220000;
      10066: inst = 32'h10408000;
      10067: inst = 32'hc404921;
      10068: inst = 32'h8220000;
      10069: inst = 32'h10408000;
      10070: inst = 32'hc404922;
      10071: inst = 32'h8220000;
      10072: inst = 32'h10408000;
      10073: inst = 32'hc404923;
      10074: inst = 32'h8220000;
      10075: inst = 32'h10408000;
      10076: inst = 32'hc40495c;
      10077: inst = 32'h8220000;
      10078: inst = 32'h10408000;
      10079: inst = 32'hc40495d;
      10080: inst = 32'h8220000;
      10081: inst = 32'h10408000;
      10082: inst = 32'hc40495e;
      10083: inst = 32'h8220000;
      10084: inst = 32'h10408000;
      10085: inst = 32'hc40495f;
      10086: inst = 32'h8220000;
      10087: inst = 32'h10408000;
      10088: inst = 32'hc404960;
      10089: inst = 32'h8220000;
      10090: inst = 32'h10408000;
      10091: inst = 32'hc404961;
      10092: inst = 32'h8220000;
      10093: inst = 32'h10408000;
      10094: inst = 32'hc404962;
      10095: inst = 32'h8220000;
      10096: inst = 32'h10408000;
      10097: inst = 32'hc404963;
      10098: inst = 32'h8220000;
      10099: inst = 32'h10408000;
      10100: inst = 32'hc404964;
      10101: inst = 32'h8220000;
      10102: inst = 32'h10408000;
      10103: inst = 32'hc404965;
      10104: inst = 32'h8220000;
      10105: inst = 32'h10408000;
      10106: inst = 32'hc404966;
      10107: inst = 32'h8220000;
      10108: inst = 32'h10408000;
      10109: inst = 32'hc404967;
      10110: inst = 32'h8220000;
      10111: inst = 32'h10408000;
      10112: inst = 32'hc404968;
      10113: inst = 32'h8220000;
      10114: inst = 32'h10408000;
      10115: inst = 32'hc404969;
      10116: inst = 32'h8220000;
      10117: inst = 32'h10408000;
      10118: inst = 32'hc40496a;
      10119: inst = 32'h8220000;
      10120: inst = 32'h10408000;
      10121: inst = 32'hc40496b;
      10122: inst = 32'h8220000;
      10123: inst = 32'h10408000;
      10124: inst = 32'hc40496c;
      10125: inst = 32'h8220000;
      10126: inst = 32'h10408000;
      10127: inst = 32'hc40496d;
      10128: inst = 32'h8220000;
      10129: inst = 32'h10408000;
      10130: inst = 32'hc40496e;
      10131: inst = 32'h8220000;
      10132: inst = 32'h10408000;
      10133: inst = 32'hc40496f;
      10134: inst = 32'h8220000;
      10135: inst = 32'h10408000;
      10136: inst = 32'hc404970;
      10137: inst = 32'h8220000;
      10138: inst = 32'h10408000;
      10139: inst = 32'hc404971;
      10140: inst = 32'h8220000;
      10141: inst = 32'h10408000;
      10142: inst = 32'hc404972;
      10143: inst = 32'h8220000;
      10144: inst = 32'h10408000;
      10145: inst = 32'hc404973;
      10146: inst = 32'h8220000;
      10147: inst = 32'h10408000;
      10148: inst = 32'hc404974;
      10149: inst = 32'h8220000;
      10150: inst = 32'h10408000;
      10151: inst = 32'hc404975;
      10152: inst = 32'h8220000;
      10153: inst = 32'h10408000;
      10154: inst = 32'hc404976;
      10155: inst = 32'h8220000;
      10156: inst = 32'h10408000;
      10157: inst = 32'hc404977;
      10158: inst = 32'h8220000;
      10159: inst = 32'h10408000;
      10160: inst = 32'hc404978;
      10161: inst = 32'h8220000;
      10162: inst = 32'h10408000;
      10163: inst = 32'hc404979;
      10164: inst = 32'h8220000;
      10165: inst = 32'h10408000;
      10166: inst = 32'hc40497a;
      10167: inst = 32'h8220000;
      10168: inst = 32'h10408000;
      10169: inst = 32'hc40497b;
      10170: inst = 32'h8220000;
      10171: inst = 32'h10408000;
      10172: inst = 32'hc40497c;
      10173: inst = 32'h8220000;
      10174: inst = 32'h10408000;
      10175: inst = 32'hc40497d;
      10176: inst = 32'h8220000;
      10177: inst = 32'h10408000;
      10178: inst = 32'hc40497e;
      10179: inst = 32'h8220000;
      10180: inst = 32'h10408000;
      10181: inst = 32'hc40497f;
      10182: inst = 32'h8220000;
      10183: inst = 32'h10408000;
      10184: inst = 32'hc404980;
      10185: inst = 32'h8220000;
      10186: inst = 32'h10408000;
      10187: inst = 32'hc404981;
      10188: inst = 32'h8220000;
      10189: inst = 32'h10408000;
      10190: inst = 32'hc404982;
      10191: inst = 32'h8220000;
      10192: inst = 32'h10408000;
      10193: inst = 32'hc404983;
      10194: inst = 32'h8220000;
      10195: inst = 32'h10408000;
      10196: inst = 32'hc404992;
      10197: inst = 32'h8220000;
      10198: inst = 32'h10408000;
      10199: inst = 32'hc4049bc;
      10200: inst = 32'h8220000;
      10201: inst = 32'h10408000;
      10202: inst = 32'hc4049bd;
      10203: inst = 32'h8220000;
      10204: inst = 32'h10408000;
      10205: inst = 32'hc4049be;
      10206: inst = 32'h8220000;
      10207: inst = 32'h10408000;
      10208: inst = 32'hc4049bf;
      10209: inst = 32'h8220000;
      10210: inst = 32'h10408000;
      10211: inst = 32'hc4049c0;
      10212: inst = 32'h8220000;
      10213: inst = 32'h10408000;
      10214: inst = 32'hc4049c1;
      10215: inst = 32'h8220000;
      10216: inst = 32'h10408000;
      10217: inst = 32'hc4049c2;
      10218: inst = 32'h8220000;
      10219: inst = 32'h10408000;
      10220: inst = 32'hc4049c3;
      10221: inst = 32'h8220000;
      10222: inst = 32'h10408000;
      10223: inst = 32'hc4049c4;
      10224: inst = 32'h8220000;
      10225: inst = 32'h10408000;
      10226: inst = 32'hc4049c5;
      10227: inst = 32'h8220000;
      10228: inst = 32'h10408000;
      10229: inst = 32'hc4049c6;
      10230: inst = 32'h8220000;
      10231: inst = 32'h10408000;
      10232: inst = 32'hc4049c7;
      10233: inst = 32'h8220000;
      10234: inst = 32'h10408000;
      10235: inst = 32'hc4049c8;
      10236: inst = 32'h8220000;
      10237: inst = 32'h10408000;
      10238: inst = 32'hc4049c9;
      10239: inst = 32'h8220000;
      10240: inst = 32'h10408000;
      10241: inst = 32'hc4049ca;
      10242: inst = 32'h8220000;
      10243: inst = 32'h10408000;
      10244: inst = 32'hc4049cb;
      10245: inst = 32'h8220000;
      10246: inst = 32'h10408000;
      10247: inst = 32'hc4049cc;
      10248: inst = 32'h8220000;
      10249: inst = 32'h10408000;
      10250: inst = 32'hc4049cd;
      10251: inst = 32'h8220000;
      10252: inst = 32'h10408000;
      10253: inst = 32'hc4049ce;
      10254: inst = 32'h8220000;
      10255: inst = 32'h10408000;
      10256: inst = 32'hc4049cf;
      10257: inst = 32'h8220000;
      10258: inst = 32'h10408000;
      10259: inst = 32'hc4049d0;
      10260: inst = 32'h8220000;
      10261: inst = 32'h10408000;
      10262: inst = 32'hc4049d1;
      10263: inst = 32'h8220000;
      10264: inst = 32'h10408000;
      10265: inst = 32'hc4049d2;
      10266: inst = 32'h8220000;
      10267: inst = 32'h10408000;
      10268: inst = 32'hc4049d3;
      10269: inst = 32'h8220000;
      10270: inst = 32'h10408000;
      10271: inst = 32'hc4049d4;
      10272: inst = 32'h8220000;
      10273: inst = 32'h10408000;
      10274: inst = 32'hc4049d5;
      10275: inst = 32'h8220000;
      10276: inst = 32'h10408000;
      10277: inst = 32'hc4049d6;
      10278: inst = 32'h8220000;
      10279: inst = 32'h10408000;
      10280: inst = 32'hc4049d7;
      10281: inst = 32'h8220000;
      10282: inst = 32'h10408000;
      10283: inst = 32'hc4049d8;
      10284: inst = 32'h8220000;
      10285: inst = 32'h10408000;
      10286: inst = 32'hc4049d9;
      10287: inst = 32'h8220000;
      10288: inst = 32'h10408000;
      10289: inst = 32'hc4049da;
      10290: inst = 32'h8220000;
      10291: inst = 32'h10408000;
      10292: inst = 32'hc4049db;
      10293: inst = 32'h8220000;
      10294: inst = 32'h10408000;
      10295: inst = 32'hc4049dc;
      10296: inst = 32'h8220000;
      10297: inst = 32'h10408000;
      10298: inst = 32'hc4049dd;
      10299: inst = 32'h8220000;
      10300: inst = 32'h10408000;
      10301: inst = 32'hc4049de;
      10302: inst = 32'h8220000;
      10303: inst = 32'h10408000;
      10304: inst = 32'hc4049df;
      10305: inst = 32'h8220000;
      10306: inst = 32'h10408000;
      10307: inst = 32'hc4049e0;
      10308: inst = 32'h8220000;
      10309: inst = 32'h10408000;
      10310: inst = 32'hc4049e1;
      10311: inst = 32'h8220000;
      10312: inst = 32'h10408000;
      10313: inst = 32'hc4049e2;
      10314: inst = 32'h8220000;
      10315: inst = 32'h10408000;
      10316: inst = 32'hc4049e3;
      10317: inst = 32'h8220000;
      10318: inst = 32'h10408000;
      10319: inst = 32'hc4049f2;
      10320: inst = 32'h8220000;
      10321: inst = 32'h10408000;
      10322: inst = 32'hc404a1c;
      10323: inst = 32'h8220000;
      10324: inst = 32'h10408000;
      10325: inst = 32'hc404a1d;
      10326: inst = 32'h8220000;
      10327: inst = 32'h10408000;
      10328: inst = 32'hc404a1e;
      10329: inst = 32'h8220000;
      10330: inst = 32'h10408000;
      10331: inst = 32'hc404a1f;
      10332: inst = 32'h8220000;
      10333: inst = 32'h10408000;
      10334: inst = 32'hc404a20;
      10335: inst = 32'h8220000;
      10336: inst = 32'h10408000;
      10337: inst = 32'hc404a21;
      10338: inst = 32'h8220000;
      10339: inst = 32'h10408000;
      10340: inst = 32'hc404a22;
      10341: inst = 32'h8220000;
      10342: inst = 32'h10408000;
      10343: inst = 32'hc404a23;
      10344: inst = 32'h8220000;
      10345: inst = 32'h10408000;
      10346: inst = 32'hc404a24;
      10347: inst = 32'h8220000;
      10348: inst = 32'h10408000;
      10349: inst = 32'hc404a25;
      10350: inst = 32'h8220000;
      10351: inst = 32'h10408000;
      10352: inst = 32'hc404a26;
      10353: inst = 32'h8220000;
      10354: inst = 32'h10408000;
      10355: inst = 32'hc404a27;
      10356: inst = 32'h8220000;
      10357: inst = 32'h10408000;
      10358: inst = 32'hc404a28;
      10359: inst = 32'h8220000;
      10360: inst = 32'h10408000;
      10361: inst = 32'hc404a29;
      10362: inst = 32'h8220000;
      10363: inst = 32'h10408000;
      10364: inst = 32'hc404a2a;
      10365: inst = 32'h8220000;
      10366: inst = 32'h10408000;
      10367: inst = 32'hc404a2b;
      10368: inst = 32'h8220000;
      10369: inst = 32'h10408000;
      10370: inst = 32'hc404a2c;
      10371: inst = 32'h8220000;
      10372: inst = 32'h10408000;
      10373: inst = 32'hc404a2d;
      10374: inst = 32'h8220000;
      10375: inst = 32'h10408000;
      10376: inst = 32'hc404a2e;
      10377: inst = 32'h8220000;
      10378: inst = 32'h10408000;
      10379: inst = 32'hc404a2f;
      10380: inst = 32'h8220000;
      10381: inst = 32'h10408000;
      10382: inst = 32'hc404a30;
      10383: inst = 32'h8220000;
      10384: inst = 32'h10408000;
      10385: inst = 32'hc404a31;
      10386: inst = 32'h8220000;
      10387: inst = 32'h10408000;
      10388: inst = 32'hc404a32;
      10389: inst = 32'h8220000;
      10390: inst = 32'h10408000;
      10391: inst = 32'hc404a33;
      10392: inst = 32'h8220000;
      10393: inst = 32'h10408000;
      10394: inst = 32'hc404a34;
      10395: inst = 32'h8220000;
      10396: inst = 32'h10408000;
      10397: inst = 32'hc404a35;
      10398: inst = 32'h8220000;
      10399: inst = 32'h10408000;
      10400: inst = 32'hc404a36;
      10401: inst = 32'h8220000;
      10402: inst = 32'h10408000;
      10403: inst = 32'hc404a37;
      10404: inst = 32'h8220000;
      10405: inst = 32'h10408000;
      10406: inst = 32'hc404a38;
      10407: inst = 32'h8220000;
      10408: inst = 32'h10408000;
      10409: inst = 32'hc404a39;
      10410: inst = 32'h8220000;
      10411: inst = 32'h10408000;
      10412: inst = 32'hc404a3a;
      10413: inst = 32'h8220000;
      10414: inst = 32'h10408000;
      10415: inst = 32'hc404a3b;
      10416: inst = 32'h8220000;
      10417: inst = 32'h10408000;
      10418: inst = 32'hc404a3c;
      10419: inst = 32'h8220000;
      10420: inst = 32'h10408000;
      10421: inst = 32'hc404a3d;
      10422: inst = 32'h8220000;
      10423: inst = 32'h10408000;
      10424: inst = 32'hc404a3e;
      10425: inst = 32'h8220000;
      10426: inst = 32'h10408000;
      10427: inst = 32'hc404a3f;
      10428: inst = 32'h8220000;
      10429: inst = 32'h10408000;
      10430: inst = 32'hc404a40;
      10431: inst = 32'h8220000;
      10432: inst = 32'h10408000;
      10433: inst = 32'hc404a41;
      10434: inst = 32'h8220000;
      10435: inst = 32'h10408000;
      10436: inst = 32'hc404a42;
      10437: inst = 32'h8220000;
      10438: inst = 32'h10408000;
      10439: inst = 32'hc404a43;
      10440: inst = 32'h8220000;
      10441: inst = 32'h10408000;
      10442: inst = 32'hc404a52;
      10443: inst = 32'h8220000;
      10444: inst = 32'h10408000;
      10445: inst = 32'hc404a7c;
      10446: inst = 32'h8220000;
      10447: inst = 32'h10408000;
      10448: inst = 32'hc404a7d;
      10449: inst = 32'h8220000;
      10450: inst = 32'h10408000;
      10451: inst = 32'hc404a7e;
      10452: inst = 32'h8220000;
      10453: inst = 32'h10408000;
      10454: inst = 32'hc404a7f;
      10455: inst = 32'h8220000;
      10456: inst = 32'h10408000;
      10457: inst = 32'hc404a80;
      10458: inst = 32'h8220000;
      10459: inst = 32'h10408000;
      10460: inst = 32'hc404a81;
      10461: inst = 32'h8220000;
      10462: inst = 32'h10408000;
      10463: inst = 32'hc404a82;
      10464: inst = 32'h8220000;
      10465: inst = 32'h10408000;
      10466: inst = 32'hc404a83;
      10467: inst = 32'h8220000;
      10468: inst = 32'h10408000;
      10469: inst = 32'hc404a84;
      10470: inst = 32'h8220000;
      10471: inst = 32'h10408000;
      10472: inst = 32'hc404a85;
      10473: inst = 32'h8220000;
      10474: inst = 32'h10408000;
      10475: inst = 32'hc404a86;
      10476: inst = 32'h8220000;
      10477: inst = 32'h10408000;
      10478: inst = 32'hc404a87;
      10479: inst = 32'h8220000;
      10480: inst = 32'h10408000;
      10481: inst = 32'hc404a88;
      10482: inst = 32'h8220000;
      10483: inst = 32'h10408000;
      10484: inst = 32'hc404a89;
      10485: inst = 32'h8220000;
      10486: inst = 32'h10408000;
      10487: inst = 32'hc404a8a;
      10488: inst = 32'h8220000;
      10489: inst = 32'h10408000;
      10490: inst = 32'hc404a8b;
      10491: inst = 32'h8220000;
      10492: inst = 32'h10408000;
      10493: inst = 32'hc404a8c;
      10494: inst = 32'h8220000;
      10495: inst = 32'h10408000;
      10496: inst = 32'hc404a8d;
      10497: inst = 32'h8220000;
      10498: inst = 32'h10408000;
      10499: inst = 32'hc404a8e;
      10500: inst = 32'h8220000;
      10501: inst = 32'h10408000;
      10502: inst = 32'hc404a8f;
      10503: inst = 32'h8220000;
      10504: inst = 32'h10408000;
      10505: inst = 32'hc404a90;
      10506: inst = 32'h8220000;
      10507: inst = 32'h10408000;
      10508: inst = 32'hc404a91;
      10509: inst = 32'h8220000;
      10510: inst = 32'h10408000;
      10511: inst = 32'hc404a92;
      10512: inst = 32'h8220000;
      10513: inst = 32'h10408000;
      10514: inst = 32'hc404a93;
      10515: inst = 32'h8220000;
      10516: inst = 32'h10408000;
      10517: inst = 32'hc404a94;
      10518: inst = 32'h8220000;
      10519: inst = 32'h10408000;
      10520: inst = 32'hc404a95;
      10521: inst = 32'h8220000;
      10522: inst = 32'h10408000;
      10523: inst = 32'hc404a96;
      10524: inst = 32'h8220000;
      10525: inst = 32'h10408000;
      10526: inst = 32'hc404a97;
      10527: inst = 32'h8220000;
      10528: inst = 32'h10408000;
      10529: inst = 32'hc404a98;
      10530: inst = 32'h8220000;
      10531: inst = 32'h10408000;
      10532: inst = 32'hc404a99;
      10533: inst = 32'h8220000;
      10534: inst = 32'h10408000;
      10535: inst = 32'hc404a9a;
      10536: inst = 32'h8220000;
      10537: inst = 32'h10408000;
      10538: inst = 32'hc404a9b;
      10539: inst = 32'h8220000;
      10540: inst = 32'h10408000;
      10541: inst = 32'hc404a9c;
      10542: inst = 32'h8220000;
      10543: inst = 32'h10408000;
      10544: inst = 32'hc404a9d;
      10545: inst = 32'h8220000;
      10546: inst = 32'h10408000;
      10547: inst = 32'hc404a9e;
      10548: inst = 32'h8220000;
      10549: inst = 32'h10408000;
      10550: inst = 32'hc404a9f;
      10551: inst = 32'h8220000;
      10552: inst = 32'h10408000;
      10553: inst = 32'hc404aa0;
      10554: inst = 32'h8220000;
      10555: inst = 32'h10408000;
      10556: inst = 32'hc404aa1;
      10557: inst = 32'h8220000;
      10558: inst = 32'h10408000;
      10559: inst = 32'hc404aa2;
      10560: inst = 32'h8220000;
      10561: inst = 32'h10408000;
      10562: inst = 32'hc404aa3;
      10563: inst = 32'h8220000;
      10564: inst = 32'h10408000;
      10565: inst = 32'hc404ab4;
      10566: inst = 32'h8220000;
      10567: inst = 32'h10408000;
      10568: inst = 32'hc404adc;
      10569: inst = 32'h8220000;
      10570: inst = 32'h10408000;
      10571: inst = 32'hc404add;
      10572: inst = 32'h8220000;
      10573: inst = 32'h10408000;
      10574: inst = 32'hc404ade;
      10575: inst = 32'h8220000;
      10576: inst = 32'h10408000;
      10577: inst = 32'hc404adf;
      10578: inst = 32'h8220000;
      10579: inst = 32'h10408000;
      10580: inst = 32'hc404ae0;
      10581: inst = 32'h8220000;
      10582: inst = 32'h10408000;
      10583: inst = 32'hc404ae1;
      10584: inst = 32'h8220000;
      10585: inst = 32'h10408000;
      10586: inst = 32'hc404ae2;
      10587: inst = 32'h8220000;
      10588: inst = 32'h10408000;
      10589: inst = 32'hc404ae3;
      10590: inst = 32'h8220000;
      10591: inst = 32'h10408000;
      10592: inst = 32'hc404ae4;
      10593: inst = 32'h8220000;
      10594: inst = 32'h10408000;
      10595: inst = 32'hc404ae5;
      10596: inst = 32'h8220000;
      10597: inst = 32'h10408000;
      10598: inst = 32'hc404ae6;
      10599: inst = 32'h8220000;
      10600: inst = 32'h10408000;
      10601: inst = 32'hc404ae7;
      10602: inst = 32'h8220000;
      10603: inst = 32'h10408000;
      10604: inst = 32'hc404ae8;
      10605: inst = 32'h8220000;
      10606: inst = 32'h10408000;
      10607: inst = 32'hc404ae9;
      10608: inst = 32'h8220000;
      10609: inst = 32'h10408000;
      10610: inst = 32'hc404aea;
      10611: inst = 32'h8220000;
      10612: inst = 32'h10408000;
      10613: inst = 32'hc404aeb;
      10614: inst = 32'h8220000;
      10615: inst = 32'h10408000;
      10616: inst = 32'hc404aec;
      10617: inst = 32'h8220000;
      10618: inst = 32'h10408000;
      10619: inst = 32'hc404aed;
      10620: inst = 32'h8220000;
      10621: inst = 32'h10408000;
      10622: inst = 32'hc404aee;
      10623: inst = 32'h8220000;
      10624: inst = 32'h10408000;
      10625: inst = 32'hc404aef;
      10626: inst = 32'h8220000;
      10627: inst = 32'h10408000;
      10628: inst = 32'hc404af0;
      10629: inst = 32'h8220000;
      10630: inst = 32'h10408000;
      10631: inst = 32'hc404af1;
      10632: inst = 32'h8220000;
      10633: inst = 32'h10408000;
      10634: inst = 32'hc404af2;
      10635: inst = 32'h8220000;
      10636: inst = 32'h10408000;
      10637: inst = 32'hc404af3;
      10638: inst = 32'h8220000;
      10639: inst = 32'h10408000;
      10640: inst = 32'hc404af4;
      10641: inst = 32'h8220000;
      10642: inst = 32'h10408000;
      10643: inst = 32'hc404af5;
      10644: inst = 32'h8220000;
      10645: inst = 32'h10408000;
      10646: inst = 32'hc404af6;
      10647: inst = 32'h8220000;
      10648: inst = 32'h10408000;
      10649: inst = 32'hc404af7;
      10650: inst = 32'h8220000;
      10651: inst = 32'h10408000;
      10652: inst = 32'hc404af8;
      10653: inst = 32'h8220000;
      10654: inst = 32'h10408000;
      10655: inst = 32'hc404af9;
      10656: inst = 32'h8220000;
      10657: inst = 32'h10408000;
      10658: inst = 32'hc404afa;
      10659: inst = 32'h8220000;
      10660: inst = 32'h10408000;
      10661: inst = 32'hc404afb;
      10662: inst = 32'h8220000;
      10663: inst = 32'h10408000;
      10664: inst = 32'hc404afc;
      10665: inst = 32'h8220000;
      10666: inst = 32'h10408000;
      10667: inst = 32'hc404afd;
      10668: inst = 32'h8220000;
      10669: inst = 32'h10408000;
      10670: inst = 32'hc404afe;
      10671: inst = 32'h8220000;
      10672: inst = 32'h10408000;
      10673: inst = 32'hc404aff;
      10674: inst = 32'h8220000;
      10675: inst = 32'h10408000;
      10676: inst = 32'hc404b00;
      10677: inst = 32'h8220000;
      10678: inst = 32'h10408000;
      10679: inst = 32'hc404b01;
      10680: inst = 32'h8220000;
      10681: inst = 32'h10408000;
      10682: inst = 32'hc404b02;
      10683: inst = 32'h8220000;
      10684: inst = 32'h10408000;
      10685: inst = 32'hc404b03;
      10686: inst = 32'h8220000;
      10687: inst = 32'h10408000;
      10688: inst = 32'hc404b14;
      10689: inst = 32'h8220000;
      10690: inst = 32'h10408000;
      10691: inst = 32'hc404b3c;
      10692: inst = 32'h8220000;
      10693: inst = 32'h10408000;
      10694: inst = 32'hc404b3d;
      10695: inst = 32'h8220000;
      10696: inst = 32'h10408000;
      10697: inst = 32'hc404b3e;
      10698: inst = 32'h8220000;
      10699: inst = 32'h10408000;
      10700: inst = 32'hc404b3f;
      10701: inst = 32'h8220000;
      10702: inst = 32'h10408000;
      10703: inst = 32'hc404b40;
      10704: inst = 32'h8220000;
      10705: inst = 32'h10408000;
      10706: inst = 32'hc404b41;
      10707: inst = 32'h8220000;
      10708: inst = 32'h10408000;
      10709: inst = 32'hc404b42;
      10710: inst = 32'h8220000;
      10711: inst = 32'h10408000;
      10712: inst = 32'hc404b43;
      10713: inst = 32'h8220000;
      10714: inst = 32'h10408000;
      10715: inst = 32'hc404b44;
      10716: inst = 32'h8220000;
      10717: inst = 32'h10408000;
      10718: inst = 32'hc404b45;
      10719: inst = 32'h8220000;
      10720: inst = 32'h10408000;
      10721: inst = 32'hc404b46;
      10722: inst = 32'h8220000;
      10723: inst = 32'h10408000;
      10724: inst = 32'hc404b47;
      10725: inst = 32'h8220000;
      10726: inst = 32'h10408000;
      10727: inst = 32'hc404b48;
      10728: inst = 32'h8220000;
      10729: inst = 32'h10408000;
      10730: inst = 32'hc404b49;
      10731: inst = 32'h8220000;
      10732: inst = 32'h10408000;
      10733: inst = 32'hc404b4a;
      10734: inst = 32'h8220000;
      10735: inst = 32'h10408000;
      10736: inst = 32'hc404b4b;
      10737: inst = 32'h8220000;
      10738: inst = 32'h10408000;
      10739: inst = 32'hc404b4c;
      10740: inst = 32'h8220000;
      10741: inst = 32'h10408000;
      10742: inst = 32'hc404b4d;
      10743: inst = 32'h8220000;
      10744: inst = 32'h10408000;
      10745: inst = 32'hc404b4e;
      10746: inst = 32'h8220000;
      10747: inst = 32'h10408000;
      10748: inst = 32'hc404b4f;
      10749: inst = 32'h8220000;
      10750: inst = 32'h10408000;
      10751: inst = 32'hc404b50;
      10752: inst = 32'h8220000;
      10753: inst = 32'h10408000;
      10754: inst = 32'hc404b51;
      10755: inst = 32'h8220000;
      10756: inst = 32'h10408000;
      10757: inst = 32'hc404b52;
      10758: inst = 32'h8220000;
      10759: inst = 32'h10408000;
      10760: inst = 32'hc404b53;
      10761: inst = 32'h8220000;
      10762: inst = 32'h10408000;
      10763: inst = 32'hc404b54;
      10764: inst = 32'h8220000;
      10765: inst = 32'h10408000;
      10766: inst = 32'hc404b55;
      10767: inst = 32'h8220000;
      10768: inst = 32'h10408000;
      10769: inst = 32'hc404b56;
      10770: inst = 32'h8220000;
      10771: inst = 32'h10408000;
      10772: inst = 32'hc404b57;
      10773: inst = 32'h8220000;
      10774: inst = 32'h10408000;
      10775: inst = 32'hc404b58;
      10776: inst = 32'h8220000;
      10777: inst = 32'h10408000;
      10778: inst = 32'hc404b59;
      10779: inst = 32'h8220000;
      10780: inst = 32'h10408000;
      10781: inst = 32'hc404b5a;
      10782: inst = 32'h8220000;
      10783: inst = 32'h10408000;
      10784: inst = 32'hc404b5b;
      10785: inst = 32'h8220000;
      10786: inst = 32'h10408000;
      10787: inst = 32'hc404b5c;
      10788: inst = 32'h8220000;
      10789: inst = 32'h10408000;
      10790: inst = 32'hc404b5d;
      10791: inst = 32'h8220000;
      10792: inst = 32'h10408000;
      10793: inst = 32'hc404b5e;
      10794: inst = 32'h8220000;
      10795: inst = 32'h10408000;
      10796: inst = 32'hc404b5f;
      10797: inst = 32'h8220000;
      10798: inst = 32'h10408000;
      10799: inst = 32'hc404b60;
      10800: inst = 32'h8220000;
      10801: inst = 32'h10408000;
      10802: inst = 32'hc404b61;
      10803: inst = 32'h8220000;
      10804: inst = 32'h10408000;
      10805: inst = 32'hc404b62;
      10806: inst = 32'h8220000;
      10807: inst = 32'h10408000;
      10808: inst = 32'hc404b63;
      10809: inst = 32'h8220000;
      10810: inst = 32'h10408000;
      10811: inst = 32'hc404b9c;
      10812: inst = 32'h8220000;
      10813: inst = 32'h10408000;
      10814: inst = 32'hc404b9d;
      10815: inst = 32'h8220000;
      10816: inst = 32'h10408000;
      10817: inst = 32'hc404b9e;
      10818: inst = 32'h8220000;
      10819: inst = 32'h10408000;
      10820: inst = 32'hc404b9f;
      10821: inst = 32'h8220000;
      10822: inst = 32'h10408000;
      10823: inst = 32'hc404ba0;
      10824: inst = 32'h8220000;
      10825: inst = 32'h10408000;
      10826: inst = 32'hc404ba1;
      10827: inst = 32'h8220000;
      10828: inst = 32'h10408000;
      10829: inst = 32'hc404ba2;
      10830: inst = 32'h8220000;
      10831: inst = 32'h10408000;
      10832: inst = 32'hc404ba3;
      10833: inst = 32'h8220000;
      10834: inst = 32'h10408000;
      10835: inst = 32'hc404ba4;
      10836: inst = 32'h8220000;
      10837: inst = 32'h10408000;
      10838: inst = 32'hc404ba5;
      10839: inst = 32'h8220000;
      10840: inst = 32'h10408000;
      10841: inst = 32'hc404ba6;
      10842: inst = 32'h8220000;
      10843: inst = 32'h10408000;
      10844: inst = 32'hc404ba7;
      10845: inst = 32'h8220000;
      10846: inst = 32'h10408000;
      10847: inst = 32'hc404ba8;
      10848: inst = 32'h8220000;
      10849: inst = 32'h10408000;
      10850: inst = 32'hc404ba9;
      10851: inst = 32'h8220000;
      10852: inst = 32'h10408000;
      10853: inst = 32'hc404baa;
      10854: inst = 32'h8220000;
      10855: inst = 32'h10408000;
      10856: inst = 32'hc404bab;
      10857: inst = 32'h8220000;
      10858: inst = 32'h10408000;
      10859: inst = 32'hc404bac;
      10860: inst = 32'h8220000;
      10861: inst = 32'h10408000;
      10862: inst = 32'hc404bad;
      10863: inst = 32'h8220000;
      10864: inst = 32'h10408000;
      10865: inst = 32'hc404bae;
      10866: inst = 32'h8220000;
      10867: inst = 32'h10408000;
      10868: inst = 32'hc404baf;
      10869: inst = 32'h8220000;
      10870: inst = 32'h10408000;
      10871: inst = 32'hc404bb0;
      10872: inst = 32'h8220000;
      10873: inst = 32'h10408000;
      10874: inst = 32'hc404bb1;
      10875: inst = 32'h8220000;
      10876: inst = 32'h10408000;
      10877: inst = 32'hc404bb2;
      10878: inst = 32'h8220000;
      10879: inst = 32'h10408000;
      10880: inst = 32'hc404bb3;
      10881: inst = 32'h8220000;
      10882: inst = 32'h10408000;
      10883: inst = 32'hc404bb4;
      10884: inst = 32'h8220000;
      10885: inst = 32'h10408000;
      10886: inst = 32'hc404bb5;
      10887: inst = 32'h8220000;
      10888: inst = 32'h10408000;
      10889: inst = 32'hc404bb6;
      10890: inst = 32'h8220000;
      10891: inst = 32'h10408000;
      10892: inst = 32'hc404bb7;
      10893: inst = 32'h8220000;
      10894: inst = 32'h10408000;
      10895: inst = 32'hc404bb8;
      10896: inst = 32'h8220000;
      10897: inst = 32'h10408000;
      10898: inst = 32'hc404bb9;
      10899: inst = 32'h8220000;
      10900: inst = 32'h10408000;
      10901: inst = 32'hc404bba;
      10902: inst = 32'h8220000;
      10903: inst = 32'h10408000;
      10904: inst = 32'hc404bbb;
      10905: inst = 32'h8220000;
      10906: inst = 32'h10408000;
      10907: inst = 32'hc404bbc;
      10908: inst = 32'h8220000;
      10909: inst = 32'h10408000;
      10910: inst = 32'hc404bbd;
      10911: inst = 32'h8220000;
      10912: inst = 32'h10408000;
      10913: inst = 32'hc404bbe;
      10914: inst = 32'h8220000;
      10915: inst = 32'h10408000;
      10916: inst = 32'hc404bbf;
      10917: inst = 32'h8220000;
      10918: inst = 32'h10408000;
      10919: inst = 32'hc404bc0;
      10920: inst = 32'h8220000;
      10921: inst = 32'h10408000;
      10922: inst = 32'hc404bc1;
      10923: inst = 32'h8220000;
      10924: inst = 32'h10408000;
      10925: inst = 32'hc404bc2;
      10926: inst = 32'h8220000;
      10927: inst = 32'h10408000;
      10928: inst = 32'hc404bc3;
      10929: inst = 32'h8220000;
      10930: inst = 32'hc20ee75;
      10931: inst = 32'h10408000;
      10932: inst = 32'hc4042ea;
      10933: inst = 32'h8220000;
      10934: inst = 32'h10408000;
      10935: inst = 32'hc4043a7;
      10936: inst = 32'h8220000;
      10937: inst = 32'hc20d42c;
      10938: inst = 32'h10408000;
      10939: inst = 32'hc4042eb;
      10940: inst = 32'h8220000;
      10941: inst = 32'h10408000;
      10942: inst = 32'hc4042ec;
      10943: inst = 32'h8220000;
      10944: inst = 32'h10408000;
      10945: inst = 32'hc4043a8;
      10946: inst = 32'h8220000;
      10947: inst = 32'hc20ee55;
      10948: inst = 32'h10408000;
      10949: inst = 32'hc4042ed;
      10950: inst = 32'h8220000;
      10951: inst = 32'h10408000;
      10952: inst = 32'hc4043b0;
      10953: inst = 32'h8220000;
      10954: inst = 32'hc20e571;
      10955: inst = 32'h10408000;
      10956: inst = 32'hc404349;
      10957: inst = 32'h8220000;
      10958: inst = 32'h10408000;
      10959: inst = 32'hc40434e;
      10960: inst = 32'h8220000;
      10961: inst = 32'h10408000;
      10962: inst = 32'hc404406;
      10963: inst = 32'h8220000;
      10964: inst = 32'h10408000;
      10965: inst = 32'hc404411;
      10966: inst = 32'h8220000;
      10967: inst = 32'hc20cb28;
      10968: inst = 32'h10408000;
      10969: inst = 32'hc40434a;
      10970: inst = 32'h8220000;
      10971: inst = 32'h10408000;
      10972: inst = 32'hc40434d;
      10973: inst = 32'h8220000;
      10974: inst = 32'h10408000;
      10975: inst = 32'hc404407;
      10976: inst = 32'h8220000;
      10977: inst = 32'h10408000;
      10978: inst = 32'hc404410;
      10979: inst = 32'h8220000;
      10980: inst = 32'hc20cac7;
      10981: inst = 32'h10408000;
      10982: inst = 32'hc40434b;
      10983: inst = 32'h8220000;
      10984: inst = 32'h10408000;
      10985: inst = 32'hc40434c;
      10986: inst = 32'h8220000;
      10987: inst = 32'h10408000;
      10988: inst = 32'hc4043a9;
      10989: inst = 32'h8220000;
      10990: inst = 32'h10408000;
      10991: inst = 32'hc4043aa;
      10992: inst = 32'h8220000;
      10993: inst = 32'h10408000;
      10994: inst = 32'hc4043ab;
      10995: inst = 32'h8220000;
      10996: inst = 32'h10408000;
      10997: inst = 32'hc4043ac;
      10998: inst = 32'h8220000;
      10999: inst = 32'h10408000;
      11000: inst = 32'hc4043ad;
      11001: inst = 32'h8220000;
      11002: inst = 32'h10408000;
      11003: inst = 32'hc4043ae;
      11004: inst = 32'h8220000;
      11005: inst = 32'h10408000;
      11006: inst = 32'hc404408;
      11007: inst = 32'h8220000;
      11008: inst = 32'h10408000;
      11009: inst = 32'hc404409;
      11010: inst = 32'h8220000;
      11011: inst = 32'h10408000;
      11012: inst = 32'hc40440a;
      11013: inst = 32'h8220000;
      11014: inst = 32'h10408000;
      11015: inst = 32'hc40440b;
      11016: inst = 32'h8220000;
      11017: inst = 32'h10408000;
      11018: inst = 32'hc40440c;
      11019: inst = 32'h8220000;
      11020: inst = 32'h10408000;
      11021: inst = 32'hc40440d;
      11022: inst = 32'h8220000;
      11023: inst = 32'h10408000;
      11024: inst = 32'hc40440e;
      11025: inst = 32'h8220000;
      11026: inst = 32'h10408000;
      11027: inst = 32'hc40440f;
      11028: inst = 32'h8220000;
      11029: inst = 32'hc20d40c;
      11030: inst = 32'h10408000;
      11031: inst = 32'hc4043af;
      11032: inst = 32'h8220000;
      11033: inst = 32'hc20ee8e;
      11034: inst = 32'h10408000;
      11035: inst = 32'hc40446a;
      11036: inst = 32'h8220000;
      11037: inst = 32'h10408000;
      11038: inst = 32'hc4044b5;
      11039: inst = 32'h8220000;
      11040: inst = 32'hc20ee48;
      11041: inst = 32'h10408000;
      11042: inst = 32'hc40446b;
      11043: inst = 32'h8220000;
      11044: inst = 32'h10408000;
      11045: inst = 32'hc40446c;
      11046: inst = 32'h8220000;
      11047: inst = 32'h10408000;
      11048: inst = 32'hc4044b3;
      11049: inst = 32'h8220000;
      11050: inst = 32'h10408000;
      11051: inst = 32'hc4044b4;
      11052: inst = 32'h8220000;
      11053: inst = 32'hc20ee90;
      11054: inst = 32'h10408000;
      11055: inst = 32'hc40446d;
      11056: inst = 32'h8220000;
      11057: inst = 32'h10408000;
      11058: inst = 32'hc4044b2;
      11059: inst = 32'h8220000;
      11060: inst = 32'hc20eeb5;
      11061: inst = 32'h10408000;
      11062: inst = 32'hc4044cb;
      11063: inst = 32'h8220000;
      11064: inst = 32'h10408000;
      11065: inst = 32'hc4044cc;
      11066: inst = 32'h8220000;
      11067: inst = 32'h10408000;
      11068: inst = 32'hc404513;
      11069: inst = 32'h8220000;
      11070: inst = 32'h10408000;
      11071: inst = 32'hc404514;
      11072: inst = 32'h8220000;
      11073: inst = 32'hc20c2e2;
      11074: inst = 32'h10408000;
      11075: inst = 32'hc4046ef;
      11076: inst = 32'h8220000;
      11077: inst = 32'h10408000;
      11078: inst = 32'hc4046f0;
      11079: inst = 32'h8220000;
      11080: inst = 32'h10408000;
      11081: inst = 32'hc4046f1;
      11082: inst = 32'h8220000;
      11083: inst = 32'h10408000;
      11084: inst = 32'hc4046f2;
      11085: inst = 32'h8220000;
      11086: inst = 32'h10408000;
      11087: inst = 32'hc4046f3;
      11088: inst = 32'h8220000;
      11089: inst = 32'h10408000;
      11090: inst = 32'hc4046f4;
      11091: inst = 32'h8220000;
      11092: inst = 32'h10408000;
      11093: inst = 32'hc4046f5;
      11094: inst = 32'h8220000;
      11095: inst = 32'h10408000;
      11096: inst = 32'hc4046f6;
      11097: inst = 32'h8220000;
      11098: inst = 32'h10408000;
      11099: inst = 32'hc4046f7;
      11100: inst = 32'h8220000;
      11101: inst = 32'h10408000;
      11102: inst = 32'hc4046f8;
      11103: inst = 32'h8220000;
      11104: inst = 32'h10408000;
      11105: inst = 32'hc4046f9;
      11106: inst = 32'h8220000;
      11107: inst = 32'h10408000;
      11108: inst = 32'hc4046fa;
      11109: inst = 32'h8220000;
      11110: inst = 32'h10408000;
      11111: inst = 32'hc4046fb;
      11112: inst = 32'h8220000;
      11113: inst = 32'h10408000;
      11114: inst = 32'hc4046fc;
      11115: inst = 32'h8220000;
      11116: inst = 32'h10408000;
      11117: inst = 32'hc4046fd;
      11118: inst = 32'h8220000;
      11119: inst = 32'h10408000;
      11120: inst = 32'hc4046fe;
      11121: inst = 32'h8220000;
      11122: inst = 32'h10408000;
      11123: inst = 32'hc4046ff;
      11124: inst = 32'h8220000;
      11125: inst = 32'h10408000;
      11126: inst = 32'hc40474f;
      11127: inst = 32'h8220000;
      11128: inst = 32'h10408000;
      11129: inst = 32'hc40475f;
      11130: inst = 32'h8220000;
      11131: inst = 32'h10408000;
      11132: inst = 32'hc4047af;
      11133: inst = 32'h8220000;
      11134: inst = 32'h10408000;
      11135: inst = 32'hc4047bf;
      11136: inst = 32'h8220000;
      11137: inst = 32'h10408000;
      11138: inst = 32'hc40480f;
      11139: inst = 32'h8220000;
      11140: inst = 32'h10408000;
      11141: inst = 32'hc40481f;
      11142: inst = 32'h8220000;
      11143: inst = 32'h10408000;
      11144: inst = 32'hc40486f;
      11145: inst = 32'h8220000;
      11146: inst = 32'h10408000;
      11147: inst = 32'hc40487f;
      11148: inst = 32'h8220000;
      11149: inst = 32'h10408000;
      11150: inst = 32'hc4048cf;
      11151: inst = 32'h8220000;
      11152: inst = 32'h10408000;
      11153: inst = 32'hc4048df;
      11154: inst = 32'h8220000;
      11155: inst = 32'h10408000;
      11156: inst = 32'hc40492f;
      11157: inst = 32'h8220000;
      11158: inst = 32'h10408000;
      11159: inst = 32'hc40493f;
      11160: inst = 32'h8220000;
      11161: inst = 32'h10408000;
      11162: inst = 32'hc40498f;
      11163: inst = 32'h8220000;
      11164: inst = 32'h10408000;
      11165: inst = 32'hc40499f;
      11166: inst = 32'h8220000;
      11167: inst = 32'h10408000;
      11168: inst = 32'hc4049ef;
      11169: inst = 32'h8220000;
      11170: inst = 32'h10408000;
      11171: inst = 32'hc4049ff;
      11172: inst = 32'h8220000;
      11173: inst = 32'h10408000;
      11174: inst = 32'hc404a4f;
      11175: inst = 32'h8220000;
      11176: inst = 32'h10408000;
      11177: inst = 32'hc404a5f;
      11178: inst = 32'h8220000;
      11179: inst = 32'h10408000;
      11180: inst = 32'hc404aaf;
      11181: inst = 32'h8220000;
      11182: inst = 32'h10408000;
      11183: inst = 32'hc404abf;
      11184: inst = 32'h8220000;
      11185: inst = 32'h10408000;
      11186: inst = 32'hc404b0f;
      11187: inst = 32'h8220000;
      11188: inst = 32'h10408000;
      11189: inst = 32'hc404b1f;
      11190: inst = 32'h8220000;
      11191: inst = 32'h10408000;
      11192: inst = 32'hc404b6f;
      11193: inst = 32'h8220000;
      11194: inst = 32'h10408000;
      11195: inst = 32'hc404b7f;
      11196: inst = 32'h8220000;
      11197: inst = 32'h10408000;
      11198: inst = 32'hc404bcf;
      11199: inst = 32'h8220000;
      11200: inst = 32'h10408000;
      11201: inst = 32'hc404bdf;
      11202: inst = 32'h8220000;
      11203: inst = 32'h10408000;
      11204: inst = 32'hc404c2f;
      11205: inst = 32'h8220000;
      11206: inst = 32'h10408000;
      11207: inst = 32'hc404c3f;
      11208: inst = 32'h8220000;
      11209: inst = 32'h10408000;
      11210: inst = 32'hc404c8f;
      11211: inst = 32'h8220000;
      11212: inst = 32'h10408000;
      11213: inst = 32'hc404c9f;
      11214: inst = 32'h8220000;
      11215: inst = 32'h10408000;
      11216: inst = 32'hc404cef;
      11217: inst = 32'h8220000;
      11218: inst = 32'h10408000;
      11219: inst = 32'hc404cff;
      11220: inst = 32'h8220000;
      11221: inst = 32'h10408000;
      11222: inst = 32'hc404d4f;
      11223: inst = 32'h8220000;
      11224: inst = 32'h10408000;
      11225: inst = 32'hc404d5f;
      11226: inst = 32'h8220000;
      11227: inst = 32'h10408000;
      11228: inst = 32'hc404daf;
      11229: inst = 32'h8220000;
      11230: inst = 32'h10408000;
      11231: inst = 32'hc404dbf;
      11232: inst = 32'h8220000;
      11233: inst = 32'h10408000;
      11234: inst = 32'hc404e0f;
      11235: inst = 32'h8220000;
      11236: inst = 32'h10408000;
      11237: inst = 32'hc404e1f;
      11238: inst = 32'h8220000;
      11239: inst = 32'h10408000;
      11240: inst = 32'hc404e6f;
      11241: inst = 32'h8220000;
      11242: inst = 32'h10408000;
      11243: inst = 32'hc404e7f;
      11244: inst = 32'h8220000;
      11245: inst = 32'h10408000;
      11246: inst = 32'hc404ecf;
      11247: inst = 32'h8220000;
      11248: inst = 32'h10408000;
      11249: inst = 32'hc404edf;
      11250: inst = 32'h8220000;
      11251: inst = 32'h10408000;
      11252: inst = 32'hc404f2f;
      11253: inst = 32'h8220000;
      11254: inst = 32'h10408000;
      11255: inst = 32'hc404f3f;
      11256: inst = 32'h8220000;
      11257: inst = 32'h10408000;
      11258: inst = 32'hc404f8f;
      11259: inst = 32'h8220000;
      11260: inst = 32'h10408000;
      11261: inst = 32'hc404f9f;
      11262: inst = 32'h8220000;
      11263: inst = 32'h10408000;
      11264: inst = 32'hc404fef;
      11265: inst = 32'h8220000;
      11266: inst = 32'h10408000;
      11267: inst = 32'hc404fff;
      11268: inst = 32'h8220000;
      11269: inst = 32'h10408000;
      11270: inst = 32'hc40504f;
      11271: inst = 32'h8220000;
      11272: inst = 32'h10408000;
      11273: inst = 32'hc40505f;
      11274: inst = 32'h8220000;
      11275: inst = 32'h10408000;
      11276: inst = 32'hc4050af;
      11277: inst = 32'h8220000;
      11278: inst = 32'h10408000;
      11279: inst = 32'hc4050bf;
      11280: inst = 32'h8220000;
      11281: inst = 32'h10408000;
      11282: inst = 32'hc40510f;
      11283: inst = 32'h8220000;
      11284: inst = 32'h10408000;
      11285: inst = 32'hc40511f;
      11286: inst = 32'h8220000;
      11287: inst = 32'h10408000;
      11288: inst = 32'hc40516f;
      11289: inst = 32'h8220000;
      11290: inst = 32'h10408000;
      11291: inst = 32'hc40517f;
      11292: inst = 32'h8220000;
      11293: inst = 32'h10408000;
      11294: inst = 32'hc4051cf;
      11295: inst = 32'h8220000;
      11296: inst = 32'h10408000;
      11297: inst = 32'hc4051df;
      11298: inst = 32'h8220000;
      11299: inst = 32'h10408000;
      11300: inst = 32'hc40522f;
      11301: inst = 32'h8220000;
      11302: inst = 32'h10408000;
      11303: inst = 32'hc40523f;
      11304: inst = 32'h8220000;
      11305: inst = 32'h10408000;
      11306: inst = 32'hc40528f;
      11307: inst = 32'h8220000;
      11308: inst = 32'h10408000;
      11309: inst = 32'hc40529f;
      11310: inst = 32'h8220000;
      11311: inst = 32'h10408000;
      11312: inst = 32'hc4052ef;
      11313: inst = 32'h8220000;
      11314: inst = 32'h10408000;
      11315: inst = 32'hc4052f0;
      11316: inst = 32'h8220000;
      11317: inst = 32'h10408000;
      11318: inst = 32'hc4052f1;
      11319: inst = 32'h8220000;
      11320: inst = 32'h10408000;
      11321: inst = 32'hc4052f2;
      11322: inst = 32'h8220000;
      11323: inst = 32'h10408000;
      11324: inst = 32'hc4052f3;
      11325: inst = 32'h8220000;
      11326: inst = 32'h10408000;
      11327: inst = 32'hc4052f4;
      11328: inst = 32'h8220000;
      11329: inst = 32'h10408000;
      11330: inst = 32'hc4052f5;
      11331: inst = 32'h8220000;
      11332: inst = 32'h10408000;
      11333: inst = 32'hc4052f6;
      11334: inst = 32'h8220000;
      11335: inst = 32'h10408000;
      11336: inst = 32'hc4052f7;
      11337: inst = 32'h8220000;
      11338: inst = 32'h10408000;
      11339: inst = 32'hc4052f8;
      11340: inst = 32'h8220000;
      11341: inst = 32'h10408000;
      11342: inst = 32'hc4052f9;
      11343: inst = 32'h8220000;
      11344: inst = 32'h10408000;
      11345: inst = 32'hc4052fa;
      11346: inst = 32'h8220000;
      11347: inst = 32'h10408000;
      11348: inst = 32'hc4052fb;
      11349: inst = 32'h8220000;
      11350: inst = 32'h10408000;
      11351: inst = 32'hc4052fc;
      11352: inst = 32'h8220000;
      11353: inst = 32'h10408000;
      11354: inst = 32'hc4052fd;
      11355: inst = 32'h8220000;
      11356: inst = 32'h10408000;
      11357: inst = 32'hc4052fe;
      11358: inst = 32'h8220000;
      11359: inst = 32'h10408000;
      11360: inst = 32'hc4052ff;
      11361: inst = 32'h8220000;
      11362: inst = 32'hc20dbc5;
      11363: inst = 32'h10408000;
      11364: inst = 32'hc404750;
      11365: inst = 32'h8220000;
      11366: inst = 32'h10408000;
      11367: inst = 32'hc404751;
      11368: inst = 32'h8220000;
      11369: inst = 32'h10408000;
      11370: inst = 32'hc404752;
      11371: inst = 32'h8220000;
      11372: inst = 32'h10408000;
      11373: inst = 32'hc404753;
      11374: inst = 32'h8220000;
      11375: inst = 32'h10408000;
      11376: inst = 32'hc404754;
      11377: inst = 32'h8220000;
      11378: inst = 32'h10408000;
      11379: inst = 32'hc404755;
      11380: inst = 32'h8220000;
      11381: inst = 32'h10408000;
      11382: inst = 32'hc404756;
      11383: inst = 32'h8220000;
      11384: inst = 32'h10408000;
      11385: inst = 32'hc404757;
      11386: inst = 32'h8220000;
      11387: inst = 32'h10408000;
      11388: inst = 32'hc404758;
      11389: inst = 32'h8220000;
      11390: inst = 32'h10408000;
      11391: inst = 32'hc404759;
      11392: inst = 32'h8220000;
      11393: inst = 32'h10408000;
      11394: inst = 32'hc40475a;
      11395: inst = 32'h8220000;
      11396: inst = 32'h10408000;
      11397: inst = 32'hc40475b;
      11398: inst = 32'h8220000;
      11399: inst = 32'h10408000;
      11400: inst = 32'hc40475c;
      11401: inst = 32'h8220000;
      11402: inst = 32'h10408000;
      11403: inst = 32'hc40475d;
      11404: inst = 32'h8220000;
      11405: inst = 32'h10408000;
      11406: inst = 32'hc40475e;
      11407: inst = 32'h8220000;
      11408: inst = 32'h10408000;
      11409: inst = 32'hc4047b0;
      11410: inst = 32'h8220000;
      11411: inst = 32'h10408000;
      11412: inst = 32'hc4047b1;
      11413: inst = 32'h8220000;
      11414: inst = 32'h10408000;
      11415: inst = 32'hc4047b2;
      11416: inst = 32'h8220000;
      11417: inst = 32'h10408000;
      11418: inst = 32'hc4047b3;
      11419: inst = 32'h8220000;
      11420: inst = 32'h10408000;
      11421: inst = 32'hc4047b4;
      11422: inst = 32'h8220000;
      11423: inst = 32'h10408000;
      11424: inst = 32'hc4047b5;
      11425: inst = 32'h8220000;
      11426: inst = 32'h10408000;
      11427: inst = 32'hc4047b6;
      11428: inst = 32'h8220000;
      11429: inst = 32'h10408000;
      11430: inst = 32'hc4047b7;
      11431: inst = 32'h8220000;
      11432: inst = 32'h10408000;
      11433: inst = 32'hc4047b8;
      11434: inst = 32'h8220000;
      11435: inst = 32'h10408000;
      11436: inst = 32'hc4047b9;
      11437: inst = 32'h8220000;
      11438: inst = 32'h10408000;
      11439: inst = 32'hc4047ba;
      11440: inst = 32'h8220000;
      11441: inst = 32'h10408000;
      11442: inst = 32'hc4047bb;
      11443: inst = 32'h8220000;
      11444: inst = 32'h10408000;
      11445: inst = 32'hc4047bc;
      11446: inst = 32'h8220000;
      11447: inst = 32'h10408000;
      11448: inst = 32'hc4047bd;
      11449: inst = 32'h8220000;
      11450: inst = 32'h10408000;
      11451: inst = 32'hc4047be;
      11452: inst = 32'h8220000;
      11453: inst = 32'h10408000;
      11454: inst = 32'hc404810;
      11455: inst = 32'h8220000;
      11456: inst = 32'h10408000;
      11457: inst = 32'hc404811;
      11458: inst = 32'h8220000;
      11459: inst = 32'h10408000;
      11460: inst = 32'hc404812;
      11461: inst = 32'h8220000;
      11462: inst = 32'h10408000;
      11463: inst = 32'hc404813;
      11464: inst = 32'h8220000;
      11465: inst = 32'h10408000;
      11466: inst = 32'hc404814;
      11467: inst = 32'h8220000;
      11468: inst = 32'h10408000;
      11469: inst = 32'hc404815;
      11470: inst = 32'h8220000;
      11471: inst = 32'h10408000;
      11472: inst = 32'hc404816;
      11473: inst = 32'h8220000;
      11474: inst = 32'h10408000;
      11475: inst = 32'hc404817;
      11476: inst = 32'h8220000;
      11477: inst = 32'h10408000;
      11478: inst = 32'hc404818;
      11479: inst = 32'h8220000;
      11480: inst = 32'h10408000;
      11481: inst = 32'hc404819;
      11482: inst = 32'h8220000;
      11483: inst = 32'h10408000;
      11484: inst = 32'hc40481a;
      11485: inst = 32'h8220000;
      11486: inst = 32'h10408000;
      11487: inst = 32'hc40481b;
      11488: inst = 32'h8220000;
      11489: inst = 32'h10408000;
      11490: inst = 32'hc40481c;
      11491: inst = 32'h8220000;
      11492: inst = 32'h10408000;
      11493: inst = 32'hc40481d;
      11494: inst = 32'h8220000;
      11495: inst = 32'h10408000;
      11496: inst = 32'hc40481e;
      11497: inst = 32'h8220000;
      11498: inst = 32'h10408000;
      11499: inst = 32'hc404870;
      11500: inst = 32'h8220000;
      11501: inst = 32'h10408000;
      11502: inst = 32'hc404871;
      11503: inst = 32'h8220000;
      11504: inst = 32'h10408000;
      11505: inst = 32'hc404872;
      11506: inst = 32'h8220000;
      11507: inst = 32'h10408000;
      11508: inst = 32'hc404873;
      11509: inst = 32'h8220000;
      11510: inst = 32'h10408000;
      11511: inst = 32'hc404874;
      11512: inst = 32'h8220000;
      11513: inst = 32'h10408000;
      11514: inst = 32'hc404875;
      11515: inst = 32'h8220000;
      11516: inst = 32'h10408000;
      11517: inst = 32'hc404876;
      11518: inst = 32'h8220000;
      11519: inst = 32'h10408000;
      11520: inst = 32'hc404877;
      11521: inst = 32'h8220000;
      11522: inst = 32'h10408000;
      11523: inst = 32'hc404878;
      11524: inst = 32'h8220000;
      11525: inst = 32'h10408000;
      11526: inst = 32'hc404879;
      11527: inst = 32'h8220000;
      11528: inst = 32'h10408000;
      11529: inst = 32'hc40487a;
      11530: inst = 32'h8220000;
      11531: inst = 32'h10408000;
      11532: inst = 32'hc40487b;
      11533: inst = 32'h8220000;
      11534: inst = 32'h10408000;
      11535: inst = 32'hc40487c;
      11536: inst = 32'h8220000;
      11537: inst = 32'h10408000;
      11538: inst = 32'hc40487d;
      11539: inst = 32'h8220000;
      11540: inst = 32'h10408000;
      11541: inst = 32'hc40487e;
      11542: inst = 32'h8220000;
      11543: inst = 32'h10408000;
      11544: inst = 32'hc4048d0;
      11545: inst = 32'h8220000;
      11546: inst = 32'h10408000;
      11547: inst = 32'hc4048d1;
      11548: inst = 32'h8220000;
      11549: inst = 32'h10408000;
      11550: inst = 32'hc4048d2;
      11551: inst = 32'h8220000;
      11552: inst = 32'h10408000;
      11553: inst = 32'hc4048d3;
      11554: inst = 32'h8220000;
      11555: inst = 32'h10408000;
      11556: inst = 32'hc4048d4;
      11557: inst = 32'h8220000;
      11558: inst = 32'h10408000;
      11559: inst = 32'hc4048d5;
      11560: inst = 32'h8220000;
      11561: inst = 32'h10408000;
      11562: inst = 32'hc4048d6;
      11563: inst = 32'h8220000;
      11564: inst = 32'h10408000;
      11565: inst = 32'hc4048d7;
      11566: inst = 32'h8220000;
      11567: inst = 32'h10408000;
      11568: inst = 32'hc4048d8;
      11569: inst = 32'h8220000;
      11570: inst = 32'h10408000;
      11571: inst = 32'hc4048d9;
      11572: inst = 32'h8220000;
      11573: inst = 32'h10408000;
      11574: inst = 32'hc4048da;
      11575: inst = 32'h8220000;
      11576: inst = 32'h10408000;
      11577: inst = 32'hc4048db;
      11578: inst = 32'h8220000;
      11579: inst = 32'h10408000;
      11580: inst = 32'hc4048dc;
      11581: inst = 32'h8220000;
      11582: inst = 32'h10408000;
      11583: inst = 32'hc4048dd;
      11584: inst = 32'h8220000;
      11585: inst = 32'h10408000;
      11586: inst = 32'hc4048de;
      11587: inst = 32'h8220000;
      11588: inst = 32'h10408000;
      11589: inst = 32'hc404930;
      11590: inst = 32'h8220000;
      11591: inst = 32'h10408000;
      11592: inst = 32'hc404931;
      11593: inst = 32'h8220000;
      11594: inst = 32'h10408000;
      11595: inst = 32'hc404936;
      11596: inst = 32'h8220000;
      11597: inst = 32'h10408000;
      11598: inst = 32'hc404937;
      11599: inst = 32'h8220000;
      11600: inst = 32'h10408000;
      11601: inst = 32'hc404938;
      11602: inst = 32'h8220000;
      11603: inst = 32'h10408000;
      11604: inst = 32'hc404939;
      11605: inst = 32'h8220000;
      11606: inst = 32'h10408000;
      11607: inst = 32'hc40493a;
      11608: inst = 32'h8220000;
      11609: inst = 32'h10408000;
      11610: inst = 32'hc40493b;
      11611: inst = 32'h8220000;
      11612: inst = 32'h10408000;
      11613: inst = 32'hc40493c;
      11614: inst = 32'h8220000;
      11615: inst = 32'h10408000;
      11616: inst = 32'hc40493d;
      11617: inst = 32'h8220000;
      11618: inst = 32'h10408000;
      11619: inst = 32'hc40493e;
      11620: inst = 32'h8220000;
      11621: inst = 32'h10408000;
      11622: inst = 32'hc404990;
      11623: inst = 32'h8220000;
      11624: inst = 32'h10408000;
      11625: inst = 32'hc404991;
      11626: inst = 32'h8220000;
      11627: inst = 32'h10408000;
      11628: inst = 32'hc404996;
      11629: inst = 32'h8220000;
      11630: inst = 32'h10408000;
      11631: inst = 32'hc404997;
      11632: inst = 32'h8220000;
      11633: inst = 32'h10408000;
      11634: inst = 32'hc404998;
      11635: inst = 32'h8220000;
      11636: inst = 32'h10408000;
      11637: inst = 32'hc404999;
      11638: inst = 32'h8220000;
      11639: inst = 32'h10408000;
      11640: inst = 32'hc40499a;
      11641: inst = 32'h8220000;
      11642: inst = 32'h10408000;
      11643: inst = 32'hc40499b;
      11644: inst = 32'h8220000;
      11645: inst = 32'h10408000;
      11646: inst = 32'hc40499c;
      11647: inst = 32'h8220000;
      11648: inst = 32'h10408000;
      11649: inst = 32'hc40499d;
      11650: inst = 32'h8220000;
      11651: inst = 32'h10408000;
      11652: inst = 32'hc40499e;
      11653: inst = 32'h8220000;
      11654: inst = 32'h10408000;
      11655: inst = 32'hc4049f0;
      11656: inst = 32'h8220000;
      11657: inst = 32'h10408000;
      11658: inst = 32'hc4049f1;
      11659: inst = 32'h8220000;
      11660: inst = 32'h10408000;
      11661: inst = 32'hc4049f6;
      11662: inst = 32'h8220000;
      11663: inst = 32'h10408000;
      11664: inst = 32'hc4049f7;
      11665: inst = 32'h8220000;
      11666: inst = 32'h10408000;
      11667: inst = 32'hc4049f8;
      11668: inst = 32'h8220000;
      11669: inst = 32'h10408000;
      11670: inst = 32'hc4049f9;
      11671: inst = 32'h8220000;
      11672: inst = 32'h10408000;
      11673: inst = 32'hc4049fa;
      11674: inst = 32'h8220000;
      11675: inst = 32'h10408000;
      11676: inst = 32'hc4049fb;
      11677: inst = 32'h8220000;
      11678: inst = 32'h10408000;
      11679: inst = 32'hc4049fc;
      11680: inst = 32'h8220000;
      11681: inst = 32'h10408000;
      11682: inst = 32'hc4049fd;
      11683: inst = 32'h8220000;
      11684: inst = 32'h10408000;
      11685: inst = 32'hc4049fe;
      11686: inst = 32'h8220000;
      11687: inst = 32'h10408000;
      11688: inst = 32'hc404a50;
      11689: inst = 32'h8220000;
      11690: inst = 32'h10408000;
      11691: inst = 32'hc404a51;
      11692: inst = 32'h8220000;
      11693: inst = 32'h10408000;
      11694: inst = 32'hc404a56;
      11695: inst = 32'h8220000;
      11696: inst = 32'h10408000;
      11697: inst = 32'hc404a57;
      11698: inst = 32'h8220000;
      11699: inst = 32'h10408000;
      11700: inst = 32'hc404a58;
      11701: inst = 32'h8220000;
      11702: inst = 32'h10408000;
      11703: inst = 32'hc404a59;
      11704: inst = 32'h8220000;
      11705: inst = 32'h10408000;
      11706: inst = 32'hc404a5a;
      11707: inst = 32'h8220000;
      11708: inst = 32'h10408000;
      11709: inst = 32'hc404a5b;
      11710: inst = 32'h8220000;
      11711: inst = 32'h10408000;
      11712: inst = 32'hc404a5c;
      11713: inst = 32'h8220000;
      11714: inst = 32'h10408000;
      11715: inst = 32'hc404a5d;
      11716: inst = 32'h8220000;
      11717: inst = 32'h10408000;
      11718: inst = 32'hc404a5e;
      11719: inst = 32'h8220000;
      11720: inst = 32'h10408000;
      11721: inst = 32'hc404ab0;
      11722: inst = 32'h8220000;
      11723: inst = 32'h10408000;
      11724: inst = 32'hc404ab1;
      11725: inst = 32'h8220000;
      11726: inst = 32'h10408000;
      11727: inst = 32'hc404ab6;
      11728: inst = 32'h8220000;
      11729: inst = 32'h10408000;
      11730: inst = 32'hc404ab7;
      11731: inst = 32'h8220000;
      11732: inst = 32'h10408000;
      11733: inst = 32'hc404ab8;
      11734: inst = 32'h8220000;
      11735: inst = 32'h10408000;
      11736: inst = 32'hc404ab9;
      11737: inst = 32'h8220000;
      11738: inst = 32'h10408000;
      11739: inst = 32'hc404aba;
      11740: inst = 32'h8220000;
      11741: inst = 32'h10408000;
      11742: inst = 32'hc404abb;
      11743: inst = 32'h8220000;
      11744: inst = 32'h10408000;
      11745: inst = 32'hc404abc;
      11746: inst = 32'h8220000;
      11747: inst = 32'h10408000;
      11748: inst = 32'hc404abd;
      11749: inst = 32'h8220000;
      11750: inst = 32'h10408000;
      11751: inst = 32'hc404abe;
      11752: inst = 32'h8220000;
      11753: inst = 32'h10408000;
      11754: inst = 32'hc404b10;
      11755: inst = 32'h8220000;
      11756: inst = 32'h10408000;
      11757: inst = 32'hc404b11;
      11758: inst = 32'h8220000;
      11759: inst = 32'h10408000;
      11760: inst = 32'hc404b16;
      11761: inst = 32'h8220000;
      11762: inst = 32'h10408000;
      11763: inst = 32'hc404b17;
      11764: inst = 32'h8220000;
      11765: inst = 32'h10408000;
      11766: inst = 32'hc404b18;
      11767: inst = 32'h8220000;
      11768: inst = 32'h10408000;
      11769: inst = 32'hc404b19;
      11770: inst = 32'h8220000;
      11771: inst = 32'h10408000;
      11772: inst = 32'hc404b1a;
      11773: inst = 32'h8220000;
      11774: inst = 32'h10408000;
      11775: inst = 32'hc404b1b;
      11776: inst = 32'h8220000;
      11777: inst = 32'h10408000;
      11778: inst = 32'hc404b1c;
      11779: inst = 32'h8220000;
      11780: inst = 32'h10408000;
      11781: inst = 32'hc404b1d;
      11782: inst = 32'h8220000;
      11783: inst = 32'h10408000;
      11784: inst = 32'hc404b1e;
      11785: inst = 32'h8220000;
      11786: inst = 32'h10408000;
      11787: inst = 32'hc404b70;
      11788: inst = 32'h8220000;
      11789: inst = 32'h10408000;
      11790: inst = 32'hc404b71;
      11791: inst = 32'h8220000;
      11792: inst = 32'h10408000;
      11793: inst = 32'hc404b76;
      11794: inst = 32'h8220000;
      11795: inst = 32'h10408000;
      11796: inst = 32'hc404b77;
      11797: inst = 32'h8220000;
      11798: inst = 32'h10408000;
      11799: inst = 32'hc404b78;
      11800: inst = 32'h8220000;
      11801: inst = 32'h10408000;
      11802: inst = 32'hc404b79;
      11803: inst = 32'h8220000;
      11804: inst = 32'h10408000;
      11805: inst = 32'hc404b7a;
      11806: inst = 32'h8220000;
      11807: inst = 32'h10408000;
      11808: inst = 32'hc404b7b;
      11809: inst = 32'h8220000;
      11810: inst = 32'h10408000;
      11811: inst = 32'hc404b7c;
      11812: inst = 32'h8220000;
      11813: inst = 32'h10408000;
      11814: inst = 32'hc404b7d;
      11815: inst = 32'h8220000;
      11816: inst = 32'h10408000;
      11817: inst = 32'hc404b7e;
      11818: inst = 32'h8220000;
      11819: inst = 32'h10408000;
      11820: inst = 32'hc404bd0;
      11821: inst = 32'h8220000;
      11822: inst = 32'h10408000;
      11823: inst = 32'hc404bd1;
      11824: inst = 32'h8220000;
      11825: inst = 32'h10408000;
      11826: inst = 32'hc404bd2;
      11827: inst = 32'h8220000;
      11828: inst = 32'h10408000;
      11829: inst = 32'hc404bd3;
      11830: inst = 32'h8220000;
      11831: inst = 32'h10408000;
      11832: inst = 32'hc404bd4;
      11833: inst = 32'h8220000;
      11834: inst = 32'h10408000;
      11835: inst = 32'hc404bd5;
      11836: inst = 32'h8220000;
      11837: inst = 32'h10408000;
      11838: inst = 32'hc404bd6;
      11839: inst = 32'h8220000;
      11840: inst = 32'h10408000;
      11841: inst = 32'hc404bd7;
      11842: inst = 32'h8220000;
      11843: inst = 32'h10408000;
      11844: inst = 32'hc404bd8;
      11845: inst = 32'h8220000;
      11846: inst = 32'h10408000;
      11847: inst = 32'hc404bd9;
      11848: inst = 32'h8220000;
      11849: inst = 32'h10408000;
      11850: inst = 32'hc404bda;
      11851: inst = 32'h8220000;
      11852: inst = 32'h10408000;
      11853: inst = 32'hc404bdb;
      11854: inst = 32'h8220000;
      11855: inst = 32'h10408000;
      11856: inst = 32'hc404bdc;
      11857: inst = 32'h8220000;
      11858: inst = 32'h10408000;
      11859: inst = 32'hc404bdd;
      11860: inst = 32'h8220000;
      11861: inst = 32'h10408000;
      11862: inst = 32'hc404bde;
      11863: inst = 32'h8220000;
      11864: inst = 32'h10408000;
      11865: inst = 32'hc404c30;
      11866: inst = 32'h8220000;
      11867: inst = 32'h10408000;
      11868: inst = 32'hc404c31;
      11869: inst = 32'h8220000;
      11870: inst = 32'h10408000;
      11871: inst = 32'hc404c32;
      11872: inst = 32'h8220000;
      11873: inst = 32'h10408000;
      11874: inst = 32'hc404c33;
      11875: inst = 32'h8220000;
      11876: inst = 32'h10408000;
      11877: inst = 32'hc404c34;
      11878: inst = 32'h8220000;
      11879: inst = 32'h10408000;
      11880: inst = 32'hc404c35;
      11881: inst = 32'h8220000;
      11882: inst = 32'h10408000;
      11883: inst = 32'hc404c36;
      11884: inst = 32'h8220000;
      11885: inst = 32'h10408000;
      11886: inst = 32'hc404c37;
      11887: inst = 32'h8220000;
      11888: inst = 32'h10408000;
      11889: inst = 32'hc404c38;
      11890: inst = 32'h8220000;
      11891: inst = 32'h10408000;
      11892: inst = 32'hc404c39;
      11893: inst = 32'h8220000;
      11894: inst = 32'h10408000;
      11895: inst = 32'hc404c3a;
      11896: inst = 32'h8220000;
      11897: inst = 32'h10408000;
      11898: inst = 32'hc404c3b;
      11899: inst = 32'h8220000;
      11900: inst = 32'h10408000;
      11901: inst = 32'hc404c3c;
      11902: inst = 32'h8220000;
      11903: inst = 32'h10408000;
      11904: inst = 32'hc404c3d;
      11905: inst = 32'h8220000;
      11906: inst = 32'h10408000;
      11907: inst = 32'hc404c3e;
      11908: inst = 32'h8220000;
      11909: inst = 32'h10408000;
      11910: inst = 32'hc404c90;
      11911: inst = 32'h8220000;
      11912: inst = 32'h10408000;
      11913: inst = 32'hc404c91;
      11914: inst = 32'h8220000;
      11915: inst = 32'h10408000;
      11916: inst = 32'hc404c92;
      11917: inst = 32'h8220000;
      11918: inst = 32'h10408000;
      11919: inst = 32'hc404c93;
      11920: inst = 32'h8220000;
      11921: inst = 32'h10408000;
      11922: inst = 32'hc404c94;
      11923: inst = 32'h8220000;
      11924: inst = 32'h10408000;
      11925: inst = 32'hc404c95;
      11926: inst = 32'h8220000;
      11927: inst = 32'h10408000;
      11928: inst = 32'hc404c96;
      11929: inst = 32'h8220000;
      11930: inst = 32'h10408000;
      11931: inst = 32'hc404c97;
      11932: inst = 32'h8220000;
      11933: inst = 32'h10408000;
      11934: inst = 32'hc404c98;
      11935: inst = 32'h8220000;
      11936: inst = 32'h10408000;
      11937: inst = 32'hc404c99;
      11938: inst = 32'h8220000;
      11939: inst = 32'h10408000;
      11940: inst = 32'hc404c9a;
      11941: inst = 32'h8220000;
      11942: inst = 32'h10408000;
      11943: inst = 32'hc404c9b;
      11944: inst = 32'h8220000;
      11945: inst = 32'h10408000;
      11946: inst = 32'hc404c9c;
      11947: inst = 32'h8220000;
      11948: inst = 32'h10408000;
      11949: inst = 32'hc404c9d;
      11950: inst = 32'h8220000;
      11951: inst = 32'h10408000;
      11952: inst = 32'hc404c9e;
      11953: inst = 32'h8220000;
      11954: inst = 32'h10408000;
      11955: inst = 32'hc404cf0;
      11956: inst = 32'h8220000;
      11957: inst = 32'h10408000;
      11958: inst = 32'hc404cf1;
      11959: inst = 32'h8220000;
      11960: inst = 32'h10408000;
      11961: inst = 32'hc404cf2;
      11962: inst = 32'h8220000;
      11963: inst = 32'h10408000;
      11964: inst = 32'hc404cf3;
      11965: inst = 32'h8220000;
      11966: inst = 32'h10408000;
      11967: inst = 32'hc404cf4;
      11968: inst = 32'h8220000;
      11969: inst = 32'h10408000;
      11970: inst = 32'hc404cf5;
      11971: inst = 32'h8220000;
      11972: inst = 32'h10408000;
      11973: inst = 32'hc404cf6;
      11974: inst = 32'h8220000;
      11975: inst = 32'h10408000;
      11976: inst = 32'hc404cf7;
      11977: inst = 32'h8220000;
      11978: inst = 32'h10408000;
      11979: inst = 32'hc404cf8;
      11980: inst = 32'h8220000;
      11981: inst = 32'h10408000;
      11982: inst = 32'hc404cf9;
      11983: inst = 32'h8220000;
      11984: inst = 32'h10408000;
      11985: inst = 32'hc404cfa;
      11986: inst = 32'h8220000;
      11987: inst = 32'h10408000;
      11988: inst = 32'hc404cfe;
      11989: inst = 32'h8220000;
      11990: inst = 32'h10408000;
      11991: inst = 32'hc404d50;
      11992: inst = 32'h8220000;
      11993: inst = 32'h10408000;
      11994: inst = 32'hc404d51;
      11995: inst = 32'h8220000;
      11996: inst = 32'h10408000;
      11997: inst = 32'hc404d52;
      11998: inst = 32'h8220000;
      11999: inst = 32'h10408000;
      12000: inst = 32'hc404d53;
      12001: inst = 32'h8220000;
      12002: inst = 32'h10408000;
      12003: inst = 32'hc404d54;
      12004: inst = 32'h8220000;
      12005: inst = 32'h10408000;
      12006: inst = 32'hc404d55;
      12007: inst = 32'h8220000;
      12008: inst = 32'h10408000;
      12009: inst = 32'hc404d56;
      12010: inst = 32'h8220000;
      12011: inst = 32'h10408000;
      12012: inst = 32'hc404d57;
      12013: inst = 32'h8220000;
      12014: inst = 32'h10408000;
      12015: inst = 32'hc404d58;
      12016: inst = 32'h8220000;
      12017: inst = 32'h10408000;
      12018: inst = 32'hc404d59;
      12019: inst = 32'h8220000;
      12020: inst = 32'h10408000;
      12021: inst = 32'hc404d5a;
      12022: inst = 32'h8220000;
      12023: inst = 32'h10408000;
      12024: inst = 32'hc404d5c;
      12025: inst = 32'h8220000;
      12026: inst = 32'h10408000;
      12027: inst = 32'hc404d5d;
      12028: inst = 32'h8220000;
      12029: inst = 32'h10408000;
      12030: inst = 32'hc404d5e;
      12031: inst = 32'h8220000;
      12032: inst = 32'h10408000;
      12033: inst = 32'hc404db0;
      12034: inst = 32'h8220000;
      12035: inst = 32'h10408000;
      12036: inst = 32'hc404db1;
      12037: inst = 32'h8220000;
      12038: inst = 32'h10408000;
      12039: inst = 32'hc404db2;
      12040: inst = 32'h8220000;
      12041: inst = 32'h10408000;
      12042: inst = 32'hc404db3;
      12043: inst = 32'h8220000;
      12044: inst = 32'h10408000;
      12045: inst = 32'hc404db4;
      12046: inst = 32'h8220000;
      12047: inst = 32'h10408000;
      12048: inst = 32'hc404db5;
      12049: inst = 32'h8220000;
      12050: inst = 32'h10408000;
      12051: inst = 32'hc404db6;
      12052: inst = 32'h8220000;
      12053: inst = 32'h10408000;
      12054: inst = 32'hc404db7;
      12055: inst = 32'h8220000;
      12056: inst = 32'h10408000;
      12057: inst = 32'hc404db8;
      12058: inst = 32'h8220000;
      12059: inst = 32'h10408000;
      12060: inst = 32'hc404db9;
      12061: inst = 32'h8220000;
      12062: inst = 32'h10408000;
      12063: inst = 32'hc404dba;
      12064: inst = 32'h8220000;
      12065: inst = 32'h10408000;
      12066: inst = 32'hc404dbb;
      12067: inst = 32'h8220000;
      12068: inst = 32'h10408000;
      12069: inst = 32'hc404dbc;
      12070: inst = 32'h8220000;
      12071: inst = 32'h10408000;
      12072: inst = 32'hc404dbd;
      12073: inst = 32'h8220000;
      12074: inst = 32'h10408000;
      12075: inst = 32'hc404dbe;
      12076: inst = 32'h8220000;
      12077: inst = 32'h10408000;
      12078: inst = 32'hc404e10;
      12079: inst = 32'h8220000;
      12080: inst = 32'h10408000;
      12081: inst = 32'hc404e11;
      12082: inst = 32'h8220000;
      12083: inst = 32'h10408000;
      12084: inst = 32'hc404e12;
      12085: inst = 32'h8220000;
      12086: inst = 32'h10408000;
      12087: inst = 32'hc404e13;
      12088: inst = 32'h8220000;
      12089: inst = 32'h10408000;
      12090: inst = 32'hc404e14;
      12091: inst = 32'h8220000;
      12092: inst = 32'h10408000;
      12093: inst = 32'hc404e15;
      12094: inst = 32'h8220000;
      12095: inst = 32'h10408000;
      12096: inst = 32'hc404e16;
      12097: inst = 32'h8220000;
      12098: inst = 32'h10408000;
      12099: inst = 32'hc404e17;
      12100: inst = 32'h8220000;
      12101: inst = 32'h10408000;
      12102: inst = 32'hc404e18;
      12103: inst = 32'h8220000;
      12104: inst = 32'h10408000;
      12105: inst = 32'hc404e19;
      12106: inst = 32'h8220000;
      12107: inst = 32'h10408000;
      12108: inst = 32'hc404e1a;
      12109: inst = 32'h8220000;
      12110: inst = 32'h10408000;
      12111: inst = 32'hc404e1b;
      12112: inst = 32'h8220000;
      12113: inst = 32'h10408000;
      12114: inst = 32'hc404e1c;
      12115: inst = 32'h8220000;
      12116: inst = 32'h10408000;
      12117: inst = 32'hc404e1d;
      12118: inst = 32'h8220000;
      12119: inst = 32'h10408000;
      12120: inst = 32'hc404e1e;
      12121: inst = 32'h8220000;
      12122: inst = 32'h10408000;
      12123: inst = 32'hc404e70;
      12124: inst = 32'h8220000;
      12125: inst = 32'h10408000;
      12126: inst = 32'hc404e71;
      12127: inst = 32'h8220000;
      12128: inst = 32'h10408000;
      12129: inst = 32'hc404e72;
      12130: inst = 32'h8220000;
      12131: inst = 32'h10408000;
      12132: inst = 32'hc404e73;
      12133: inst = 32'h8220000;
      12134: inst = 32'h10408000;
      12135: inst = 32'hc404e74;
      12136: inst = 32'h8220000;
      12137: inst = 32'h10408000;
      12138: inst = 32'hc404e75;
      12139: inst = 32'h8220000;
      12140: inst = 32'h10408000;
      12141: inst = 32'hc404e76;
      12142: inst = 32'h8220000;
      12143: inst = 32'h10408000;
      12144: inst = 32'hc404e77;
      12145: inst = 32'h8220000;
      12146: inst = 32'h10408000;
      12147: inst = 32'hc404e78;
      12148: inst = 32'h8220000;
      12149: inst = 32'h10408000;
      12150: inst = 32'hc404e79;
      12151: inst = 32'h8220000;
      12152: inst = 32'h10408000;
      12153: inst = 32'hc404e7a;
      12154: inst = 32'h8220000;
      12155: inst = 32'h10408000;
      12156: inst = 32'hc404e7b;
      12157: inst = 32'h8220000;
      12158: inst = 32'h10408000;
      12159: inst = 32'hc404e7c;
      12160: inst = 32'h8220000;
      12161: inst = 32'h10408000;
      12162: inst = 32'hc404e7d;
      12163: inst = 32'h8220000;
      12164: inst = 32'h10408000;
      12165: inst = 32'hc404e7e;
      12166: inst = 32'h8220000;
      12167: inst = 32'h10408000;
      12168: inst = 32'hc404ed0;
      12169: inst = 32'h8220000;
      12170: inst = 32'h10408000;
      12171: inst = 32'hc404ed1;
      12172: inst = 32'h8220000;
      12173: inst = 32'h10408000;
      12174: inst = 32'hc404ed2;
      12175: inst = 32'h8220000;
      12176: inst = 32'h10408000;
      12177: inst = 32'hc404ed3;
      12178: inst = 32'h8220000;
      12179: inst = 32'h10408000;
      12180: inst = 32'hc404ed4;
      12181: inst = 32'h8220000;
      12182: inst = 32'h10408000;
      12183: inst = 32'hc404ed5;
      12184: inst = 32'h8220000;
      12185: inst = 32'h10408000;
      12186: inst = 32'hc404ed6;
      12187: inst = 32'h8220000;
      12188: inst = 32'h10408000;
      12189: inst = 32'hc404ed7;
      12190: inst = 32'h8220000;
      12191: inst = 32'h10408000;
      12192: inst = 32'hc404ed8;
      12193: inst = 32'h8220000;
      12194: inst = 32'h10408000;
      12195: inst = 32'hc404ed9;
      12196: inst = 32'h8220000;
      12197: inst = 32'h10408000;
      12198: inst = 32'hc404eda;
      12199: inst = 32'h8220000;
      12200: inst = 32'h10408000;
      12201: inst = 32'hc404edb;
      12202: inst = 32'h8220000;
      12203: inst = 32'h10408000;
      12204: inst = 32'hc404edc;
      12205: inst = 32'h8220000;
      12206: inst = 32'h10408000;
      12207: inst = 32'hc404edd;
      12208: inst = 32'h8220000;
      12209: inst = 32'h10408000;
      12210: inst = 32'hc404ede;
      12211: inst = 32'h8220000;
      12212: inst = 32'h10408000;
      12213: inst = 32'hc404f30;
      12214: inst = 32'h8220000;
      12215: inst = 32'h10408000;
      12216: inst = 32'hc404f31;
      12217: inst = 32'h8220000;
      12218: inst = 32'h10408000;
      12219: inst = 32'hc404f32;
      12220: inst = 32'h8220000;
      12221: inst = 32'h10408000;
      12222: inst = 32'hc404f33;
      12223: inst = 32'h8220000;
      12224: inst = 32'h10408000;
      12225: inst = 32'hc404f34;
      12226: inst = 32'h8220000;
      12227: inst = 32'h10408000;
      12228: inst = 32'hc404f35;
      12229: inst = 32'h8220000;
      12230: inst = 32'h10408000;
      12231: inst = 32'hc404f36;
      12232: inst = 32'h8220000;
      12233: inst = 32'h10408000;
      12234: inst = 32'hc404f37;
      12235: inst = 32'h8220000;
      12236: inst = 32'h10408000;
      12237: inst = 32'hc404f38;
      12238: inst = 32'h8220000;
      12239: inst = 32'h10408000;
      12240: inst = 32'hc404f39;
      12241: inst = 32'h8220000;
      12242: inst = 32'h10408000;
      12243: inst = 32'hc404f3a;
      12244: inst = 32'h8220000;
      12245: inst = 32'h10408000;
      12246: inst = 32'hc404f3b;
      12247: inst = 32'h8220000;
      12248: inst = 32'h10408000;
      12249: inst = 32'hc404f3c;
      12250: inst = 32'h8220000;
      12251: inst = 32'h10408000;
      12252: inst = 32'hc404f3d;
      12253: inst = 32'h8220000;
      12254: inst = 32'h10408000;
      12255: inst = 32'hc404f3e;
      12256: inst = 32'h8220000;
      12257: inst = 32'h10408000;
      12258: inst = 32'hc404f90;
      12259: inst = 32'h8220000;
      12260: inst = 32'h10408000;
      12261: inst = 32'hc404f91;
      12262: inst = 32'h8220000;
      12263: inst = 32'h10408000;
      12264: inst = 32'hc404f92;
      12265: inst = 32'h8220000;
      12266: inst = 32'h10408000;
      12267: inst = 32'hc404f93;
      12268: inst = 32'h8220000;
      12269: inst = 32'h10408000;
      12270: inst = 32'hc404f94;
      12271: inst = 32'h8220000;
      12272: inst = 32'h10408000;
      12273: inst = 32'hc404f95;
      12274: inst = 32'h8220000;
      12275: inst = 32'h10408000;
      12276: inst = 32'hc404f96;
      12277: inst = 32'h8220000;
      12278: inst = 32'h10408000;
      12279: inst = 32'hc404f97;
      12280: inst = 32'h8220000;
      12281: inst = 32'h10408000;
      12282: inst = 32'hc404f98;
      12283: inst = 32'h8220000;
      12284: inst = 32'h10408000;
      12285: inst = 32'hc404f99;
      12286: inst = 32'h8220000;
      12287: inst = 32'h10408000;
      12288: inst = 32'hc404f9a;
      12289: inst = 32'h8220000;
      12290: inst = 32'h10408000;
      12291: inst = 32'hc404f9b;
      12292: inst = 32'h8220000;
      12293: inst = 32'h10408000;
      12294: inst = 32'hc404f9c;
      12295: inst = 32'h8220000;
      12296: inst = 32'h10408000;
      12297: inst = 32'hc404f9d;
      12298: inst = 32'h8220000;
      12299: inst = 32'h10408000;
      12300: inst = 32'hc404f9e;
      12301: inst = 32'h8220000;
      12302: inst = 32'h10408000;
      12303: inst = 32'hc404ff0;
      12304: inst = 32'h8220000;
      12305: inst = 32'h10408000;
      12306: inst = 32'hc404ff1;
      12307: inst = 32'h8220000;
      12308: inst = 32'h10408000;
      12309: inst = 32'hc404ff2;
      12310: inst = 32'h8220000;
      12311: inst = 32'h10408000;
      12312: inst = 32'hc404ff3;
      12313: inst = 32'h8220000;
      12314: inst = 32'h10408000;
      12315: inst = 32'hc404ff4;
      12316: inst = 32'h8220000;
      12317: inst = 32'h10408000;
      12318: inst = 32'hc404ff5;
      12319: inst = 32'h8220000;
      12320: inst = 32'h10408000;
      12321: inst = 32'hc404ff6;
      12322: inst = 32'h8220000;
      12323: inst = 32'h10408000;
      12324: inst = 32'hc404ff7;
      12325: inst = 32'h8220000;
      12326: inst = 32'h10408000;
      12327: inst = 32'hc404ff8;
      12328: inst = 32'h8220000;
      12329: inst = 32'h10408000;
      12330: inst = 32'hc404ff9;
      12331: inst = 32'h8220000;
      12332: inst = 32'h10408000;
      12333: inst = 32'hc404ffa;
      12334: inst = 32'h8220000;
      12335: inst = 32'h10408000;
      12336: inst = 32'hc404ffb;
      12337: inst = 32'h8220000;
      12338: inst = 32'h10408000;
      12339: inst = 32'hc404ffc;
      12340: inst = 32'h8220000;
      12341: inst = 32'h10408000;
      12342: inst = 32'hc404ffd;
      12343: inst = 32'h8220000;
      12344: inst = 32'h10408000;
      12345: inst = 32'hc404ffe;
      12346: inst = 32'h8220000;
      12347: inst = 32'h10408000;
      12348: inst = 32'hc405050;
      12349: inst = 32'h8220000;
      12350: inst = 32'h10408000;
      12351: inst = 32'hc405051;
      12352: inst = 32'h8220000;
      12353: inst = 32'h10408000;
      12354: inst = 32'hc405052;
      12355: inst = 32'h8220000;
      12356: inst = 32'h10408000;
      12357: inst = 32'hc405053;
      12358: inst = 32'h8220000;
      12359: inst = 32'h10408000;
      12360: inst = 32'hc405054;
      12361: inst = 32'h8220000;
      12362: inst = 32'h10408000;
      12363: inst = 32'hc405055;
      12364: inst = 32'h8220000;
      12365: inst = 32'h10408000;
      12366: inst = 32'hc405056;
      12367: inst = 32'h8220000;
      12368: inst = 32'h10408000;
      12369: inst = 32'hc405057;
      12370: inst = 32'h8220000;
      12371: inst = 32'h10408000;
      12372: inst = 32'hc405058;
      12373: inst = 32'h8220000;
      12374: inst = 32'h10408000;
      12375: inst = 32'hc405059;
      12376: inst = 32'h8220000;
      12377: inst = 32'h10408000;
      12378: inst = 32'hc40505a;
      12379: inst = 32'h8220000;
      12380: inst = 32'h10408000;
      12381: inst = 32'hc40505b;
      12382: inst = 32'h8220000;
      12383: inst = 32'h10408000;
      12384: inst = 32'hc40505c;
      12385: inst = 32'h8220000;
      12386: inst = 32'h10408000;
      12387: inst = 32'hc40505d;
      12388: inst = 32'h8220000;
      12389: inst = 32'h10408000;
      12390: inst = 32'hc40505e;
      12391: inst = 32'h8220000;
      12392: inst = 32'h10408000;
      12393: inst = 32'hc4050b0;
      12394: inst = 32'h8220000;
      12395: inst = 32'h10408000;
      12396: inst = 32'hc4050b1;
      12397: inst = 32'h8220000;
      12398: inst = 32'h10408000;
      12399: inst = 32'hc4050b2;
      12400: inst = 32'h8220000;
      12401: inst = 32'h10408000;
      12402: inst = 32'hc4050b3;
      12403: inst = 32'h8220000;
      12404: inst = 32'h10408000;
      12405: inst = 32'hc4050b4;
      12406: inst = 32'h8220000;
      12407: inst = 32'h10408000;
      12408: inst = 32'hc4050b5;
      12409: inst = 32'h8220000;
      12410: inst = 32'h10408000;
      12411: inst = 32'hc4050b6;
      12412: inst = 32'h8220000;
      12413: inst = 32'h10408000;
      12414: inst = 32'hc4050b7;
      12415: inst = 32'h8220000;
      12416: inst = 32'h10408000;
      12417: inst = 32'hc4050b8;
      12418: inst = 32'h8220000;
      12419: inst = 32'h10408000;
      12420: inst = 32'hc4050b9;
      12421: inst = 32'h8220000;
      12422: inst = 32'h10408000;
      12423: inst = 32'hc4050ba;
      12424: inst = 32'h8220000;
      12425: inst = 32'h10408000;
      12426: inst = 32'hc4050bb;
      12427: inst = 32'h8220000;
      12428: inst = 32'h10408000;
      12429: inst = 32'hc4050bc;
      12430: inst = 32'h8220000;
      12431: inst = 32'h10408000;
      12432: inst = 32'hc4050bd;
      12433: inst = 32'h8220000;
      12434: inst = 32'h10408000;
      12435: inst = 32'hc4050be;
      12436: inst = 32'h8220000;
      12437: inst = 32'h10408000;
      12438: inst = 32'hc405110;
      12439: inst = 32'h8220000;
      12440: inst = 32'h10408000;
      12441: inst = 32'hc405111;
      12442: inst = 32'h8220000;
      12443: inst = 32'h10408000;
      12444: inst = 32'hc405112;
      12445: inst = 32'h8220000;
      12446: inst = 32'h10408000;
      12447: inst = 32'hc405113;
      12448: inst = 32'h8220000;
      12449: inst = 32'h10408000;
      12450: inst = 32'hc405114;
      12451: inst = 32'h8220000;
      12452: inst = 32'h10408000;
      12453: inst = 32'hc405115;
      12454: inst = 32'h8220000;
      12455: inst = 32'h10408000;
      12456: inst = 32'hc405116;
      12457: inst = 32'h8220000;
      12458: inst = 32'h10408000;
      12459: inst = 32'hc405117;
      12460: inst = 32'h8220000;
      12461: inst = 32'h10408000;
      12462: inst = 32'hc405118;
      12463: inst = 32'h8220000;
      12464: inst = 32'h10408000;
      12465: inst = 32'hc405119;
      12466: inst = 32'h8220000;
      12467: inst = 32'h10408000;
      12468: inst = 32'hc40511a;
      12469: inst = 32'h8220000;
      12470: inst = 32'h10408000;
      12471: inst = 32'hc40511b;
      12472: inst = 32'h8220000;
      12473: inst = 32'h10408000;
      12474: inst = 32'hc40511c;
      12475: inst = 32'h8220000;
      12476: inst = 32'h10408000;
      12477: inst = 32'hc40511d;
      12478: inst = 32'h8220000;
      12479: inst = 32'h10408000;
      12480: inst = 32'hc40511e;
      12481: inst = 32'h8220000;
      12482: inst = 32'h10408000;
      12483: inst = 32'hc405170;
      12484: inst = 32'h8220000;
      12485: inst = 32'h10408000;
      12486: inst = 32'hc405171;
      12487: inst = 32'h8220000;
      12488: inst = 32'h10408000;
      12489: inst = 32'hc405172;
      12490: inst = 32'h8220000;
      12491: inst = 32'h10408000;
      12492: inst = 32'hc405173;
      12493: inst = 32'h8220000;
      12494: inst = 32'h10408000;
      12495: inst = 32'hc405174;
      12496: inst = 32'h8220000;
      12497: inst = 32'h10408000;
      12498: inst = 32'hc405175;
      12499: inst = 32'h8220000;
      12500: inst = 32'h10408000;
      12501: inst = 32'hc405176;
      12502: inst = 32'h8220000;
      12503: inst = 32'h10408000;
      12504: inst = 32'hc405177;
      12505: inst = 32'h8220000;
      12506: inst = 32'h10408000;
      12507: inst = 32'hc405178;
      12508: inst = 32'h8220000;
      12509: inst = 32'h10408000;
      12510: inst = 32'hc405179;
      12511: inst = 32'h8220000;
      12512: inst = 32'h10408000;
      12513: inst = 32'hc40517a;
      12514: inst = 32'h8220000;
      12515: inst = 32'h10408000;
      12516: inst = 32'hc40517b;
      12517: inst = 32'h8220000;
      12518: inst = 32'h10408000;
      12519: inst = 32'hc40517c;
      12520: inst = 32'h8220000;
      12521: inst = 32'h10408000;
      12522: inst = 32'hc40517d;
      12523: inst = 32'h8220000;
      12524: inst = 32'h10408000;
      12525: inst = 32'hc40517e;
      12526: inst = 32'h8220000;
      12527: inst = 32'h10408000;
      12528: inst = 32'hc4051d0;
      12529: inst = 32'h8220000;
      12530: inst = 32'h10408000;
      12531: inst = 32'hc4051d1;
      12532: inst = 32'h8220000;
      12533: inst = 32'h10408000;
      12534: inst = 32'hc4051d2;
      12535: inst = 32'h8220000;
      12536: inst = 32'h10408000;
      12537: inst = 32'hc4051d3;
      12538: inst = 32'h8220000;
      12539: inst = 32'h10408000;
      12540: inst = 32'hc4051d4;
      12541: inst = 32'h8220000;
      12542: inst = 32'h10408000;
      12543: inst = 32'hc4051d5;
      12544: inst = 32'h8220000;
      12545: inst = 32'h10408000;
      12546: inst = 32'hc4051d6;
      12547: inst = 32'h8220000;
      12548: inst = 32'h10408000;
      12549: inst = 32'hc4051d7;
      12550: inst = 32'h8220000;
      12551: inst = 32'h10408000;
      12552: inst = 32'hc4051d8;
      12553: inst = 32'h8220000;
      12554: inst = 32'h10408000;
      12555: inst = 32'hc4051d9;
      12556: inst = 32'h8220000;
      12557: inst = 32'h10408000;
      12558: inst = 32'hc4051da;
      12559: inst = 32'h8220000;
      12560: inst = 32'h10408000;
      12561: inst = 32'hc4051db;
      12562: inst = 32'h8220000;
      12563: inst = 32'h10408000;
      12564: inst = 32'hc4051dc;
      12565: inst = 32'h8220000;
      12566: inst = 32'h10408000;
      12567: inst = 32'hc4051dd;
      12568: inst = 32'h8220000;
      12569: inst = 32'h10408000;
      12570: inst = 32'hc4051de;
      12571: inst = 32'h8220000;
      12572: inst = 32'h10408000;
      12573: inst = 32'hc405230;
      12574: inst = 32'h8220000;
      12575: inst = 32'h10408000;
      12576: inst = 32'hc405231;
      12577: inst = 32'h8220000;
      12578: inst = 32'h10408000;
      12579: inst = 32'hc405232;
      12580: inst = 32'h8220000;
      12581: inst = 32'h10408000;
      12582: inst = 32'hc405233;
      12583: inst = 32'h8220000;
      12584: inst = 32'h10408000;
      12585: inst = 32'hc405234;
      12586: inst = 32'h8220000;
      12587: inst = 32'h10408000;
      12588: inst = 32'hc405235;
      12589: inst = 32'h8220000;
      12590: inst = 32'h10408000;
      12591: inst = 32'hc405236;
      12592: inst = 32'h8220000;
      12593: inst = 32'h10408000;
      12594: inst = 32'hc405237;
      12595: inst = 32'h8220000;
      12596: inst = 32'h10408000;
      12597: inst = 32'hc405238;
      12598: inst = 32'h8220000;
      12599: inst = 32'h10408000;
      12600: inst = 32'hc405239;
      12601: inst = 32'h8220000;
      12602: inst = 32'h10408000;
      12603: inst = 32'hc40523a;
      12604: inst = 32'h8220000;
      12605: inst = 32'h10408000;
      12606: inst = 32'hc40523b;
      12607: inst = 32'h8220000;
      12608: inst = 32'h10408000;
      12609: inst = 32'hc40523c;
      12610: inst = 32'h8220000;
      12611: inst = 32'h10408000;
      12612: inst = 32'hc40523d;
      12613: inst = 32'h8220000;
      12614: inst = 32'h10408000;
      12615: inst = 32'hc40523e;
      12616: inst = 32'h8220000;
      12617: inst = 32'h10408000;
      12618: inst = 32'hc405290;
      12619: inst = 32'h8220000;
      12620: inst = 32'h10408000;
      12621: inst = 32'hc405291;
      12622: inst = 32'h8220000;
      12623: inst = 32'h10408000;
      12624: inst = 32'hc405292;
      12625: inst = 32'h8220000;
      12626: inst = 32'h10408000;
      12627: inst = 32'hc405293;
      12628: inst = 32'h8220000;
      12629: inst = 32'h10408000;
      12630: inst = 32'hc405294;
      12631: inst = 32'h8220000;
      12632: inst = 32'h10408000;
      12633: inst = 32'hc405295;
      12634: inst = 32'h8220000;
      12635: inst = 32'h10408000;
      12636: inst = 32'hc405296;
      12637: inst = 32'h8220000;
      12638: inst = 32'h10408000;
      12639: inst = 32'hc405297;
      12640: inst = 32'h8220000;
      12641: inst = 32'h10408000;
      12642: inst = 32'hc405298;
      12643: inst = 32'h8220000;
      12644: inst = 32'h10408000;
      12645: inst = 32'hc405299;
      12646: inst = 32'h8220000;
      12647: inst = 32'h10408000;
      12648: inst = 32'hc40529a;
      12649: inst = 32'h8220000;
      12650: inst = 32'h10408000;
      12651: inst = 32'hc40529b;
      12652: inst = 32'h8220000;
      12653: inst = 32'h10408000;
      12654: inst = 32'hc40529c;
      12655: inst = 32'h8220000;
      12656: inst = 32'h10408000;
      12657: inst = 32'hc40529d;
      12658: inst = 32'h8220000;
      12659: inst = 32'h10408000;
      12660: inst = 32'hc40529e;
      12661: inst = 32'h8220000;
      12662: inst = 32'hc20ef7c;
      12663: inst = 32'h10408000;
      12664: inst = 32'hc404932;
      12665: inst = 32'h8220000;
      12666: inst = 32'h10408000;
      12667: inst = 32'hc404933;
      12668: inst = 32'h8220000;
      12669: inst = 32'h10408000;
      12670: inst = 32'hc404934;
      12671: inst = 32'h8220000;
      12672: inst = 32'h10408000;
      12673: inst = 32'hc404935;
      12674: inst = 32'h8220000;
      12675: inst = 32'h10408000;
      12676: inst = 32'hc404993;
      12677: inst = 32'h8220000;
      12678: inst = 32'h10408000;
      12679: inst = 32'hc404994;
      12680: inst = 32'h8220000;
      12681: inst = 32'h10408000;
      12682: inst = 32'hc404995;
      12683: inst = 32'h8220000;
      12684: inst = 32'h10408000;
      12685: inst = 32'hc4049f3;
      12686: inst = 32'h8220000;
      12687: inst = 32'h10408000;
      12688: inst = 32'hc4049f4;
      12689: inst = 32'h8220000;
      12690: inst = 32'h10408000;
      12691: inst = 32'hc4049f5;
      12692: inst = 32'h8220000;
      12693: inst = 32'h10408000;
      12694: inst = 32'hc404a53;
      12695: inst = 32'h8220000;
      12696: inst = 32'h10408000;
      12697: inst = 32'hc404a54;
      12698: inst = 32'h8220000;
      12699: inst = 32'h10408000;
      12700: inst = 32'hc404a55;
      12701: inst = 32'h8220000;
      12702: inst = 32'h10408000;
      12703: inst = 32'hc404ab2;
      12704: inst = 32'h8220000;
      12705: inst = 32'h10408000;
      12706: inst = 32'hc404ab3;
      12707: inst = 32'h8220000;
      12708: inst = 32'h10408000;
      12709: inst = 32'hc404ab5;
      12710: inst = 32'h8220000;
      12711: inst = 32'h10408000;
      12712: inst = 32'hc404b12;
      12713: inst = 32'h8220000;
      12714: inst = 32'h10408000;
      12715: inst = 32'hc404b13;
      12716: inst = 32'h8220000;
      12717: inst = 32'h10408000;
      12718: inst = 32'hc404b15;
      12719: inst = 32'h8220000;
      12720: inst = 32'h10408000;
      12721: inst = 32'hc404b72;
      12722: inst = 32'h8220000;
      12723: inst = 32'h10408000;
      12724: inst = 32'hc404b73;
      12725: inst = 32'h8220000;
      12726: inst = 32'h10408000;
      12727: inst = 32'hc404b74;
      12728: inst = 32'h8220000;
      12729: inst = 32'h10408000;
      12730: inst = 32'hc404b75;
      12731: inst = 32'h8220000;
      12732: inst = 32'hc20eed7;
      12733: inst = 32'h10408000;
      12734: inst = 32'hc404a08;
      12735: inst = 32'h8220000;
      12736: inst = 32'h10408000;
      12737: inst = 32'hc404a0e;
      12738: inst = 32'h8220000;
      12739: inst = 32'hc20e6fa;
      12740: inst = 32'h10408000;
      12741: inst = 32'hc404a09;
      12742: inst = 32'h8220000;
      12743: inst = 32'h10408000;
      12744: inst = 32'hc404a0d;
      12745: inst = 32'h8220000;
      12746: inst = 32'h10408000;
      12747: inst = 32'hc404be7;
      12748: inst = 32'h8220000;
      12749: inst = 32'hc20e6fb;
      12750: inst = 32'h10408000;
      12751: inst = 32'hc404a0a;
      12752: inst = 32'h8220000;
      12753: inst = 32'h10408000;
      12754: inst = 32'hc404a0c;
      12755: inst = 32'h8220000;
      12756: inst = 32'h10408000;
      12757: inst = 32'hc404ac7;
      12758: inst = 32'h8220000;
      12759: inst = 32'h10408000;
      12760: inst = 32'hc404acf;
      12761: inst = 32'h8220000;
      12762: inst = 32'h10408000;
      12763: inst = 32'hc404b87;
      12764: inst = 32'h8220000;
      12765: inst = 32'h10408000;
      12766: inst = 32'hc404b8f;
      12767: inst = 32'h8220000;
      12768: inst = 32'h10408000;
      12769: inst = 32'hc404c4d;
      12770: inst = 32'h8220000;
      12771: inst = 32'hc20defb;
      12772: inst = 32'h10408000;
      12773: inst = 32'hc404a0b;
      12774: inst = 32'h8220000;
      12775: inst = 32'h10408000;
      12776: inst = 32'hc404a68;
      12777: inst = 32'h8220000;
      12778: inst = 32'h10408000;
      12779: inst = 32'hc404a69;
      12780: inst = 32'h8220000;
      12781: inst = 32'h10408000;
      12782: inst = 32'hc404a6a;
      12783: inst = 32'h8220000;
      12784: inst = 32'h10408000;
      12785: inst = 32'hc404a6b;
      12786: inst = 32'h8220000;
      12787: inst = 32'h10408000;
      12788: inst = 32'hc404a6c;
      12789: inst = 32'h8220000;
      12790: inst = 32'h10408000;
      12791: inst = 32'hc404a6d;
      12792: inst = 32'h8220000;
      12793: inst = 32'h10408000;
      12794: inst = 32'hc404a6e;
      12795: inst = 32'h8220000;
      12796: inst = 32'h10408000;
      12797: inst = 32'hc404ac8;
      12798: inst = 32'h8220000;
      12799: inst = 32'h10408000;
      12800: inst = 32'hc404ac9;
      12801: inst = 32'h8220000;
      12802: inst = 32'h10408000;
      12803: inst = 32'hc404aca;
      12804: inst = 32'h8220000;
      12805: inst = 32'h10408000;
      12806: inst = 32'hc404acb;
      12807: inst = 32'h8220000;
      12808: inst = 32'h10408000;
      12809: inst = 32'hc404acc;
      12810: inst = 32'h8220000;
      12811: inst = 32'h10408000;
      12812: inst = 32'hc404acd;
      12813: inst = 32'h8220000;
      12814: inst = 32'h10408000;
      12815: inst = 32'hc404ace;
      12816: inst = 32'h8220000;
      12817: inst = 32'h10408000;
      12818: inst = 32'hc404b27;
      12819: inst = 32'h8220000;
      12820: inst = 32'h10408000;
      12821: inst = 32'hc404b2a;
      12822: inst = 32'h8220000;
      12823: inst = 32'h10408000;
      12824: inst = 32'hc404b2d;
      12825: inst = 32'h8220000;
      12826: inst = 32'h10408000;
      12827: inst = 32'hc404b2e;
      12828: inst = 32'h8220000;
      12829: inst = 32'h10408000;
      12830: inst = 32'hc404b2f;
      12831: inst = 32'h8220000;
      12832: inst = 32'h10408000;
      12833: inst = 32'hc404b8a;
      12834: inst = 32'h8220000;
      12835: inst = 32'h10408000;
      12836: inst = 32'hc404b8d;
      12837: inst = 32'h8220000;
      12838: inst = 32'h10408000;
      12839: inst = 32'hc404b8e;
      12840: inst = 32'h8220000;
      12841: inst = 32'h10408000;
      12842: inst = 32'hc404be8;
      12843: inst = 32'h8220000;
      12844: inst = 32'h10408000;
      12845: inst = 32'hc404be9;
      12846: inst = 32'h8220000;
      12847: inst = 32'h10408000;
      12848: inst = 32'hc404bea;
      12849: inst = 32'h8220000;
      12850: inst = 32'h10408000;
      12851: inst = 32'hc404beb;
      12852: inst = 32'h8220000;
      12853: inst = 32'h10408000;
      12854: inst = 32'hc404bec;
      12855: inst = 32'h8220000;
      12856: inst = 32'h10408000;
      12857: inst = 32'hc404bed;
      12858: inst = 32'h8220000;
      12859: inst = 32'h10408000;
      12860: inst = 32'hc404bee;
      12861: inst = 32'h8220000;
      12862: inst = 32'h10408000;
      12863: inst = 32'hc404c49;
      12864: inst = 32'h8220000;
      12865: inst = 32'h10408000;
      12866: inst = 32'hc404c4b;
      12867: inst = 32'h8220000;
      12868: inst = 32'h10408000;
      12869: inst = 32'hc404ca9;
      12870: inst = 32'h8220000;
      12871: inst = 32'h10408000;
      12872: inst = 32'hc404cab;
      12873: inst = 32'h8220000;
      12874: inst = 32'hc20eed8;
      12875: inst = 32'h10408000;
      12876: inst = 32'hc404a67;
      12877: inst = 32'h8220000;
      12878: inst = 32'h10408000;
      12879: inst = 32'hc404a6f;
      12880: inst = 32'h8220000;
      12881: inst = 32'hc204a69;
      12882: inst = 32'h10408000;
      12883: inst = 32'hc404b28;
      12884: inst = 32'h8220000;
      12885: inst = 32'h10408000;
      12886: inst = 32'hc404b29;
      12887: inst = 32'h8220000;
      12888: inst = 32'h10408000;
      12889: inst = 32'hc404b2b;
      12890: inst = 32'h8220000;
      12891: inst = 32'h10408000;
      12892: inst = 32'hc404b2c;
      12893: inst = 32'h8220000;
      12894: inst = 32'h10408000;
      12895: inst = 32'hc404b88;
      12896: inst = 32'h8220000;
      12897: inst = 32'h10408000;
      12898: inst = 32'hc404b89;
      12899: inst = 32'h8220000;
      12900: inst = 32'h10408000;
      12901: inst = 32'hc404b8b;
      12902: inst = 32'h8220000;
      12903: inst = 32'h10408000;
      12904: inst = 32'hc404b8c;
      12905: inst = 32'h8220000;
      12906: inst = 32'h10408000;
      12907: inst = 32'hc404c48;
      12908: inst = 32'h8220000;
      12909: inst = 32'h10408000;
      12910: inst = 32'hc404c4a;
      12911: inst = 32'h8220000;
      12912: inst = 32'h10408000;
      12913: inst = 32'hc404c4c;
      12914: inst = 32'h8220000;
      12915: inst = 32'h10408000;
      12916: inst = 32'hc404ca8;
      12917: inst = 32'h8220000;
      12918: inst = 32'h10408000;
      12919: inst = 32'hc404caa;
      12920: inst = 32'h8220000;
      12921: inst = 32'h10408000;
      12922: inst = 32'hc404cac;
      12923: inst = 32'h8220000;
      12924: inst = 32'h10408000;
      12925: inst = 32'hc405085;
      12926: inst = 32'h8220000;
      12927: inst = 32'h10408000;
      12928: inst = 32'hc40509a;
      12929: inst = 32'h8220000;
      12930: inst = 32'h10408000;
      12931: inst = 32'hc4050e4;
      12932: inst = 32'h8220000;
      12933: inst = 32'h10408000;
      12934: inst = 32'hc4050e5;
      12935: inst = 32'h8220000;
      12936: inst = 32'h10408000;
      12937: inst = 32'hc4050fa;
      12938: inst = 32'h8220000;
      12939: inst = 32'h10408000;
      12940: inst = 32'hc4050fb;
      12941: inst = 32'h8220000;
      12942: inst = 32'h10408000;
      12943: inst = 32'hc405143;
      12944: inst = 32'h8220000;
      12945: inst = 32'h10408000;
      12946: inst = 32'hc405144;
      12947: inst = 32'h8220000;
      12948: inst = 32'h10408000;
      12949: inst = 32'hc405145;
      12950: inst = 32'h8220000;
      12951: inst = 32'h10408000;
      12952: inst = 32'hc40515a;
      12953: inst = 32'h8220000;
      12954: inst = 32'h10408000;
      12955: inst = 32'hc40515b;
      12956: inst = 32'h8220000;
      12957: inst = 32'h10408000;
      12958: inst = 32'hc40515c;
      12959: inst = 32'h8220000;
      12960: inst = 32'h10408000;
      12961: inst = 32'hc4051a2;
      12962: inst = 32'h8220000;
      12963: inst = 32'h10408000;
      12964: inst = 32'hc4051a3;
      12965: inst = 32'h8220000;
      12966: inst = 32'h10408000;
      12967: inst = 32'hc4051a4;
      12968: inst = 32'h8220000;
      12969: inst = 32'h10408000;
      12970: inst = 32'hc4051a5;
      12971: inst = 32'h8220000;
      12972: inst = 32'h10408000;
      12973: inst = 32'hc4051ba;
      12974: inst = 32'h8220000;
      12975: inst = 32'h10408000;
      12976: inst = 32'hc4051bb;
      12977: inst = 32'h8220000;
      12978: inst = 32'h10408000;
      12979: inst = 32'hc4051bc;
      12980: inst = 32'h8220000;
      12981: inst = 32'h10408000;
      12982: inst = 32'hc4051bd;
      12983: inst = 32'h8220000;
      12984: inst = 32'h10408000;
      12985: inst = 32'hc405202;
      12986: inst = 32'h8220000;
      12987: inst = 32'h10408000;
      12988: inst = 32'hc405203;
      12989: inst = 32'h8220000;
      12990: inst = 32'h10408000;
      12991: inst = 32'hc405204;
      12992: inst = 32'h8220000;
      12993: inst = 32'h10408000;
      12994: inst = 32'hc405205;
      12995: inst = 32'h8220000;
      12996: inst = 32'h10408000;
      12997: inst = 32'hc40521a;
      12998: inst = 32'h8220000;
      12999: inst = 32'h10408000;
      13000: inst = 32'hc40521b;
      13001: inst = 32'h8220000;
      13002: inst = 32'h10408000;
      13003: inst = 32'hc40521c;
      13004: inst = 32'h8220000;
      13005: inst = 32'h10408000;
      13006: inst = 32'hc40521d;
      13007: inst = 32'h8220000;
      13008: inst = 32'h10408000;
      13009: inst = 32'hc405262;
      13010: inst = 32'h8220000;
      13011: inst = 32'h10408000;
      13012: inst = 32'hc405263;
      13013: inst = 32'h8220000;
      13014: inst = 32'h10408000;
      13015: inst = 32'hc405264;
      13016: inst = 32'h8220000;
      13017: inst = 32'h10408000;
      13018: inst = 32'hc405265;
      13019: inst = 32'h8220000;
      13020: inst = 32'h10408000;
      13021: inst = 32'hc40527a;
      13022: inst = 32'h8220000;
      13023: inst = 32'h10408000;
      13024: inst = 32'hc40527b;
      13025: inst = 32'h8220000;
      13026: inst = 32'h10408000;
      13027: inst = 32'hc40527c;
      13028: inst = 32'h8220000;
      13029: inst = 32'h10408000;
      13030: inst = 32'hc40527d;
      13031: inst = 32'h8220000;
      13032: inst = 32'h10408000;
      13033: inst = 32'hc4052c2;
      13034: inst = 32'h8220000;
      13035: inst = 32'h10408000;
      13036: inst = 32'hc4052c3;
      13037: inst = 32'h8220000;
      13038: inst = 32'h10408000;
      13039: inst = 32'hc4052c4;
      13040: inst = 32'h8220000;
      13041: inst = 32'h10408000;
      13042: inst = 32'hc4052db;
      13043: inst = 32'h8220000;
      13044: inst = 32'h10408000;
      13045: inst = 32'hc4052dc;
      13046: inst = 32'h8220000;
      13047: inst = 32'h10408000;
      13048: inst = 32'hc4052dd;
      13049: inst = 32'h8220000;
      13050: inst = 32'h10408000;
      13051: inst = 32'hc405322;
      13052: inst = 32'h8220000;
      13053: inst = 32'h10408000;
      13054: inst = 32'hc405323;
      13055: inst = 32'h8220000;
      13056: inst = 32'h10408000;
      13057: inst = 32'hc405324;
      13058: inst = 32'h8220000;
      13059: inst = 32'h10408000;
      13060: inst = 32'hc40533b;
      13061: inst = 32'h8220000;
      13062: inst = 32'h10408000;
      13063: inst = 32'hc40533c;
      13064: inst = 32'h8220000;
      13065: inst = 32'h10408000;
      13066: inst = 32'hc40533d;
      13067: inst = 32'h8220000;
      13068: inst = 32'h10408000;
      13069: inst = 32'hc40537f;
      13070: inst = 32'h8220000;
      13071: inst = 32'h10408000;
      13072: inst = 32'hc405382;
      13073: inst = 32'h8220000;
      13074: inst = 32'h10408000;
      13075: inst = 32'hc405383;
      13076: inst = 32'h8220000;
      13077: inst = 32'h10408000;
      13078: inst = 32'hc405384;
      13079: inst = 32'h8220000;
      13080: inst = 32'h10408000;
      13081: inst = 32'hc40539b;
      13082: inst = 32'h8220000;
      13083: inst = 32'h10408000;
      13084: inst = 32'hc40539c;
      13085: inst = 32'h8220000;
      13086: inst = 32'h10408000;
      13087: inst = 32'hc40539d;
      13088: inst = 32'h8220000;
      13089: inst = 32'h10408000;
      13090: inst = 32'hc4053a0;
      13091: inst = 32'h8220000;
      13092: inst = 32'h10408000;
      13093: inst = 32'hc4053de;
      13094: inst = 32'h8220000;
      13095: inst = 32'h10408000;
      13096: inst = 32'hc4053df;
      13097: inst = 32'h8220000;
      13098: inst = 32'h10408000;
      13099: inst = 32'hc4053e2;
      13100: inst = 32'h8220000;
      13101: inst = 32'h10408000;
      13102: inst = 32'hc4053e3;
      13103: inst = 32'h8220000;
      13104: inst = 32'h10408000;
      13105: inst = 32'hc4053fc;
      13106: inst = 32'h8220000;
      13107: inst = 32'h10408000;
      13108: inst = 32'hc4053fd;
      13109: inst = 32'h8220000;
      13110: inst = 32'h10408000;
      13111: inst = 32'hc405400;
      13112: inst = 32'h8220000;
      13113: inst = 32'h10408000;
      13114: inst = 32'hc405401;
      13115: inst = 32'h8220000;
      13116: inst = 32'h10408000;
      13117: inst = 32'hc40543d;
      13118: inst = 32'h8220000;
      13119: inst = 32'h10408000;
      13120: inst = 32'hc40543e;
      13121: inst = 32'h8220000;
      13122: inst = 32'h10408000;
      13123: inst = 32'hc40543f;
      13124: inst = 32'h8220000;
      13125: inst = 32'h10408000;
      13126: inst = 32'hc405442;
      13127: inst = 32'h8220000;
      13128: inst = 32'h10408000;
      13129: inst = 32'hc405443;
      13130: inst = 32'h8220000;
      13131: inst = 32'h10408000;
      13132: inst = 32'hc40545c;
      13133: inst = 32'h8220000;
      13134: inst = 32'h10408000;
      13135: inst = 32'hc40545d;
      13136: inst = 32'h8220000;
      13137: inst = 32'h10408000;
      13138: inst = 32'hc405460;
      13139: inst = 32'h8220000;
      13140: inst = 32'h10408000;
      13141: inst = 32'hc405461;
      13142: inst = 32'h8220000;
      13143: inst = 32'h10408000;
      13144: inst = 32'hc405462;
      13145: inst = 32'h8220000;
      13146: inst = 32'h10408000;
      13147: inst = 32'hc40549d;
      13148: inst = 32'h8220000;
      13149: inst = 32'h10408000;
      13150: inst = 32'hc40549e;
      13151: inst = 32'h8220000;
      13152: inst = 32'h10408000;
      13153: inst = 32'hc4054a0;
      13154: inst = 32'h8220000;
      13155: inst = 32'h10408000;
      13156: inst = 32'hc4054a1;
      13157: inst = 32'h8220000;
      13158: inst = 32'h10408000;
      13159: inst = 32'hc4054a2;
      13160: inst = 32'h8220000;
      13161: inst = 32'h10408000;
      13162: inst = 32'hc4054a3;
      13163: inst = 32'h8220000;
      13164: inst = 32'h10408000;
      13165: inst = 32'hc4054bc;
      13166: inst = 32'h8220000;
      13167: inst = 32'h10408000;
      13168: inst = 32'hc4054bd;
      13169: inst = 32'h8220000;
      13170: inst = 32'h10408000;
      13171: inst = 32'hc4054be;
      13172: inst = 32'h8220000;
      13173: inst = 32'h10408000;
      13174: inst = 32'hc4054bf;
      13175: inst = 32'h8220000;
      13176: inst = 32'h10408000;
      13177: inst = 32'hc4054c1;
      13178: inst = 32'h8220000;
      13179: inst = 32'h10408000;
      13180: inst = 32'hc4054c2;
      13181: inst = 32'h8220000;
      13182: inst = 32'h10408000;
      13183: inst = 32'hc4054fc;
      13184: inst = 32'h8220000;
      13185: inst = 32'h10408000;
      13186: inst = 32'hc4054fd;
      13187: inst = 32'h8220000;
      13188: inst = 32'h10408000;
      13189: inst = 32'hc4054fe;
      13190: inst = 32'h8220000;
      13191: inst = 32'h10408000;
      13192: inst = 32'hc405502;
      13193: inst = 32'h8220000;
      13194: inst = 32'h10408000;
      13195: inst = 32'hc40551d;
      13196: inst = 32'h8220000;
      13197: inst = 32'h10408000;
      13198: inst = 32'hc405521;
      13199: inst = 32'h8220000;
      13200: inst = 32'h10408000;
      13201: inst = 32'hc405522;
      13202: inst = 32'h8220000;
      13203: inst = 32'h10408000;
      13204: inst = 32'hc405523;
      13205: inst = 32'h8220000;
      13206: inst = 32'h10408000;
      13207: inst = 32'hc40555b;
      13208: inst = 32'h8220000;
      13209: inst = 32'h10408000;
      13210: inst = 32'hc40555c;
      13211: inst = 32'h8220000;
      13212: inst = 32'h10408000;
      13213: inst = 32'hc40555d;
      13214: inst = 32'h8220000;
      13215: inst = 32'h10408000;
      13216: inst = 32'hc405562;
      13217: inst = 32'h8220000;
      13218: inst = 32'h10408000;
      13219: inst = 32'hc40557d;
      13220: inst = 32'h8220000;
      13221: inst = 32'h10408000;
      13222: inst = 32'hc405582;
      13223: inst = 32'h8220000;
      13224: inst = 32'h10408000;
      13225: inst = 32'hc405583;
      13226: inst = 32'h8220000;
      13227: inst = 32'h10408000;
      13228: inst = 32'hc405584;
      13229: inst = 32'h8220000;
      13230: inst = 32'h10408000;
      13231: inst = 32'hc4055ba;
      13232: inst = 32'h8220000;
      13233: inst = 32'h10408000;
      13234: inst = 32'hc4055bb;
      13235: inst = 32'h8220000;
      13236: inst = 32'h10408000;
      13237: inst = 32'hc4055bc;
      13238: inst = 32'h8220000;
      13239: inst = 32'h10408000;
      13240: inst = 32'hc4055bd;
      13241: inst = 32'h8220000;
      13242: inst = 32'h10408000;
      13243: inst = 32'hc4055c2;
      13244: inst = 32'h8220000;
      13245: inst = 32'h10408000;
      13246: inst = 32'hc4055dd;
      13247: inst = 32'h8220000;
      13248: inst = 32'h10408000;
      13249: inst = 32'hc4055e2;
      13250: inst = 32'h8220000;
      13251: inst = 32'h10408000;
      13252: inst = 32'hc4055e3;
      13253: inst = 32'h8220000;
      13254: inst = 32'h10408000;
      13255: inst = 32'hc4055e4;
      13256: inst = 32'h8220000;
      13257: inst = 32'h10408000;
      13258: inst = 32'hc4055e5;
      13259: inst = 32'h8220000;
      13260: inst = 32'h10408000;
      13261: inst = 32'hc40561a;
      13262: inst = 32'h8220000;
      13263: inst = 32'h10408000;
      13264: inst = 32'hc40561b;
      13265: inst = 32'h8220000;
      13266: inst = 32'h10408000;
      13267: inst = 32'hc40561c;
      13268: inst = 32'h8220000;
      13269: inst = 32'h10408000;
      13270: inst = 32'hc40561d;
      13271: inst = 32'h8220000;
      13272: inst = 32'h10408000;
      13273: inst = 32'hc405642;
      13274: inst = 32'h8220000;
      13275: inst = 32'h10408000;
      13276: inst = 32'hc405643;
      13277: inst = 32'h8220000;
      13278: inst = 32'h10408000;
      13279: inst = 32'hc405644;
      13280: inst = 32'h8220000;
      13281: inst = 32'h10408000;
      13282: inst = 32'hc405645;
      13283: inst = 32'h8220000;
      13284: inst = 32'h10408000;
      13285: inst = 32'hc405679;
      13286: inst = 32'h8220000;
      13287: inst = 32'h10408000;
      13288: inst = 32'hc40567a;
      13289: inst = 32'h8220000;
      13290: inst = 32'h10408000;
      13291: inst = 32'hc40567b;
      13292: inst = 32'h8220000;
      13293: inst = 32'h10408000;
      13294: inst = 32'hc40567c;
      13295: inst = 32'h8220000;
      13296: inst = 32'h10408000;
      13297: inst = 32'hc4056a3;
      13298: inst = 32'h8220000;
      13299: inst = 32'h10408000;
      13300: inst = 32'hc4056a4;
      13301: inst = 32'h8220000;
      13302: inst = 32'h10408000;
      13303: inst = 32'hc4056a5;
      13304: inst = 32'h8220000;
      13305: inst = 32'h10408000;
      13306: inst = 32'hc4056a6;
      13307: inst = 32'h8220000;
      13308: inst = 32'hc20e6d9;
      13309: inst = 32'h10408000;
      13310: inst = 32'hc404bef;
      13311: inst = 32'h8220000;
      13312: inst = 32'h10408000;
      13313: inst = 32'hc404c4e;
      13314: inst = 32'h8220000;
      13315: inst = 32'hc20eeb7;
      13316: inst = 32'h10408000;
      13317: inst = 32'hc404c47;
      13318: inst = 32'h8220000;
      13319: inst = 32'hc20d615;
      13320: inst = 32'h10408000;
      13321: inst = 32'hc404ca2;
      13322: inst = 32'h8220000;
      13323: inst = 32'h10408000;
      13324: inst = 32'hc404d00;
      13325: inst = 32'h8220000;
      13326: inst = 32'hc209c91;
      13327: inst = 32'h10408000;
      13328: inst = 32'hc404ca3;
      13329: inst = 32'h8220000;
      13330: inst = 32'h10408000;
      13331: inst = 32'hc404d01;
      13332: inst = 32'h8220000;
      13333: inst = 32'hc207bf0;
      13334: inst = 32'h10408000;
      13335: inst = 32'hc404ca4;
      13336: inst = 32'h8220000;
      13337: inst = 32'h10408000;
      13338: inst = 32'hc404ca5;
      13339: inst = 32'h8220000;
      13340: inst = 32'h10408000;
      13341: inst = 32'hc404ca6;
      13342: inst = 32'h8220000;
      13343: inst = 32'h10408000;
      13344: inst = 32'hc404ca7;
      13345: inst = 32'h8220000;
      13346: inst = 32'h10408000;
      13347: inst = 32'hc404d02;
      13348: inst = 32'h8220000;
      13349: inst = 32'h10408000;
      13350: inst = 32'hc404d03;
      13351: inst = 32'h8220000;
      13352: inst = 32'h10408000;
      13353: inst = 32'hc404d04;
      13354: inst = 32'h8220000;
      13355: inst = 32'h10408000;
      13356: inst = 32'hc404d05;
      13357: inst = 32'h8220000;
      13358: inst = 32'h10408000;
      13359: inst = 32'hc404d06;
      13360: inst = 32'h8220000;
      13361: inst = 32'h10408000;
      13362: inst = 32'hc404d07;
      13363: inst = 32'h8220000;
      13364: inst = 32'h10408000;
      13365: inst = 32'hc404d08;
      13366: inst = 32'h8220000;
      13367: inst = 32'h10408000;
      13368: inst = 32'hc404d09;
      13369: inst = 32'h8220000;
      13370: inst = 32'h10408000;
      13371: inst = 32'hc404d0a;
      13372: inst = 32'h8220000;
      13373: inst = 32'h10408000;
      13374: inst = 32'hc404d0b;
      13375: inst = 32'h8220000;
      13376: inst = 32'h10408000;
      13377: inst = 32'hc404d0c;
      13378: inst = 32'h8220000;
      13379: inst = 32'h10408000;
      13380: inst = 32'hc404d0d;
      13381: inst = 32'h8220000;
      13382: inst = 32'h10408000;
      13383: inst = 32'hc404d0e;
      13384: inst = 32'h8220000;
      13385: inst = 32'h10408000;
      13386: inst = 32'hc404d0f;
      13387: inst = 32'h8220000;
      13388: inst = 32'h10408000;
      13389: inst = 32'hc404d10;
      13390: inst = 32'h8220000;
      13391: inst = 32'h10408000;
      13392: inst = 32'hc404d11;
      13393: inst = 32'h8220000;
      13394: inst = 32'h10408000;
      13395: inst = 32'hc404d12;
      13396: inst = 32'h8220000;
      13397: inst = 32'h10408000;
      13398: inst = 32'hc404d13;
      13399: inst = 32'h8220000;
      13400: inst = 32'h10408000;
      13401: inst = 32'hc404d14;
      13402: inst = 32'h8220000;
      13403: inst = 32'h10408000;
      13404: inst = 32'hc4055c3;
      13405: inst = 32'h8220000;
      13406: inst = 32'h10408000;
      13407: inst = 32'hc4055dc;
      13408: inst = 32'h8220000;
      13409: inst = 32'hc20ad55;
      13410: inst = 32'h10408000;
      13411: inst = 32'hc404cad;
      13412: inst = 32'h8220000;
      13413: inst = 32'hc208410;
      13414: inst = 32'h10408000;
      13415: inst = 32'hc404cae;
      13416: inst = 32'h8220000;
      13417: inst = 32'h10408000;
      13418: inst = 32'hc404caf;
      13419: inst = 32'h8220000;
      13420: inst = 32'h10408000;
      13421: inst = 32'hc404cb0;
      13422: inst = 32'h8220000;
      13423: inst = 32'h10408000;
      13424: inst = 32'hc404cb1;
      13425: inst = 32'h8220000;
      13426: inst = 32'h10408000;
      13427: inst = 32'hc404cb2;
      13428: inst = 32'h8220000;
      13429: inst = 32'h10408000;
      13430: inst = 32'hc404cb3;
      13431: inst = 32'h8220000;
      13432: inst = 32'h10408000;
      13433: inst = 32'hc404cb4;
      13434: inst = 32'h8220000;
      13435: inst = 32'h10408000;
      13436: inst = 32'hc404cb5;
      13437: inst = 32'h8220000;
      13438: inst = 32'h10408000;
      13439: inst = 32'hc40537d;
      13440: inst = 32'h8220000;
      13441: inst = 32'h10408000;
      13442: inst = 32'hc405385;
      13443: inst = 32'h8220000;
      13444: inst = 32'h10408000;
      13445: inst = 32'hc40539a;
      13446: inst = 32'h8220000;
      13447: inst = 32'h10408000;
      13448: inst = 32'hc4053a2;
      13449: inst = 32'h8220000;
      13450: inst = 32'h10408000;
      13451: inst = 32'hc4054a4;
      13452: inst = 32'h8220000;
      13453: inst = 32'h10408000;
      13454: inst = 32'hc4054bb;
      13455: inst = 32'h8220000;
      13456: inst = 32'h10408000;
      13457: inst = 32'hc405741;
      13458: inst = 32'h8220000;
      13459: inst = 32'h10408000;
      13460: inst = 32'hc40575e;
      13461: inst = 32'h8220000;
      13462: inst = 32'hc209470;
      13463: inst = 32'h10408000;
      13464: inst = 32'hc404cb6;
      13465: inst = 32'h8220000;
      13466: inst = 32'h10408000;
      13467: inst = 32'hc404d15;
      13468: inst = 32'h8220000;
      13469: inst = 32'hc20a534;
      13470: inst = 32'h10408000;
      13471: inst = 32'hc404cfb;
      13472: inst = 32'h8220000;
      13473: inst = 32'hc208c51;
      13474: inst = 32'h10408000;
      13475: inst = 32'hc404cfc;
      13476: inst = 32'h8220000;
      13477: inst = 32'h10408000;
      13478: inst = 32'hc404cfd;
      13479: inst = 32'h8220000;
      13480: inst = 32'h10408000;
      13481: inst = 32'hc4053da;
      13482: inst = 32'h8220000;
      13483: inst = 32'h10408000;
      13484: inst = 32'hc4053dc;
      13485: inst = 32'h8220000;
      13486: inst = 32'h10408000;
      13487: inst = 32'hc405403;
      13488: inst = 32'h8220000;
      13489: inst = 32'h10408000;
      13490: inst = 32'hc405405;
      13491: inst = 32'h8220000;
      13492: inst = 32'h10408000;
      13493: inst = 32'hc4054fa;
      13494: inst = 32'h8220000;
      13495: inst = 32'h10408000;
      13496: inst = 32'hc405525;
      13497: inst = 32'h8220000;
      13498: inst = 32'h10408000;
      13499: inst = 32'hc405557;
      13500: inst = 32'h8220000;
      13501: inst = 32'h10408000;
      13502: inst = 32'hc40555f;
      13503: inst = 32'h8220000;
      13504: inst = 32'h10408000;
      13505: inst = 32'hc405580;
      13506: inst = 32'h8220000;
      13507: inst = 32'h10408000;
      13508: inst = 32'hc405588;
      13509: inst = 32'h8220000;
      13510: inst = 32'h10408000;
      13511: inst = 32'hc405618;
      13512: inst = 32'h8220000;
      13513: inst = 32'h10408000;
      13514: inst = 32'hc405627;
      13515: inst = 32'h8220000;
      13516: inst = 32'h10408000;
      13517: inst = 32'hc405638;
      13518: inst = 32'h8220000;
      13519: inst = 32'h10408000;
      13520: inst = 32'hc405647;
      13521: inst = 32'h8220000;
      13522: inst = 32'h10408000;
      13523: inst = 32'hc40570b;
      13524: inst = 32'h8220000;
      13525: inst = 32'hc206b6d;
      13526: inst = 32'h10408000;
      13527: inst = 32'hc404d16;
      13528: inst = 32'h8220000;
      13529: inst = 32'h10408000;
      13530: inst = 32'hc404d75;
      13531: inst = 32'h8220000;
      13532: inst = 32'h10408000;
      13533: inst = 32'hc404d76;
      13534: inst = 32'h8220000;
      13535: inst = 32'h10408000;
      13536: inst = 32'hc404dd5;
      13537: inst = 32'h8220000;
      13538: inst = 32'h10408000;
      13539: inst = 32'hc404dd6;
      13540: inst = 32'h8220000;
      13541: inst = 32'h10408000;
      13542: inst = 32'hc404e35;
      13543: inst = 32'h8220000;
      13544: inst = 32'h10408000;
      13545: inst = 32'hc404e36;
      13546: inst = 32'h8220000;
      13547: inst = 32'h10408000;
      13548: inst = 32'hc404e95;
      13549: inst = 32'h8220000;
      13550: inst = 32'h10408000;
      13551: inst = 32'hc404e96;
      13552: inst = 32'h8220000;
      13553: inst = 32'h10408000;
      13554: inst = 32'hc404ef5;
      13555: inst = 32'h8220000;
      13556: inst = 32'h10408000;
      13557: inst = 32'hc404ef6;
      13558: inst = 32'h8220000;
      13559: inst = 32'h10408000;
      13560: inst = 32'hc404f55;
      13561: inst = 32'h8220000;
      13562: inst = 32'h10408000;
      13563: inst = 32'hc404f56;
      13564: inst = 32'h8220000;
      13565: inst = 32'h10408000;
      13566: inst = 32'hc404fb5;
      13567: inst = 32'h8220000;
      13568: inst = 32'h10408000;
      13569: inst = 32'hc404fb6;
      13570: inst = 32'h8220000;
      13571: inst = 32'h10408000;
      13572: inst = 32'hc405015;
      13573: inst = 32'h8220000;
      13574: inst = 32'h10408000;
      13575: inst = 32'hc405016;
      13576: inst = 32'h8220000;
      13577: inst = 32'h10408000;
      13578: inst = 32'hc405075;
      13579: inst = 32'h8220000;
      13580: inst = 32'h10408000;
      13581: inst = 32'hc405076;
      13582: inst = 32'h8220000;
      13583: inst = 32'h10408000;
      13584: inst = 32'hc4050d5;
      13585: inst = 32'h8220000;
      13586: inst = 32'h10408000;
      13587: inst = 32'hc4050d6;
      13588: inst = 32'h8220000;
      13589: inst = 32'h10408000;
      13590: inst = 32'hc405135;
      13591: inst = 32'h8220000;
      13592: inst = 32'h10408000;
      13593: inst = 32'hc405136;
      13594: inst = 32'h8220000;
      13595: inst = 32'h10408000;
      13596: inst = 32'hc405195;
      13597: inst = 32'h8220000;
      13598: inst = 32'h10408000;
      13599: inst = 32'hc405196;
      13600: inst = 32'h8220000;
      13601: inst = 32'h10408000;
      13602: inst = 32'hc4051f5;
      13603: inst = 32'h8220000;
      13604: inst = 32'h10408000;
      13605: inst = 32'hc4051f6;
      13606: inst = 32'h8220000;
      13607: inst = 32'h10408000;
      13608: inst = 32'hc405255;
      13609: inst = 32'h8220000;
      13610: inst = 32'h10408000;
      13611: inst = 32'hc405256;
      13612: inst = 32'h8220000;
      13613: inst = 32'h10408000;
      13614: inst = 32'hc4052b5;
      13615: inst = 32'h8220000;
      13616: inst = 32'h10408000;
      13617: inst = 32'hc4052b6;
      13618: inst = 32'h8220000;
      13619: inst = 32'h10408000;
      13620: inst = 32'hc405325;
      13621: inst = 32'h8220000;
      13622: inst = 32'h10408000;
      13623: inst = 32'hc40533a;
      13624: inst = 32'h8220000;
      13625: inst = 32'hc20c638;
      13626: inst = 32'h10408000;
      13627: inst = 32'hc404d5b;
      13628: inst = 32'h8220000;
      13629: inst = 32'hc208c71;
      13630: inst = 32'h10408000;
      13631: inst = 32'hc404d60;
      13632: inst = 32'h8220000;
      13633: inst = 32'h10408000;
      13634: inst = 32'hc404d61;
      13635: inst = 32'h8220000;
      13636: inst = 32'h10408000;
      13637: inst = 32'hc404d62;
      13638: inst = 32'h8220000;
      13639: inst = 32'h10408000;
      13640: inst = 32'hc404d63;
      13641: inst = 32'h8220000;
      13642: inst = 32'h10408000;
      13643: inst = 32'hc404d64;
      13644: inst = 32'h8220000;
      13645: inst = 32'h10408000;
      13646: inst = 32'hc404d65;
      13647: inst = 32'h8220000;
      13648: inst = 32'h10408000;
      13649: inst = 32'hc404d66;
      13650: inst = 32'h8220000;
      13651: inst = 32'h10408000;
      13652: inst = 32'hc404d67;
      13653: inst = 32'h8220000;
      13654: inst = 32'h10408000;
      13655: inst = 32'hc404d68;
      13656: inst = 32'h8220000;
      13657: inst = 32'h10408000;
      13658: inst = 32'hc404d69;
      13659: inst = 32'h8220000;
      13660: inst = 32'h10408000;
      13661: inst = 32'hc404d6a;
      13662: inst = 32'h8220000;
      13663: inst = 32'h10408000;
      13664: inst = 32'hc404d6b;
      13665: inst = 32'h8220000;
      13666: inst = 32'h10408000;
      13667: inst = 32'hc404d6c;
      13668: inst = 32'h8220000;
      13669: inst = 32'h10408000;
      13670: inst = 32'hc404d6d;
      13671: inst = 32'h8220000;
      13672: inst = 32'h10408000;
      13673: inst = 32'hc404d6e;
      13674: inst = 32'h8220000;
      13675: inst = 32'h10408000;
      13676: inst = 32'hc404d6f;
      13677: inst = 32'h8220000;
      13678: inst = 32'h10408000;
      13679: inst = 32'hc404d70;
      13680: inst = 32'h8220000;
      13681: inst = 32'h10408000;
      13682: inst = 32'hc404d71;
      13683: inst = 32'h8220000;
      13684: inst = 32'h10408000;
      13685: inst = 32'hc404d72;
      13686: inst = 32'h8220000;
      13687: inst = 32'h10408000;
      13688: inst = 32'hc404d73;
      13689: inst = 32'h8220000;
      13690: inst = 32'h10408000;
      13691: inst = 32'hc404d74;
      13692: inst = 32'h8220000;
      13693: inst = 32'h10408000;
      13694: inst = 32'hc404dc0;
      13695: inst = 32'h8220000;
      13696: inst = 32'h10408000;
      13697: inst = 32'hc404dca;
      13698: inst = 32'h8220000;
      13699: inst = 32'h10408000;
      13700: inst = 32'hc404dd4;
      13701: inst = 32'h8220000;
      13702: inst = 32'h10408000;
      13703: inst = 32'hc404e20;
      13704: inst = 32'h8220000;
      13705: inst = 32'h10408000;
      13706: inst = 32'hc404e2a;
      13707: inst = 32'h8220000;
      13708: inst = 32'h10408000;
      13709: inst = 32'hc404e34;
      13710: inst = 32'h8220000;
      13711: inst = 32'h10408000;
      13712: inst = 32'hc404e80;
      13713: inst = 32'h8220000;
      13714: inst = 32'h10408000;
      13715: inst = 32'hc404e8a;
      13716: inst = 32'h8220000;
      13717: inst = 32'h10408000;
      13718: inst = 32'hc404e94;
      13719: inst = 32'h8220000;
      13720: inst = 32'h10408000;
      13721: inst = 32'hc404ee0;
      13722: inst = 32'h8220000;
      13723: inst = 32'h10408000;
      13724: inst = 32'hc404eea;
      13725: inst = 32'h8220000;
      13726: inst = 32'h10408000;
      13727: inst = 32'hc404ef4;
      13728: inst = 32'h8220000;
      13729: inst = 32'h10408000;
      13730: inst = 32'hc404f40;
      13731: inst = 32'h8220000;
      13732: inst = 32'h10408000;
      13733: inst = 32'hc404f4a;
      13734: inst = 32'h8220000;
      13735: inst = 32'h10408000;
      13736: inst = 32'hc404f54;
      13737: inst = 32'h8220000;
      13738: inst = 32'h10408000;
      13739: inst = 32'hc404fa0;
      13740: inst = 32'h8220000;
      13741: inst = 32'h10408000;
      13742: inst = 32'hc404faa;
      13743: inst = 32'h8220000;
      13744: inst = 32'h10408000;
      13745: inst = 32'hc404fb4;
      13746: inst = 32'h8220000;
      13747: inst = 32'h10408000;
      13748: inst = 32'hc405000;
      13749: inst = 32'h8220000;
      13750: inst = 32'h10408000;
      13751: inst = 32'hc40500a;
      13752: inst = 32'h8220000;
      13753: inst = 32'h10408000;
      13754: inst = 32'hc405014;
      13755: inst = 32'h8220000;
      13756: inst = 32'h10408000;
      13757: inst = 32'hc405060;
      13758: inst = 32'h8220000;
      13759: inst = 32'h10408000;
      13760: inst = 32'hc40506a;
      13761: inst = 32'h8220000;
      13762: inst = 32'h10408000;
      13763: inst = 32'hc405074;
      13764: inst = 32'h8220000;
      13765: inst = 32'h10408000;
      13766: inst = 32'hc4050c0;
      13767: inst = 32'h8220000;
      13768: inst = 32'h10408000;
      13769: inst = 32'hc4050ca;
      13770: inst = 32'h8220000;
      13771: inst = 32'h10408000;
      13772: inst = 32'hc4050d4;
      13773: inst = 32'h8220000;
      13774: inst = 32'h10408000;
      13775: inst = 32'hc405120;
      13776: inst = 32'h8220000;
      13777: inst = 32'h10408000;
      13778: inst = 32'hc40512a;
      13779: inst = 32'h8220000;
      13780: inst = 32'h10408000;
      13781: inst = 32'hc405134;
      13782: inst = 32'h8220000;
      13783: inst = 32'h10408000;
      13784: inst = 32'hc405180;
      13785: inst = 32'h8220000;
      13786: inst = 32'h10408000;
      13787: inst = 32'hc40518a;
      13788: inst = 32'h8220000;
      13789: inst = 32'h10408000;
      13790: inst = 32'hc405194;
      13791: inst = 32'h8220000;
      13792: inst = 32'h10408000;
      13793: inst = 32'hc4051a8;
      13794: inst = 32'h8220000;
      13795: inst = 32'h10408000;
      13796: inst = 32'hc4051a9;
      13797: inst = 32'h8220000;
      13798: inst = 32'h10408000;
      13799: inst = 32'hc4051b7;
      13800: inst = 32'h8220000;
      13801: inst = 32'h10408000;
      13802: inst = 32'hc4051e0;
      13803: inst = 32'h8220000;
      13804: inst = 32'h10408000;
      13805: inst = 32'hc4051ea;
      13806: inst = 32'h8220000;
      13807: inst = 32'h10408000;
      13808: inst = 32'hc4051f4;
      13809: inst = 32'h8220000;
      13810: inst = 32'h10408000;
      13811: inst = 32'hc405208;
      13812: inst = 32'h8220000;
      13813: inst = 32'h10408000;
      13814: inst = 32'hc405217;
      13815: inst = 32'h8220000;
      13816: inst = 32'h10408000;
      13817: inst = 32'hc405240;
      13818: inst = 32'h8220000;
      13819: inst = 32'h10408000;
      13820: inst = 32'hc40524a;
      13821: inst = 32'h8220000;
      13822: inst = 32'h10408000;
      13823: inst = 32'hc405254;
      13824: inst = 32'h8220000;
      13825: inst = 32'h10408000;
      13826: inst = 32'hc40525e;
      13827: inst = 32'h8220000;
      13828: inst = 32'h10408000;
      13829: inst = 32'hc405268;
      13830: inst = 32'h8220000;
      13831: inst = 32'h10408000;
      13832: inst = 32'hc405277;
      13833: inst = 32'h8220000;
      13834: inst = 32'h10408000;
      13835: inst = 32'hc405281;
      13836: inst = 32'h8220000;
      13837: inst = 32'h10408000;
      13838: inst = 32'hc4052a0;
      13839: inst = 32'h8220000;
      13840: inst = 32'h10408000;
      13841: inst = 32'hc4052a1;
      13842: inst = 32'h8220000;
      13843: inst = 32'h10408000;
      13844: inst = 32'hc4052a2;
      13845: inst = 32'h8220000;
      13846: inst = 32'h10408000;
      13847: inst = 32'hc4052a3;
      13848: inst = 32'h8220000;
      13849: inst = 32'h10408000;
      13850: inst = 32'hc4052a4;
      13851: inst = 32'h8220000;
      13852: inst = 32'h10408000;
      13853: inst = 32'hc4052a5;
      13854: inst = 32'h8220000;
      13855: inst = 32'h10408000;
      13856: inst = 32'hc4052a6;
      13857: inst = 32'h8220000;
      13858: inst = 32'h10408000;
      13859: inst = 32'hc4052a7;
      13860: inst = 32'h8220000;
      13861: inst = 32'h10408000;
      13862: inst = 32'hc4052a8;
      13863: inst = 32'h8220000;
      13864: inst = 32'h10408000;
      13865: inst = 32'hc4052a9;
      13866: inst = 32'h8220000;
      13867: inst = 32'h10408000;
      13868: inst = 32'hc4052aa;
      13869: inst = 32'h8220000;
      13870: inst = 32'h10408000;
      13871: inst = 32'hc4052ab;
      13872: inst = 32'h8220000;
      13873: inst = 32'h10408000;
      13874: inst = 32'hc4052ac;
      13875: inst = 32'h8220000;
      13876: inst = 32'h10408000;
      13877: inst = 32'hc4052ad;
      13878: inst = 32'h8220000;
      13879: inst = 32'h10408000;
      13880: inst = 32'hc4052ae;
      13881: inst = 32'h8220000;
      13882: inst = 32'h10408000;
      13883: inst = 32'hc4052af;
      13884: inst = 32'h8220000;
      13885: inst = 32'h10408000;
      13886: inst = 32'hc4052b0;
      13887: inst = 32'h8220000;
      13888: inst = 32'h10408000;
      13889: inst = 32'hc4052b1;
      13890: inst = 32'h8220000;
      13891: inst = 32'h10408000;
      13892: inst = 32'hc4052b2;
      13893: inst = 32'h8220000;
      13894: inst = 32'h10408000;
      13895: inst = 32'hc4052b3;
      13896: inst = 32'h8220000;
      13897: inst = 32'h10408000;
      13898: inst = 32'hc4052b4;
      13899: inst = 32'h8220000;
      13900: inst = 32'h10408000;
      13901: inst = 32'hc4052bd;
      13902: inst = 32'h8220000;
      13903: inst = 32'h10408000;
      13904: inst = 32'hc4052be;
      13905: inst = 32'h8220000;
      13906: inst = 32'h10408000;
      13907: inst = 32'hc4052c8;
      13908: inst = 32'h8220000;
      13909: inst = 32'h10408000;
      13910: inst = 32'hc4052d7;
      13911: inst = 32'h8220000;
      13912: inst = 32'h10408000;
      13913: inst = 32'hc4052e1;
      13914: inst = 32'h8220000;
      13915: inst = 32'h10408000;
      13916: inst = 32'hc4052e2;
      13917: inst = 32'h8220000;
      13918: inst = 32'h10408000;
      13919: inst = 32'hc40531c;
      13920: inst = 32'h8220000;
      13921: inst = 32'h10408000;
      13922: inst = 32'hc40531d;
      13923: inst = 32'h8220000;
      13924: inst = 32'h10408000;
      13925: inst = 32'hc40531e;
      13926: inst = 32'h8220000;
      13927: inst = 32'h10408000;
      13928: inst = 32'hc40531f;
      13929: inst = 32'h8220000;
      13930: inst = 32'h10408000;
      13931: inst = 32'hc405320;
      13932: inst = 32'h8220000;
      13933: inst = 32'h10408000;
      13934: inst = 32'hc405326;
      13935: inst = 32'h8220000;
      13936: inst = 32'h10408000;
      13937: inst = 32'hc405327;
      13938: inst = 32'h8220000;
      13939: inst = 32'h10408000;
      13940: inst = 32'hc405328;
      13941: inst = 32'h8220000;
      13942: inst = 32'h10408000;
      13943: inst = 32'hc405337;
      13944: inst = 32'h8220000;
      13945: inst = 32'h10408000;
      13946: inst = 32'hc405338;
      13947: inst = 32'h8220000;
      13948: inst = 32'h10408000;
      13949: inst = 32'hc405339;
      13950: inst = 32'h8220000;
      13951: inst = 32'h10408000;
      13952: inst = 32'hc40533f;
      13953: inst = 32'h8220000;
      13954: inst = 32'h10408000;
      13955: inst = 32'hc405340;
      13956: inst = 32'h8220000;
      13957: inst = 32'h10408000;
      13958: inst = 32'hc405341;
      13959: inst = 32'h8220000;
      13960: inst = 32'h10408000;
      13961: inst = 32'hc405342;
      13962: inst = 32'h8220000;
      13963: inst = 32'h10408000;
      13964: inst = 32'hc405343;
      13965: inst = 32'h8220000;
      13966: inst = 32'h10408000;
      13967: inst = 32'hc40537b;
      13968: inst = 32'h8220000;
      13969: inst = 32'h10408000;
      13970: inst = 32'hc40537c;
      13971: inst = 32'h8220000;
      13972: inst = 32'h10408000;
      13973: inst = 32'hc405386;
      13974: inst = 32'h8220000;
      13975: inst = 32'h10408000;
      13976: inst = 32'hc405387;
      13977: inst = 32'h8220000;
      13978: inst = 32'h10408000;
      13979: inst = 32'hc405388;
      13980: inst = 32'h8220000;
      13981: inst = 32'h10408000;
      13982: inst = 32'hc405397;
      13983: inst = 32'h8220000;
      13984: inst = 32'h10408000;
      13985: inst = 32'hc405398;
      13986: inst = 32'h8220000;
      13987: inst = 32'h10408000;
      13988: inst = 32'hc405399;
      13989: inst = 32'h8220000;
      13990: inst = 32'h10408000;
      13991: inst = 32'hc4053a3;
      13992: inst = 32'h8220000;
      13993: inst = 32'h10408000;
      13994: inst = 32'hc4053a4;
      13995: inst = 32'h8220000;
      13996: inst = 32'h10408000;
      13997: inst = 32'hc4053db;
      13998: inst = 32'h8220000;
      13999: inst = 32'h10408000;
      14000: inst = 32'hc4053e5;
      14001: inst = 32'h8220000;
      14002: inst = 32'h10408000;
      14003: inst = 32'hc4053e6;
      14004: inst = 32'h8220000;
      14005: inst = 32'h10408000;
      14006: inst = 32'hc4053e7;
      14007: inst = 32'h8220000;
      14008: inst = 32'h10408000;
      14009: inst = 32'hc4053f8;
      14010: inst = 32'h8220000;
      14011: inst = 32'h10408000;
      14012: inst = 32'hc4053f9;
      14013: inst = 32'h8220000;
      14014: inst = 32'h10408000;
      14015: inst = 32'hc4053fa;
      14016: inst = 32'h8220000;
      14017: inst = 32'h10408000;
      14018: inst = 32'hc405404;
      14019: inst = 32'h8220000;
      14020: inst = 32'h10408000;
      14021: inst = 32'hc40543a;
      14022: inst = 32'h8220000;
      14023: inst = 32'h10408000;
      14024: inst = 32'hc40543b;
      14025: inst = 32'h8220000;
      14026: inst = 32'h10408000;
      14027: inst = 32'hc405445;
      14028: inst = 32'h8220000;
      14029: inst = 32'h10408000;
      14030: inst = 32'hc405446;
      14031: inst = 32'h8220000;
      14032: inst = 32'h10408000;
      14033: inst = 32'hc405447;
      14034: inst = 32'h8220000;
      14035: inst = 32'h10408000;
      14036: inst = 32'hc405458;
      14037: inst = 32'h8220000;
      14038: inst = 32'h10408000;
      14039: inst = 32'hc405459;
      14040: inst = 32'h8220000;
      14041: inst = 32'h10408000;
      14042: inst = 32'hc40545a;
      14043: inst = 32'h8220000;
      14044: inst = 32'h10408000;
      14045: inst = 32'hc405464;
      14046: inst = 32'h8220000;
      14047: inst = 32'h10408000;
      14048: inst = 32'hc405465;
      14049: inst = 32'h8220000;
      14050: inst = 32'h10408000;
      14051: inst = 32'hc405499;
      14052: inst = 32'h8220000;
      14053: inst = 32'h10408000;
      14054: inst = 32'hc40549a;
      14055: inst = 32'h8220000;
      14056: inst = 32'h10408000;
      14057: inst = 32'hc4054a5;
      14058: inst = 32'h8220000;
      14059: inst = 32'h10408000;
      14060: inst = 32'hc4054a6;
      14061: inst = 32'h8220000;
      14062: inst = 32'h10408000;
      14063: inst = 32'hc4054a7;
      14064: inst = 32'h8220000;
      14065: inst = 32'h10408000;
      14066: inst = 32'hc4054b8;
      14067: inst = 32'h8220000;
      14068: inst = 32'h10408000;
      14069: inst = 32'hc4054b9;
      14070: inst = 32'h8220000;
      14071: inst = 32'h10408000;
      14072: inst = 32'hc4054ba;
      14073: inst = 32'h8220000;
      14074: inst = 32'h10408000;
      14075: inst = 32'hc4054c5;
      14076: inst = 32'h8220000;
      14077: inst = 32'h10408000;
      14078: inst = 32'hc4054c6;
      14079: inst = 32'h8220000;
      14080: inst = 32'h10408000;
      14081: inst = 32'hc4054f8;
      14082: inst = 32'h8220000;
      14083: inst = 32'h10408000;
      14084: inst = 32'hc4054f9;
      14085: inst = 32'h8220000;
      14086: inst = 32'h10408000;
      14087: inst = 32'hc405500;
      14088: inst = 32'h8220000;
      14089: inst = 32'h10408000;
      14090: inst = 32'hc405504;
      14091: inst = 32'h8220000;
      14092: inst = 32'h10408000;
      14093: inst = 32'hc405505;
      14094: inst = 32'h8220000;
      14095: inst = 32'h10408000;
      14096: inst = 32'hc405506;
      14097: inst = 32'h8220000;
      14098: inst = 32'h10408000;
      14099: inst = 32'hc405507;
      14100: inst = 32'h8220000;
      14101: inst = 32'h10408000;
      14102: inst = 32'hc405518;
      14103: inst = 32'h8220000;
      14104: inst = 32'h10408000;
      14105: inst = 32'hc405519;
      14106: inst = 32'h8220000;
      14107: inst = 32'h10408000;
      14108: inst = 32'hc40551a;
      14109: inst = 32'h8220000;
      14110: inst = 32'h10408000;
      14111: inst = 32'hc40551b;
      14112: inst = 32'h8220000;
      14113: inst = 32'h10408000;
      14114: inst = 32'hc40551f;
      14115: inst = 32'h8220000;
      14116: inst = 32'h10408000;
      14117: inst = 32'hc405526;
      14118: inst = 32'h8220000;
      14119: inst = 32'h10408000;
      14120: inst = 32'hc405527;
      14121: inst = 32'h8220000;
      14122: inst = 32'h10408000;
      14123: inst = 32'hc405558;
      14124: inst = 32'h8220000;
      14125: inst = 32'h10408000;
      14126: inst = 32'hc405559;
      14127: inst = 32'h8220000;
      14128: inst = 32'h10408000;
      14129: inst = 32'hc405560;
      14130: inst = 32'h8220000;
      14131: inst = 32'h10408000;
      14132: inst = 32'hc405564;
      14133: inst = 32'h8220000;
      14134: inst = 32'h10408000;
      14135: inst = 32'hc405565;
      14136: inst = 32'h8220000;
      14137: inst = 32'h10408000;
      14138: inst = 32'hc405566;
      14139: inst = 32'h8220000;
      14140: inst = 32'h10408000;
      14141: inst = 32'hc405567;
      14142: inst = 32'h8220000;
      14143: inst = 32'h10408000;
      14144: inst = 32'hc405578;
      14145: inst = 32'h8220000;
      14146: inst = 32'h10408000;
      14147: inst = 32'hc405579;
      14148: inst = 32'h8220000;
      14149: inst = 32'h10408000;
      14150: inst = 32'hc40557a;
      14151: inst = 32'h8220000;
      14152: inst = 32'h10408000;
      14153: inst = 32'hc40557b;
      14154: inst = 32'h8220000;
      14155: inst = 32'h10408000;
      14156: inst = 32'hc40557f;
      14157: inst = 32'h8220000;
      14158: inst = 32'h10408000;
      14159: inst = 32'hc405586;
      14160: inst = 32'h8220000;
      14161: inst = 32'h10408000;
      14162: inst = 32'hc405587;
      14163: inst = 32'h8220000;
      14164: inst = 32'h10408000;
      14165: inst = 32'hc4055b7;
      14166: inst = 32'h8220000;
      14167: inst = 32'h10408000;
      14168: inst = 32'hc4055b8;
      14169: inst = 32'h8220000;
      14170: inst = 32'h10408000;
      14171: inst = 32'hc4055bf;
      14172: inst = 32'h8220000;
      14173: inst = 32'h10408000;
      14174: inst = 32'hc4055c0;
      14175: inst = 32'h8220000;
      14176: inst = 32'h10408000;
      14177: inst = 32'hc4055c4;
      14178: inst = 32'h8220000;
      14179: inst = 32'h10408000;
      14180: inst = 32'hc4055c5;
      14181: inst = 32'h8220000;
      14182: inst = 32'h10408000;
      14183: inst = 32'hc4055c6;
      14184: inst = 32'h8220000;
      14185: inst = 32'h10408000;
      14186: inst = 32'hc4055c7;
      14187: inst = 32'h8220000;
      14188: inst = 32'h10408000;
      14189: inst = 32'hc4055d8;
      14190: inst = 32'h8220000;
      14191: inst = 32'h10408000;
      14192: inst = 32'hc4055d9;
      14193: inst = 32'h8220000;
      14194: inst = 32'h10408000;
      14195: inst = 32'hc4055da;
      14196: inst = 32'h8220000;
      14197: inst = 32'h10408000;
      14198: inst = 32'hc4055db;
      14199: inst = 32'h8220000;
      14200: inst = 32'h10408000;
      14201: inst = 32'hc4055df;
      14202: inst = 32'h8220000;
      14203: inst = 32'h10408000;
      14204: inst = 32'hc4055e0;
      14205: inst = 32'h8220000;
      14206: inst = 32'h10408000;
      14207: inst = 32'hc4055e7;
      14208: inst = 32'h8220000;
      14209: inst = 32'h10408000;
      14210: inst = 32'hc4055e8;
      14211: inst = 32'h8220000;
      14212: inst = 32'h10408000;
      14213: inst = 32'hc405616;
      14214: inst = 32'h8220000;
      14215: inst = 32'h10408000;
      14216: inst = 32'hc405617;
      14217: inst = 32'h8220000;
      14218: inst = 32'h10408000;
      14219: inst = 32'hc40561f;
      14220: inst = 32'h8220000;
      14221: inst = 32'h10408000;
      14222: inst = 32'hc405620;
      14223: inst = 32'h8220000;
      14224: inst = 32'h10408000;
      14225: inst = 32'hc405623;
      14226: inst = 32'h8220000;
      14227: inst = 32'h10408000;
      14228: inst = 32'hc405624;
      14229: inst = 32'h8220000;
      14230: inst = 32'h10408000;
      14231: inst = 32'hc405625;
      14232: inst = 32'h8220000;
      14233: inst = 32'h10408000;
      14234: inst = 32'hc405626;
      14235: inst = 32'h8220000;
      14236: inst = 32'h10408000;
      14237: inst = 32'hc405639;
      14238: inst = 32'h8220000;
      14239: inst = 32'h10408000;
      14240: inst = 32'hc40563a;
      14241: inst = 32'h8220000;
      14242: inst = 32'h10408000;
      14243: inst = 32'hc40563b;
      14244: inst = 32'h8220000;
      14245: inst = 32'h10408000;
      14246: inst = 32'hc40563c;
      14247: inst = 32'h8220000;
      14248: inst = 32'h10408000;
      14249: inst = 32'hc40563f;
      14250: inst = 32'h8220000;
      14251: inst = 32'h10408000;
      14252: inst = 32'hc405640;
      14253: inst = 32'h8220000;
      14254: inst = 32'h10408000;
      14255: inst = 32'hc405648;
      14256: inst = 32'h8220000;
      14257: inst = 32'h10408000;
      14258: inst = 32'hc405649;
      14259: inst = 32'h8220000;
      14260: inst = 32'h10408000;
      14261: inst = 32'hc405675;
      14262: inst = 32'h8220000;
      14263: inst = 32'h10408000;
      14264: inst = 32'hc405676;
      14265: inst = 32'h8220000;
      14266: inst = 32'h10408000;
      14267: inst = 32'hc405677;
      14268: inst = 32'h8220000;
      14269: inst = 32'h10408000;
      14270: inst = 32'hc40567e;
      14271: inst = 32'h8220000;
      14272: inst = 32'h10408000;
      14273: inst = 32'hc40567f;
      14274: inst = 32'h8220000;
      14275: inst = 32'h10408000;
      14276: inst = 32'hc405680;
      14277: inst = 32'h8220000;
      14278: inst = 32'h10408000;
      14279: inst = 32'hc405683;
      14280: inst = 32'h8220000;
      14281: inst = 32'h10408000;
      14282: inst = 32'hc405684;
      14283: inst = 32'h8220000;
      14284: inst = 32'h10408000;
      14285: inst = 32'hc405685;
      14286: inst = 32'h8220000;
      14287: inst = 32'h10408000;
      14288: inst = 32'hc405686;
      14289: inst = 32'h8220000;
      14290: inst = 32'h10408000;
      14291: inst = 32'hc405699;
      14292: inst = 32'h8220000;
      14293: inst = 32'h10408000;
      14294: inst = 32'hc40569a;
      14295: inst = 32'h8220000;
      14296: inst = 32'h10408000;
      14297: inst = 32'hc40569b;
      14298: inst = 32'h8220000;
      14299: inst = 32'h10408000;
      14300: inst = 32'hc40569c;
      14301: inst = 32'h8220000;
      14302: inst = 32'h10408000;
      14303: inst = 32'hc40569f;
      14304: inst = 32'h8220000;
      14305: inst = 32'h10408000;
      14306: inst = 32'hc4056a0;
      14307: inst = 32'h8220000;
      14308: inst = 32'h10408000;
      14309: inst = 32'hc4056a1;
      14310: inst = 32'h8220000;
      14311: inst = 32'h10408000;
      14312: inst = 32'hc4056a8;
      14313: inst = 32'h8220000;
      14314: inst = 32'h10408000;
      14315: inst = 32'hc4056a9;
      14316: inst = 32'h8220000;
      14317: inst = 32'h10408000;
      14318: inst = 32'hc4056aa;
      14319: inst = 32'h8220000;
      14320: inst = 32'h10408000;
      14321: inst = 32'hc4056d4;
      14322: inst = 32'h8220000;
      14323: inst = 32'h10408000;
      14324: inst = 32'hc4056d5;
      14325: inst = 32'h8220000;
      14326: inst = 32'h10408000;
      14327: inst = 32'hc4056d6;
      14328: inst = 32'h8220000;
      14329: inst = 32'h10408000;
      14330: inst = 32'hc4056d7;
      14331: inst = 32'h8220000;
      14332: inst = 32'h10408000;
      14333: inst = 32'hc4056d8;
      14334: inst = 32'h8220000;
      14335: inst = 32'h10408000;
      14336: inst = 32'hc4056d9;
      14337: inst = 32'h8220000;
      14338: inst = 32'h10408000;
      14339: inst = 32'hc4056da;
      14340: inst = 32'h8220000;
      14341: inst = 32'h10408000;
      14342: inst = 32'hc4056db;
      14343: inst = 32'h8220000;
      14344: inst = 32'h10408000;
      14345: inst = 32'hc4056dc;
      14346: inst = 32'h8220000;
      14347: inst = 32'h10408000;
      14348: inst = 32'hc4056dd;
      14349: inst = 32'h8220000;
      14350: inst = 32'h10408000;
      14351: inst = 32'hc4056de;
      14352: inst = 32'h8220000;
      14353: inst = 32'h10408000;
      14354: inst = 32'hc4056df;
      14355: inst = 32'h8220000;
      14356: inst = 32'h10408000;
      14357: inst = 32'hc4056e0;
      14358: inst = 32'h8220000;
      14359: inst = 32'h10408000;
      14360: inst = 32'hc4056e3;
      14361: inst = 32'h8220000;
      14362: inst = 32'h10408000;
      14363: inst = 32'hc4056e4;
      14364: inst = 32'h8220000;
      14365: inst = 32'h10408000;
      14366: inst = 32'hc4056e5;
      14367: inst = 32'h8220000;
      14368: inst = 32'h10408000;
      14369: inst = 32'hc4056e6;
      14370: inst = 32'h8220000;
      14371: inst = 32'h10408000;
      14372: inst = 32'hc4056f9;
      14373: inst = 32'h8220000;
      14374: inst = 32'h10408000;
      14375: inst = 32'hc4056fa;
      14376: inst = 32'h8220000;
      14377: inst = 32'h10408000;
      14378: inst = 32'hc4056fb;
      14379: inst = 32'h8220000;
      14380: inst = 32'h10408000;
      14381: inst = 32'hc4056fc;
      14382: inst = 32'h8220000;
      14383: inst = 32'h10408000;
      14384: inst = 32'hc4056ff;
      14385: inst = 32'h8220000;
      14386: inst = 32'h10408000;
      14387: inst = 32'hc405700;
      14388: inst = 32'h8220000;
      14389: inst = 32'h10408000;
      14390: inst = 32'hc405701;
      14391: inst = 32'h8220000;
      14392: inst = 32'h10408000;
      14393: inst = 32'hc405702;
      14394: inst = 32'h8220000;
      14395: inst = 32'h10408000;
      14396: inst = 32'hc405703;
      14397: inst = 32'h8220000;
      14398: inst = 32'h10408000;
      14399: inst = 32'hc405704;
      14400: inst = 32'h8220000;
      14401: inst = 32'h10408000;
      14402: inst = 32'hc405705;
      14403: inst = 32'h8220000;
      14404: inst = 32'h10408000;
      14405: inst = 32'hc405706;
      14406: inst = 32'h8220000;
      14407: inst = 32'h10408000;
      14408: inst = 32'hc405707;
      14409: inst = 32'h8220000;
      14410: inst = 32'h10408000;
      14411: inst = 32'hc405708;
      14412: inst = 32'h8220000;
      14413: inst = 32'h10408000;
      14414: inst = 32'hc405709;
      14415: inst = 32'h8220000;
      14416: inst = 32'h10408000;
      14417: inst = 32'hc40570a;
      14418: inst = 32'h8220000;
      14419: inst = 32'h10408000;
      14420: inst = 32'hc405734;
      14421: inst = 32'h8220000;
      14422: inst = 32'h10408000;
      14423: inst = 32'hc405735;
      14424: inst = 32'h8220000;
      14425: inst = 32'h10408000;
      14426: inst = 32'hc405736;
      14427: inst = 32'h8220000;
      14428: inst = 32'h10408000;
      14429: inst = 32'hc405737;
      14430: inst = 32'h8220000;
      14431: inst = 32'h10408000;
      14432: inst = 32'hc405738;
      14433: inst = 32'h8220000;
      14434: inst = 32'h10408000;
      14435: inst = 32'hc405739;
      14436: inst = 32'h8220000;
      14437: inst = 32'h10408000;
      14438: inst = 32'hc40573a;
      14439: inst = 32'h8220000;
      14440: inst = 32'h10408000;
      14441: inst = 32'hc40573b;
      14442: inst = 32'h8220000;
      14443: inst = 32'h10408000;
      14444: inst = 32'hc40573c;
      14445: inst = 32'h8220000;
      14446: inst = 32'h10408000;
      14447: inst = 32'hc40573d;
      14448: inst = 32'h8220000;
      14449: inst = 32'h10408000;
      14450: inst = 32'hc40573e;
      14451: inst = 32'h8220000;
      14452: inst = 32'h10408000;
      14453: inst = 32'hc40573f;
      14454: inst = 32'h8220000;
      14455: inst = 32'h10408000;
      14456: inst = 32'hc405740;
      14457: inst = 32'h8220000;
      14458: inst = 32'h10408000;
      14459: inst = 32'hc405742;
      14460: inst = 32'h8220000;
      14461: inst = 32'h10408000;
      14462: inst = 32'hc405743;
      14463: inst = 32'h8220000;
      14464: inst = 32'h10408000;
      14465: inst = 32'hc405744;
      14466: inst = 32'h8220000;
      14467: inst = 32'h10408000;
      14468: inst = 32'hc405745;
      14469: inst = 32'h8220000;
      14470: inst = 32'h10408000;
      14471: inst = 32'hc405746;
      14472: inst = 32'h8220000;
      14473: inst = 32'h10408000;
      14474: inst = 32'hc405759;
      14475: inst = 32'h8220000;
      14476: inst = 32'h10408000;
      14477: inst = 32'hc40575a;
      14478: inst = 32'h8220000;
      14479: inst = 32'h10408000;
      14480: inst = 32'hc40575b;
      14481: inst = 32'h8220000;
      14482: inst = 32'h10408000;
      14483: inst = 32'hc40575c;
      14484: inst = 32'h8220000;
      14485: inst = 32'h10408000;
      14486: inst = 32'hc40575d;
      14487: inst = 32'h8220000;
      14488: inst = 32'h10408000;
      14489: inst = 32'hc40575f;
      14490: inst = 32'h8220000;
      14491: inst = 32'h10408000;
      14492: inst = 32'hc405760;
      14493: inst = 32'h8220000;
      14494: inst = 32'h10408000;
      14495: inst = 32'hc405761;
      14496: inst = 32'h8220000;
      14497: inst = 32'h10408000;
      14498: inst = 32'hc405762;
      14499: inst = 32'h8220000;
      14500: inst = 32'h10408000;
      14501: inst = 32'hc405763;
      14502: inst = 32'h8220000;
      14503: inst = 32'h10408000;
      14504: inst = 32'hc405764;
      14505: inst = 32'h8220000;
      14506: inst = 32'h10408000;
      14507: inst = 32'hc405765;
      14508: inst = 32'h8220000;
      14509: inst = 32'h10408000;
      14510: inst = 32'hc405766;
      14511: inst = 32'h8220000;
      14512: inst = 32'h10408000;
      14513: inst = 32'hc405767;
      14514: inst = 32'h8220000;
      14515: inst = 32'h10408000;
      14516: inst = 32'hc405768;
      14517: inst = 32'h8220000;
      14518: inst = 32'h10408000;
      14519: inst = 32'hc405769;
      14520: inst = 32'h8220000;
      14521: inst = 32'h10408000;
      14522: inst = 32'hc40576a;
      14523: inst = 32'h8220000;
      14524: inst = 32'h10408000;
      14525: inst = 32'hc40576b;
      14526: inst = 32'h8220000;
      14527: inst = 32'h10408000;
      14528: inst = 32'hc405793;
      14529: inst = 32'h8220000;
      14530: inst = 32'h10408000;
      14531: inst = 32'hc405794;
      14532: inst = 32'h8220000;
      14533: inst = 32'h10408000;
      14534: inst = 32'hc405795;
      14535: inst = 32'h8220000;
      14536: inst = 32'h10408000;
      14537: inst = 32'hc405796;
      14538: inst = 32'h8220000;
      14539: inst = 32'h10408000;
      14540: inst = 32'hc405797;
      14541: inst = 32'h8220000;
      14542: inst = 32'h10408000;
      14543: inst = 32'hc405798;
      14544: inst = 32'h8220000;
      14545: inst = 32'h10408000;
      14546: inst = 32'hc405799;
      14547: inst = 32'h8220000;
      14548: inst = 32'h10408000;
      14549: inst = 32'hc40579a;
      14550: inst = 32'h8220000;
      14551: inst = 32'h10408000;
      14552: inst = 32'hc40579b;
      14553: inst = 32'h8220000;
      14554: inst = 32'h10408000;
      14555: inst = 32'hc40579c;
      14556: inst = 32'h8220000;
      14557: inst = 32'h10408000;
      14558: inst = 32'hc40579d;
      14559: inst = 32'h8220000;
      14560: inst = 32'h10408000;
      14561: inst = 32'hc40579e;
      14562: inst = 32'h8220000;
      14563: inst = 32'h10408000;
      14564: inst = 32'hc40579f;
      14565: inst = 32'h8220000;
      14566: inst = 32'h10408000;
      14567: inst = 32'hc4057a0;
      14568: inst = 32'h8220000;
      14569: inst = 32'h10408000;
      14570: inst = 32'hc4057a1;
      14571: inst = 32'h8220000;
      14572: inst = 32'h10408000;
      14573: inst = 32'hc4057a2;
      14574: inst = 32'h8220000;
      14575: inst = 32'h10408000;
      14576: inst = 32'hc4057a3;
      14577: inst = 32'h8220000;
      14578: inst = 32'h10408000;
      14579: inst = 32'hc4057a4;
      14580: inst = 32'h8220000;
      14581: inst = 32'h10408000;
      14582: inst = 32'hc4057a5;
      14583: inst = 32'h8220000;
      14584: inst = 32'h10408000;
      14585: inst = 32'hc4057a6;
      14586: inst = 32'h8220000;
      14587: inst = 32'h10408000;
      14588: inst = 32'hc4057b9;
      14589: inst = 32'h8220000;
      14590: inst = 32'h10408000;
      14591: inst = 32'hc4057ba;
      14592: inst = 32'h8220000;
      14593: inst = 32'h10408000;
      14594: inst = 32'hc4057bb;
      14595: inst = 32'h8220000;
      14596: inst = 32'h10408000;
      14597: inst = 32'hc4057bc;
      14598: inst = 32'h8220000;
      14599: inst = 32'h10408000;
      14600: inst = 32'hc4057bd;
      14601: inst = 32'h8220000;
      14602: inst = 32'h10408000;
      14603: inst = 32'hc4057be;
      14604: inst = 32'h8220000;
      14605: inst = 32'h10408000;
      14606: inst = 32'hc4057bf;
      14607: inst = 32'h8220000;
      14608: inst = 32'h10408000;
      14609: inst = 32'hc4057c0;
      14610: inst = 32'h8220000;
      14611: inst = 32'h10408000;
      14612: inst = 32'hc4057c1;
      14613: inst = 32'h8220000;
      14614: inst = 32'h10408000;
      14615: inst = 32'hc4057c2;
      14616: inst = 32'h8220000;
      14617: inst = 32'h10408000;
      14618: inst = 32'hc4057c3;
      14619: inst = 32'h8220000;
      14620: inst = 32'h10408000;
      14621: inst = 32'hc4057c4;
      14622: inst = 32'h8220000;
      14623: inst = 32'h10408000;
      14624: inst = 32'hc4057c5;
      14625: inst = 32'h8220000;
      14626: inst = 32'h10408000;
      14627: inst = 32'hc4057c6;
      14628: inst = 32'h8220000;
      14629: inst = 32'h10408000;
      14630: inst = 32'hc4057c7;
      14631: inst = 32'h8220000;
      14632: inst = 32'h10408000;
      14633: inst = 32'hc4057c8;
      14634: inst = 32'h8220000;
      14635: inst = 32'h10408000;
      14636: inst = 32'hc4057c9;
      14637: inst = 32'h8220000;
      14638: inst = 32'h10408000;
      14639: inst = 32'hc4057ca;
      14640: inst = 32'h8220000;
      14641: inst = 32'h10408000;
      14642: inst = 32'hc4057cb;
      14643: inst = 32'h8220000;
      14644: inst = 32'h10408000;
      14645: inst = 32'hc4057cc;
      14646: inst = 32'h8220000;
      14647: inst = 32'hc20bdd7;
      14648: inst = 32'h10408000;
      14649: inst = 32'hc404dc1;
      14650: inst = 32'h8220000;
      14651: inst = 32'h10408000;
      14652: inst = 32'hc404dc2;
      14653: inst = 32'h8220000;
      14654: inst = 32'h10408000;
      14655: inst = 32'hc404dc3;
      14656: inst = 32'h8220000;
      14657: inst = 32'h10408000;
      14658: inst = 32'hc404dc4;
      14659: inst = 32'h8220000;
      14660: inst = 32'h10408000;
      14661: inst = 32'hc404dc5;
      14662: inst = 32'h8220000;
      14663: inst = 32'h10408000;
      14664: inst = 32'hc404dc6;
      14665: inst = 32'h8220000;
      14666: inst = 32'h10408000;
      14667: inst = 32'hc404dc7;
      14668: inst = 32'h8220000;
      14669: inst = 32'h10408000;
      14670: inst = 32'hc404dc8;
      14671: inst = 32'h8220000;
      14672: inst = 32'h10408000;
      14673: inst = 32'hc404dc9;
      14674: inst = 32'h8220000;
      14675: inst = 32'h10408000;
      14676: inst = 32'hc404dcb;
      14677: inst = 32'h8220000;
      14678: inst = 32'h10408000;
      14679: inst = 32'hc404dcc;
      14680: inst = 32'h8220000;
      14681: inst = 32'h10408000;
      14682: inst = 32'hc404dcd;
      14683: inst = 32'h8220000;
      14684: inst = 32'h10408000;
      14685: inst = 32'hc404dce;
      14686: inst = 32'h8220000;
      14687: inst = 32'h10408000;
      14688: inst = 32'hc404dcf;
      14689: inst = 32'h8220000;
      14690: inst = 32'h10408000;
      14691: inst = 32'hc404dd0;
      14692: inst = 32'h8220000;
      14693: inst = 32'h10408000;
      14694: inst = 32'hc404dd1;
      14695: inst = 32'h8220000;
      14696: inst = 32'h10408000;
      14697: inst = 32'hc404dd2;
      14698: inst = 32'h8220000;
      14699: inst = 32'h10408000;
      14700: inst = 32'hc404dd3;
      14701: inst = 32'h8220000;
      14702: inst = 32'h10408000;
      14703: inst = 32'hc404e21;
      14704: inst = 32'h8220000;
      14705: inst = 32'h10408000;
      14706: inst = 32'hc404e22;
      14707: inst = 32'h8220000;
      14708: inst = 32'h10408000;
      14709: inst = 32'hc404e23;
      14710: inst = 32'h8220000;
      14711: inst = 32'h10408000;
      14712: inst = 32'hc404e24;
      14713: inst = 32'h8220000;
      14714: inst = 32'h10408000;
      14715: inst = 32'hc404e25;
      14716: inst = 32'h8220000;
      14717: inst = 32'h10408000;
      14718: inst = 32'hc404e26;
      14719: inst = 32'h8220000;
      14720: inst = 32'h10408000;
      14721: inst = 32'hc404e27;
      14722: inst = 32'h8220000;
      14723: inst = 32'h10408000;
      14724: inst = 32'hc404e28;
      14725: inst = 32'h8220000;
      14726: inst = 32'h10408000;
      14727: inst = 32'hc404e29;
      14728: inst = 32'h8220000;
      14729: inst = 32'h10408000;
      14730: inst = 32'hc404e2b;
      14731: inst = 32'h8220000;
      14732: inst = 32'h10408000;
      14733: inst = 32'hc404e2c;
      14734: inst = 32'h8220000;
      14735: inst = 32'h10408000;
      14736: inst = 32'hc404e2d;
      14737: inst = 32'h8220000;
      14738: inst = 32'h10408000;
      14739: inst = 32'hc404e2e;
      14740: inst = 32'h8220000;
      14741: inst = 32'h10408000;
      14742: inst = 32'hc404e2f;
      14743: inst = 32'h8220000;
      14744: inst = 32'h10408000;
      14745: inst = 32'hc404e30;
      14746: inst = 32'h8220000;
      14747: inst = 32'h10408000;
      14748: inst = 32'hc404e31;
      14749: inst = 32'h8220000;
      14750: inst = 32'h10408000;
      14751: inst = 32'hc404e32;
      14752: inst = 32'h8220000;
      14753: inst = 32'h10408000;
      14754: inst = 32'hc404e33;
      14755: inst = 32'h8220000;
      14756: inst = 32'h10408000;
      14757: inst = 32'hc404e81;
      14758: inst = 32'h8220000;
      14759: inst = 32'h10408000;
      14760: inst = 32'hc404e82;
      14761: inst = 32'h8220000;
      14762: inst = 32'h10408000;
      14763: inst = 32'hc404e83;
      14764: inst = 32'h8220000;
      14765: inst = 32'h10408000;
      14766: inst = 32'hc404e84;
      14767: inst = 32'h8220000;
      14768: inst = 32'h10408000;
      14769: inst = 32'hc404e85;
      14770: inst = 32'h8220000;
      14771: inst = 32'h10408000;
      14772: inst = 32'hc404e86;
      14773: inst = 32'h8220000;
      14774: inst = 32'h10408000;
      14775: inst = 32'hc404e87;
      14776: inst = 32'h8220000;
      14777: inst = 32'h10408000;
      14778: inst = 32'hc404e88;
      14779: inst = 32'h8220000;
      14780: inst = 32'h10408000;
      14781: inst = 32'hc404e89;
      14782: inst = 32'h8220000;
      14783: inst = 32'h10408000;
      14784: inst = 32'hc404e8b;
      14785: inst = 32'h8220000;
      14786: inst = 32'h10408000;
      14787: inst = 32'hc404e8c;
      14788: inst = 32'h8220000;
      14789: inst = 32'h10408000;
      14790: inst = 32'hc404e8d;
      14791: inst = 32'h8220000;
      14792: inst = 32'h10408000;
      14793: inst = 32'hc404e8e;
      14794: inst = 32'h8220000;
      14795: inst = 32'h10408000;
      14796: inst = 32'hc404e8f;
      14797: inst = 32'h8220000;
      14798: inst = 32'h10408000;
      14799: inst = 32'hc404e90;
      14800: inst = 32'h8220000;
      14801: inst = 32'h10408000;
      14802: inst = 32'hc404e91;
      14803: inst = 32'h8220000;
      14804: inst = 32'h10408000;
      14805: inst = 32'hc404e92;
      14806: inst = 32'h8220000;
      14807: inst = 32'h10408000;
      14808: inst = 32'hc404e93;
      14809: inst = 32'h8220000;
      14810: inst = 32'h10408000;
      14811: inst = 32'hc404ee1;
      14812: inst = 32'h8220000;
      14813: inst = 32'h10408000;
      14814: inst = 32'hc404ee2;
      14815: inst = 32'h8220000;
      14816: inst = 32'h10408000;
      14817: inst = 32'hc404ee3;
      14818: inst = 32'h8220000;
      14819: inst = 32'h10408000;
      14820: inst = 32'hc404ee4;
      14821: inst = 32'h8220000;
      14822: inst = 32'h10408000;
      14823: inst = 32'hc404ee5;
      14824: inst = 32'h8220000;
      14825: inst = 32'h10408000;
      14826: inst = 32'hc404ee6;
      14827: inst = 32'h8220000;
      14828: inst = 32'h10408000;
      14829: inst = 32'hc404ee7;
      14830: inst = 32'h8220000;
      14831: inst = 32'h10408000;
      14832: inst = 32'hc404ee8;
      14833: inst = 32'h8220000;
      14834: inst = 32'h10408000;
      14835: inst = 32'hc404ee9;
      14836: inst = 32'h8220000;
      14837: inst = 32'h10408000;
      14838: inst = 32'hc404eeb;
      14839: inst = 32'h8220000;
      14840: inst = 32'h10408000;
      14841: inst = 32'hc404eec;
      14842: inst = 32'h8220000;
      14843: inst = 32'h10408000;
      14844: inst = 32'hc404eed;
      14845: inst = 32'h8220000;
      14846: inst = 32'h10408000;
      14847: inst = 32'hc404eee;
      14848: inst = 32'h8220000;
      14849: inst = 32'h10408000;
      14850: inst = 32'hc404eef;
      14851: inst = 32'h8220000;
      14852: inst = 32'h10408000;
      14853: inst = 32'hc404ef0;
      14854: inst = 32'h8220000;
      14855: inst = 32'h10408000;
      14856: inst = 32'hc404ef1;
      14857: inst = 32'h8220000;
      14858: inst = 32'h10408000;
      14859: inst = 32'hc404ef2;
      14860: inst = 32'h8220000;
      14861: inst = 32'h10408000;
      14862: inst = 32'hc404ef3;
      14863: inst = 32'h8220000;
      14864: inst = 32'h10408000;
      14865: inst = 32'hc404f41;
      14866: inst = 32'h8220000;
      14867: inst = 32'h10408000;
      14868: inst = 32'hc404f42;
      14869: inst = 32'h8220000;
      14870: inst = 32'h10408000;
      14871: inst = 32'hc404f43;
      14872: inst = 32'h8220000;
      14873: inst = 32'h10408000;
      14874: inst = 32'hc404f44;
      14875: inst = 32'h8220000;
      14876: inst = 32'h10408000;
      14877: inst = 32'hc404f45;
      14878: inst = 32'h8220000;
      14879: inst = 32'h10408000;
      14880: inst = 32'hc404f46;
      14881: inst = 32'h8220000;
      14882: inst = 32'h10408000;
      14883: inst = 32'hc404f47;
      14884: inst = 32'h8220000;
      14885: inst = 32'h10408000;
      14886: inst = 32'hc404f48;
      14887: inst = 32'h8220000;
      14888: inst = 32'h10408000;
      14889: inst = 32'hc404f49;
      14890: inst = 32'h8220000;
      14891: inst = 32'h10408000;
      14892: inst = 32'hc404f4b;
      14893: inst = 32'h8220000;
      14894: inst = 32'h10408000;
      14895: inst = 32'hc404f4c;
      14896: inst = 32'h8220000;
      14897: inst = 32'h10408000;
      14898: inst = 32'hc404f4d;
      14899: inst = 32'h8220000;
      14900: inst = 32'h10408000;
      14901: inst = 32'hc404f4e;
      14902: inst = 32'h8220000;
      14903: inst = 32'h10408000;
      14904: inst = 32'hc404f4f;
      14905: inst = 32'h8220000;
      14906: inst = 32'h10408000;
      14907: inst = 32'hc404f50;
      14908: inst = 32'h8220000;
      14909: inst = 32'h10408000;
      14910: inst = 32'hc404f51;
      14911: inst = 32'h8220000;
      14912: inst = 32'h10408000;
      14913: inst = 32'hc404f52;
      14914: inst = 32'h8220000;
      14915: inst = 32'h10408000;
      14916: inst = 32'hc404f53;
      14917: inst = 32'h8220000;
      14918: inst = 32'h10408000;
      14919: inst = 32'hc404fa1;
      14920: inst = 32'h8220000;
      14921: inst = 32'h10408000;
      14922: inst = 32'hc404fa2;
      14923: inst = 32'h8220000;
      14924: inst = 32'h10408000;
      14925: inst = 32'hc404fa3;
      14926: inst = 32'h8220000;
      14927: inst = 32'h10408000;
      14928: inst = 32'hc404fa4;
      14929: inst = 32'h8220000;
      14930: inst = 32'h10408000;
      14931: inst = 32'hc404fa5;
      14932: inst = 32'h8220000;
      14933: inst = 32'h10408000;
      14934: inst = 32'hc404fa6;
      14935: inst = 32'h8220000;
      14936: inst = 32'h10408000;
      14937: inst = 32'hc404fa7;
      14938: inst = 32'h8220000;
      14939: inst = 32'h10408000;
      14940: inst = 32'hc404fa9;
      14941: inst = 32'h8220000;
      14942: inst = 32'h10408000;
      14943: inst = 32'hc404fab;
      14944: inst = 32'h8220000;
      14945: inst = 32'h10408000;
      14946: inst = 32'hc404fad;
      14947: inst = 32'h8220000;
      14948: inst = 32'h10408000;
      14949: inst = 32'hc404fae;
      14950: inst = 32'h8220000;
      14951: inst = 32'h10408000;
      14952: inst = 32'hc404faf;
      14953: inst = 32'h8220000;
      14954: inst = 32'h10408000;
      14955: inst = 32'hc404fb0;
      14956: inst = 32'h8220000;
      14957: inst = 32'h10408000;
      14958: inst = 32'hc404fb1;
      14959: inst = 32'h8220000;
      14960: inst = 32'h10408000;
      14961: inst = 32'hc404fb2;
      14962: inst = 32'h8220000;
      14963: inst = 32'h10408000;
      14964: inst = 32'hc404fb3;
      14965: inst = 32'h8220000;
      14966: inst = 32'h10408000;
      14967: inst = 32'hc405001;
      14968: inst = 32'h8220000;
      14969: inst = 32'h10408000;
      14970: inst = 32'hc405002;
      14971: inst = 32'h8220000;
      14972: inst = 32'h10408000;
      14973: inst = 32'hc405003;
      14974: inst = 32'h8220000;
      14975: inst = 32'h10408000;
      14976: inst = 32'hc405004;
      14977: inst = 32'h8220000;
      14978: inst = 32'h10408000;
      14979: inst = 32'hc405005;
      14980: inst = 32'h8220000;
      14981: inst = 32'h10408000;
      14982: inst = 32'hc405006;
      14983: inst = 32'h8220000;
      14984: inst = 32'h10408000;
      14985: inst = 32'hc405007;
      14986: inst = 32'h8220000;
      14987: inst = 32'h10408000;
      14988: inst = 32'hc405009;
      14989: inst = 32'h8220000;
      14990: inst = 32'h10408000;
      14991: inst = 32'hc40500b;
      14992: inst = 32'h8220000;
      14993: inst = 32'h10408000;
      14994: inst = 32'hc40500d;
      14995: inst = 32'h8220000;
      14996: inst = 32'h10408000;
      14997: inst = 32'hc40500e;
      14998: inst = 32'h8220000;
      14999: inst = 32'h10408000;
      15000: inst = 32'hc40500f;
      15001: inst = 32'h8220000;
      15002: inst = 32'h10408000;
      15003: inst = 32'hc405010;
      15004: inst = 32'h8220000;
      15005: inst = 32'h10408000;
      15006: inst = 32'hc405011;
      15007: inst = 32'h8220000;
      15008: inst = 32'h10408000;
      15009: inst = 32'hc405012;
      15010: inst = 32'h8220000;
      15011: inst = 32'h10408000;
      15012: inst = 32'hc405013;
      15013: inst = 32'h8220000;
      15014: inst = 32'h10408000;
      15015: inst = 32'hc405061;
      15016: inst = 32'h8220000;
      15017: inst = 32'h10408000;
      15018: inst = 32'hc405062;
      15019: inst = 32'h8220000;
      15020: inst = 32'h10408000;
      15021: inst = 32'hc405063;
      15022: inst = 32'h8220000;
      15023: inst = 32'h10408000;
      15024: inst = 32'hc405064;
      15025: inst = 32'h8220000;
      15026: inst = 32'h10408000;
      15027: inst = 32'hc405065;
      15028: inst = 32'h8220000;
      15029: inst = 32'h10408000;
      15030: inst = 32'hc405066;
      15031: inst = 32'h8220000;
      15032: inst = 32'h10408000;
      15033: inst = 32'hc405067;
      15034: inst = 32'h8220000;
      15035: inst = 32'h10408000;
      15036: inst = 32'hc405068;
      15037: inst = 32'h8220000;
      15038: inst = 32'h10408000;
      15039: inst = 32'hc405069;
      15040: inst = 32'h8220000;
      15041: inst = 32'h10408000;
      15042: inst = 32'hc40506b;
      15043: inst = 32'h8220000;
      15044: inst = 32'h10408000;
      15045: inst = 32'hc40506c;
      15046: inst = 32'h8220000;
      15047: inst = 32'h10408000;
      15048: inst = 32'hc40506d;
      15049: inst = 32'h8220000;
      15050: inst = 32'h10408000;
      15051: inst = 32'hc40506e;
      15052: inst = 32'h8220000;
      15053: inst = 32'h10408000;
      15054: inst = 32'hc40506f;
      15055: inst = 32'h8220000;
      15056: inst = 32'h10408000;
      15057: inst = 32'hc405070;
      15058: inst = 32'h8220000;
      15059: inst = 32'h10408000;
      15060: inst = 32'hc405071;
      15061: inst = 32'h8220000;
      15062: inst = 32'h10408000;
      15063: inst = 32'hc405072;
      15064: inst = 32'h8220000;
      15065: inst = 32'h10408000;
      15066: inst = 32'hc405073;
      15067: inst = 32'h8220000;
      15068: inst = 32'h10408000;
      15069: inst = 32'hc4050c1;
      15070: inst = 32'h8220000;
      15071: inst = 32'h10408000;
      15072: inst = 32'hc4050c2;
      15073: inst = 32'h8220000;
      15074: inst = 32'h10408000;
      15075: inst = 32'hc4050c3;
      15076: inst = 32'h8220000;
      15077: inst = 32'h10408000;
      15078: inst = 32'hc4050c4;
      15079: inst = 32'h8220000;
      15080: inst = 32'h10408000;
      15081: inst = 32'hc4050c5;
      15082: inst = 32'h8220000;
      15083: inst = 32'h10408000;
      15084: inst = 32'hc4050c6;
      15085: inst = 32'h8220000;
      15086: inst = 32'h10408000;
      15087: inst = 32'hc4050c7;
      15088: inst = 32'h8220000;
      15089: inst = 32'h10408000;
      15090: inst = 32'hc4050c8;
      15091: inst = 32'h8220000;
      15092: inst = 32'h10408000;
      15093: inst = 32'hc4050c9;
      15094: inst = 32'h8220000;
      15095: inst = 32'h10408000;
      15096: inst = 32'hc4050cb;
      15097: inst = 32'h8220000;
      15098: inst = 32'h10408000;
      15099: inst = 32'hc4050cc;
      15100: inst = 32'h8220000;
      15101: inst = 32'h10408000;
      15102: inst = 32'hc4050cd;
      15103: inst = 32'h8220000;
      15104: inst = 32'h10408000;
      15105: inst = 32'hc4050ce;
      15106: inst = 32'h8220000;
      15107: inst = 32'h10408000;
      15108: inst = 32'hc4050cf;
      15109: inst = 32'h8220000;
      15110: inst = 32'h10408000;
      15111: inst = 32'hc4050d0;
      15112: inst = 32'h8220000;
      15113: inst = 32'h10408000;
      15114: inst = 32'hc4050d1;
      15115: inst = 32'h8220000;
      15116: inst = 32'h10408000;
      15117: inst = 32'hc4050d2;
      15118: inst = 32'h8220000;
      15119: inst = 32'h10408000;
      15120: inst = 32'hc4050d3;
      15121: inst = 32'h8220000;
      15122: inst = 32'h10408000;
      15123: inst = 32'hc405121;
      15124: inst = 32'h8220000;
      15125: inst = 32'h10408000;
      15126: inst = 32'hc405122;
      15127: inst = 32'h8220000;
      15128: inst = 32'h10408000;
      15129: inst = 32'hc405123;
      15130: inst = 32'h8220000;
      15131: inst = 32'h10408000;
      15132: inst = 32'hc405124;
      15133: inst = 32'h8220000;
      15134: inst = 32'h10408000;
      15135: inst = 32'hc405125;
      15136: inst = 32'h8220000;
      15137: inst = 32'h10408000;
      15138: inst = 32'hc405126;
      15139: inst = 32'h8220000;
      15140: inst = 32'h10408000;
      15141: inst = 32'hc405127;
      15142: inst = 32'h8220000;
      15143: inst = 32'h10408000;
      15144: inst = 32'hc405128;
      15145: inst = 32'h8220000;
      15146: inst = 32'h10408000;
      15147: inst = 32'hc405129;
      15148: inst = 32'h8220000;
      15149: inst = 32'h10408000;
      15150: inst = 32'hc40512b;
      15151: inst = 32'h8220000;
      15152: inst = 32'h10408000;
      15153: inst = 32'hc40512c;
      15154: inst = 32'h8220000;
      15155: inst = 32'h10408000;
      15156: inst = 32'hc40512d;
      15157: inst = 32'h8220000;
      15158: inst = 32'h10408000;
      15159: inst = 32'hc40512e;
      15160: inst = 32'h8220000;
      15161: inst = 32'h10408000;
      15162: inst = 32'hc40512f;
      15163: inst = 32'h8220000;
      15164: inst = 32'h10408000;
      15165: inst = 32'hc405130;
      15166: inst = 32'h8220000;
      15167: inst = 32'h10408000;
      15168: inst = 32'hc405131;
      15169: inst = 32'h8220000;
      15170: inst = 32'h10408000;
      15171: inst = 32'hc405132;
      15172: inst = 32'h8220000;
      15173: inst = 32'h10408000;
      15174: inst = 32'hc405133;
      15175: inst = 32'h8220000;
      15176: inst = 32'h10408000;
      15177: inst = 32'hc405181;
      15178: inst = 32'h8220000;
      15179: inst = 32'h10408000;
      15180: inst = 32'hc405182;
      15181: inst = 32'h8220000;
      15182: inst = 32'h10408000;
      15183: inst = 32'hc405183;
      15184: inst = 32'h8220000;
      15185: inst = 32'h10408000;
      15186: inst = 32'hc405184;
      15187: inst = 32'h8220000;
      15188: inst = 32'h10408000;
      15189: inst = 32'hc405185;
      15190: inst = 32'h8220000;
      15191: inst = 32'h10408000;
      15192: inst = 32'hc405186;
      15193: inst = 32'h8220000;
      15194: inst = 32'h10408000;
      15195: inst = 32'hc405187;
      15196: inst = 32'h8220000;
      15197: inst = 32'h10408000;
      15198: inst = 32'hc405188;
      15199: inst = 32'h8220000;
      15200: inst = 32'h10408000;
      15201: inst = 32'hc405189;
      15202: inst = 32'h8220000;
      15203: inst = 32'h10408000;
      15204: inst = 32'hc40518b;
      15205: inst = 32'h8220000;
      15206: inst = 32'h10408000;
      15207: inst = 32'hc40518c;
      15208: inst = 32'h8220000;
      15209: inst = 32'h10408000;
      15210: inst = 32'hc40518d;
      15211: inst = 32'h8220000;
      15212: inst = 32'h10408000;
      15213: inst = 32'hc40518e;
      15214: inst = 32'h8220000;
      15215: inst = 32'h10408000;
      15216: inst = 32'hc40518f;
      15217: inst = 32'h8220000;
      15218: inst = 32'h10408000;
      15219: inst = 32'hc405190;
      15220: inst = 32'h8220000;
      15221: inst = 32'h10408000;
      15222: inst = 32'hc405191;
      15223: inst = 32'h8220000;
      15224: inst = 32'h10408000;
      15225: inst = 32'hc405192;
      15226: inst = 32'h8220000;
      15227: inst = 32'h10408000;
      15228: inst = 32'hc405193;
      15229: inst = 32'h8220000;
      15230: inst = 32'h10408000;
      15231: inst = 32'hc4051e1;
      15232: inst = 32'h8220000;
      15233: inst = 32'h10408000;
      15234: inst = 32'hc4051e2;
      15235: inst = 32'h8220000;
      15236: inst = 32'h10408000;
      15237: inst = 32'hc4051e3;
      15238: inst = 32'h8220000;
      15239: inst = 32'h10408000;
      15240: inst = 32'hc4051e4;
      15241: inst = 32'h8220000;
      15242: inst = 32'h10408000;
      15243: inst = 32'hc4051e5;
      15244: inst = 32'h8220000;
      15245: inst = 32'h10408000;
      15246: inst = 32'hc4051e6;
      15247: inst = 32'h8220000;
      15248: inst = 32'h10408000;
      15249: inst = 32'hc4051e7;
      15250: inst = 32'h8220000;
      15251: inst = 32'h10408000;
      15252: inst = 32'hc4051e8;
      15253: inst = 32'h8220000;
      15254: inst = 32'h10408000;
      15255: inst = 32'hc4051e9;
      15256: inst = 32'h8220000;
      15257: inst = 32'h10408000;
      15258: inst = 32'hc4051eb;
      15259: inst = 32'h8220000;
      15260: inst = 32'h10408000;
      15261: inst = 32'hc4051ec;
      15262: inst = 32'h8220000;
      15263: inst = 32'h10408000;
      15264: inst = 32'hc4051ed;
      15265: inst = 32'h8220000;
      15266: inst = 32'h10408000;
      15267: inst = 32'hc4051ee;
      15268: inst = 32'h8220000;
      15269: inst = 32'h10408000;
      15270: inst = 32'hc4051ef;
      15271: inst = 32'h8220000;
      15272: inst = 32'h10408000;
      15273: inst = 32'hc4051f0;
      15274: inst = 32'h8220000;
      15275: inst = 32'h10408000;
      15276: inst = 32'hc4051f1;
      15277: inst = 32'h8220000;
      15278: inst = 32'h10408000;
      15279: inst = 32'hc4051f2;
      15280: inst = 32'h8220000;
      15281: inst = 32'h10408000;
      15282: inst = 32'hc4051f3;
      15283: inst = 32'h8220000;
      15284: inst = 32'h10408000;
      15285: inst = 32'hc405241;
      15286: inst = 32'h8220000;
      15287: inst = 32'h10408000;
      15288: inst = 32'hc405242;
      15289: inst = 32'h8220000;
      15290: inst = 32'h10408000;
      15291: inst = 32'hc405243;
      15292: inst = 32'h8220000;
      15293: inst = 32'h10408000;
      15294: inst = 32'hc405244;
      15295: inst = 32'h8220000;
      15296: inst = 32'h10408000;
      15297: inst = 32'hc405245;
      15298: inst = 32'h8220000;
      15299: inst = 32'h10408000;
      15300: inst = 32'hc405246;
      15301: inst = 32'h8220000;
      15302: inst = 32'h10408000;
      15303: inst = 32'hc405247;
      15304: inst = 32'h8220000;
      15305: inst = 32'h10408000;
      15306: inst = 32'hc405248;
      15307: inst = 32'h8220000;
      15308: inst = 32'h10408000;
      15309: inst = 32'hc405249;
      15310: inst = 32'h8220000;
      15311: inst = 32'h10408000;
      15312: inst = 32'hc40524b;
      15313: inst = 32'h8220000;
      15314: inst = 32'h10408000;
      15315: inst = 32'hc40524c;
      15316: inst = 32'h8220000;
      15317: inst = 32'h10408000;
      15318: inst = 32'hc40524d;
      15319: inst = 32'h8220000;
      15320: inst = 32'h10408000;
      15321: inst = 32'hc40524e;
      15322: inst = 32'h8220000;
      15323: inst = 32'h10408000;
      15324: inst = 32'hc40524f;
      15325: inst = 32'h8220000;
      15326: inst = 32'h10408000;
      15327: inst = 32'hc405250;
      15328: inst = 32'h8220000;
      15329: inst = 32'h10408000;
      15330: inst = 32'hc405251;
      15331: inst = 32'h8220000;
      15332: inst = 32'h10408000;
      15333: inst = 32'hc405252;
      15334: inst = 32'h8220000;
      15335: inst = 32'h10408000;
      15336: inst = 32'hc405253;
      15337: inst = 32'h8220000;
      15338: inst = 32'hc20bd73;
      15339: inst = 32'h10408000;
      15340: inst = 32'hc404e9f;
      15341: inst = 32'h8220000;
      15342: inst = 32'h10408000;
      15343: inst = 32'hc404ec0;
      15344: inst = 32'h8220000;
      15345: inst = 32'hc205aed;
      15346: inst = 32'h10408000;
      15347: inst = 32'hc404ea0;
      15348: inst = 32'h8220000;
      15349: inst = 32'h10408000;
      15350: inst = 32'hc404ea1;
      15351: inst = 32'h8220000;
      15352: inst = 32'h10408000;
      15353: inst = 32'hc404ea2;
      15354: inst = 32'h8220000;
      15355: inst = 32'h10408000;
      15356: inst = 32'hc404ea3;
      15357: inst = 32'h8220000;
      15358: inst = 32'h10408000;
      15359: inst = 32'hc404ea4;
      15360: inst = 32'h8220000;
      15361: inst = 32'h10408000;
      15362: inst = 32'hc404ebb;
      15363: inst = 32'h8220000;
      15364: inst = 32'h10408000;
      15365: inst = 32'hc404ebc;
      15366: inst = 32'h8220000;
      15367: inst = 32'h10408000;
      15368: inst = 32'hc404ebd;
      15369: inst = 32'h8220000;
      15370: inst = 32'h10408000;
      15371: inst = 32'hc404ebe;
      15372: inst = 32'h8220000;
      15373: inst = 32'h10408000;
      15374: inst = 32'hc404ebf;
      15375: inst = 32'h8220000;
      15376: inst = 32'h10408000;
      15377: inst = 32'hc404f00;
      15378: inst = 32'h8220000;
      15379: inst = 32'h10408000;
      15380: inst = 32'hc404f01;
      15381: inst = 32'h8220000;
      15382: inst = 32'h10408000;
      15383: inst = 32'hc404f02;
      15384: inst = 32'h8220000;
      15385: inst = 32'h10408000;
      15386: inst = 32'hc404f03;
      15387: inst = 32'h8220000;
      15388: inst = 32'h10408000;
      15389: inst = 32'hc404f04;
      15390: inst = 32'h8220000;
      15391: inst = 32'h10408000;
      15392: inst = 32'hc404f05;
      15393: inst = 32'h8220000;
      15394: inst = 32'h10408000;
      15395: inst = 32'hc404f1a;
      15396: inst = 32'h8220000;
      15397: inst = 32'h10408000;
      15398: inst = 32'hc404f1b;
      15399: inst = 32'h8220000;
      15400: inst = 32'h10408000;
      15401: inst = 32'hc404f1c;
      15402: inst = 32'h8220000;
      15403: inst = 32'h10408000;
      15404: inst = 32'hc404f1d;
      15405: inst = 32'h8220000;
      15406: inst = 32'h10408000;
      15407: inst = 32'hc404f1e;
      15408: inst = 32'h8220000;
      15409: inst = 32'h10408000;
      15410: inst = 32'hc404f1f;
      15411: inst = 32'h8220000;
      15412: inst = 32'h10408000;
      15413: inst = 32'hc404f60;
      15414: inst = 32'h8220000;
      15415: inst = 32'h10408000;
      15416: inst = 32'hc404f61;
      15417: inst = 32'h8220000;
      15418: inst = 32'h10408000;
      15419: inst = 32'hc404f62;
      15420: inst = 32'h8220000;
      15421: inst = 32'h10408000;
      15422: inst = 32'hc404f63;
      15423: inst = 32'h8220000;
      15424: inst = 32'h10408000;
      15425: inst = 32'hc404f64;
      15426: inst = 32'h8220000;
      15427: inst = 32'h10408000;
      15428: inst = 32'hc404f65;
      15429: inst = 32'h8220000;
      15430: inst = 32'h10408000;
      15431: inst = 32'hc404f66;
      15432: inst = 32'h8220000;
      15433: inst = 32'h10408000;
      15434: inst = 32'hc404f67;
      15435: inst = 32'h8220000;
      15436: inst = 32'h10408000;
      15437: inst = 32'hc404f78;
      15438: inst = 32'h8220000;
      15439: inst = 32'h10408000;
      15440: inst = 32'hc404f79;
      15441: inst = 32'h8220000;
      15442: inst = 32'h10408000;
      15443: inst = 32'hc404f7a;
      15444: inst = 32'h8220000;
      15445: inst = 32'h10408000;
      15446: inst = 32'hc404f7b;
      15447: inst = 32'h8220000;
      15448: inst = 32'h10408000;
      15449: inst = 32'hc404f7c;
      15450: inst = 32'h8220000;
      15451: inst = 32'h10408000;
      15452: inst = 32'hc404f7d;
      15453: inst = 32'h8220000;
      15454: inst = 32'h10408000;
      15455: inst = 32'hc404f7e;
      15456: inst = 32'h8220000;
      15457: inst = 32'h10408000;
      15458: inst = 32'hc404f7f;
      15459: inst = 32'h8220000;
      15460: inst = 32'h10408000;
      15461: inst = 32'hc404fc0;
      15462: inst = 32'h8220000;
      15463: inst = 32'h10408000;
      15464: inst = 32'hc404fc1;
      15465: inst = 32'h8220000;
      15466: inst = 32'h10408000;
      15467: inst = 32'hc404fc2;
      15468: inst = 32'h8220000;
      15469: inst = 32'h10408000;
      15470: inst = 32'hc404fc3;
      15471: inst = 32'h8220000;
      15472: inst = 32'h10408000;
      15473: inst = 32'hc404fc4;
      15474: inst = 32'h8220000;
      15475: inst = 32'h10408000;
      15476: inst = 32'hc404fc6;
      15477: inst = 32'h8220000;
      15478: inst = 32'h10408000;
      15479: inst = 32'hc404fc7;
      15480: inst = 32'h8220000;
      15481: inst = 32'h10408000;
      15482: inst = 32'hc404fd8;
      15483: inst = 32'h8220000;
      15484: inst = 32'h10408000;
      15485: inst = 32'hc404fd9;
      15486: inst = 32'h8220000;
      15487: inst = 32'h10408000;
      15488: inst = 32'hc404fdb;
      15489: inst = 32'h8220000;
      15490: inst = 32'h10408000;
      15491: inst = 32'hc404fdc;
      15492: inst = 32'h8220000;
      15493: inst = 32'h10408000;
      15494: inst = 32'hc404fdd;
      15495: inst = 32'h8220000;
      15496: inst = 32'h10408000;
      15497: inst = 32'hc404fde;
      15498: inst = 32'h8220000;
      15499: inst = 32'h10408000;
      15500: inst = 32'hc404fdf;
      15501: inst = 32'h8220000;
      15502: inst = 32'h10408000;
      15503: inst = 32'hc405020;
      15504: inst = 32'h8220000;
      15505: inst = 32'h10408000;
      15506: inst = 32'hc405021;
      15507: inst = 32'h8220000;
      15508: inst = 32'h10408000;
      15509: inst = 32'hc405022;
      15510: inst = 32'h8220000;
      15511: inst = 32'h10408000;
      15512: inst = 32'hc405023;
      15513: inst = 32'h8220000;
      15514: inst = 32'h10408000;
      15515: inst = 32'hc405026;
      15516: inst = 32'h8220000;
      15517: inst = 32'h10408000;
      15518: inst = 32'hc405027;
      15519: inst = 32'h8220000;
      15520: inst = 32'h10408000;
      15521: inst = 32'hc405038;
      15522: inst = 32'h8220000;
      15523: inst = 32'h10408000;
      15524: inst = 32'hc405039;
      15525: inst = 32'h8220000;
      15526: inst = 32'h10408000;
      15527: inst = 32'hc40503c;
      15528: inst = 32'h8220000;
      15529: inst = 32'h10408000;
      15530: inst = 32'hc40503d;
      15531: inst = 32'h8220000;
      15532: inst = 32'h10408000;
      15533: inst = 32'hc40503e;
      15534: inst = 32'h8220000;
      15535: inst = 32'h10408000;
      15536: inst = 32'hc40503f;
      15537: inst = 32'h8220000;
      15538: inst = 32'h10408000;
      15539: inst = 32'hc40507f;
      15540: inst = 32'h8220000;
      15541: inst = 32'h10408000;
      15542: inst = 32'hc405080;
      15543: inst = 32'h8220000;
      15544: inst = 32'h10408000;
      15545: inst = 32'hc405081;
      15546: inst = 32'h8220000;
      15547: inst = 32'h10408000;
      15548: inst = 32'hc405082;
      15549: inst = 32'h8220000;
      15550: inst = 32'h10408000;
      15551: inst = 32'hc405086;
      15552: inst = 32'h8220000;
      15553: inst = 32'h10408000;
      15554: inst = 32'hc405087;
      15555: inst = 32'h8220000;
      15556: inst = 32'h10408000;
      15557: inst = 32'hc405098;
      15558: inst = 32'h8220000;
      15559: inst = 32'h10408000;
      15560: inst = 32'hc405099;
      15561: inst = 32'h8220000;
      15562: inst = 32'h10408000;
      15563: inst = 32'hc40509d;
      15564: inst = 32'h8220000;
      15565: inst = 32'h10408000;
      15566: inst = 32'hc40509e;
      15567: inst = 32'h8220000;
      15568: inst = 32'h10408000;
      15569: inst = 32'hc40509f;
      15570: inst = 32'h8220000;
      15571: inst = 32'h10408000;
      15572: inst = 32'hc4050a0;
      15573: inst = 32'h8220000;
      15574: inst = 32'h10408000;
      15575: inst = 32'hc4050df;
      15576: inst = 32'h8220000;
      15577: inst = 32'h10408000;
      15578: inst = 32'hc4050e0;
      15579: inst = 32'h8220000;
      15580: inst = 32'h10408000;
      15581: inst = 32'hc4050e1;
      15582: inst = 32'h8220000;
      15583: inst = 32'h10408000;
      15584: inst = 32'hc4050e2;
      15585: inst = 32'h8220000;
      15586: inst = 32'h10408000;
      15587: inst = 32'hc4050e6;
      15588: inst = 32'h8220000;
      15589: inst = 32'h10408000;
      15590: inst = 32'hc4050e7;
      15591: inst = 32'h8220000;
      15592: inst = 32'h10408000;
      15593: inst = 32'hc4050f8;
      15594: inst = 32'h8220000;
      15595: inst = 32'h10408000;
      15596: inst = 32'hc4050f9;
      15597: inst = 32'h8220000;
      15598: inst = 32'h10408000;
      15599: inst = 32'hc4050fd;
      15600: inst = 32'h8220000;
      15601: inst = 32'h10408000;
      15602: inst = 32'hc4050fe;
      15603: inst = 32'h8220000;
      15604: inst = 32'h10408000;
      15605: inst = 32'hc4050ff;
      15606: inst = 32'h8220000;
      15607: inst = 32'h10408000;
      15608: inst = 32'hc405100;
      15609: inst = 32'h8220000;
      15610: inst = 32'h10408000;
      15611: inst = 32'hc40513f;
      15612: inst = 32'h8220000;
      15613: inst = 32'h10408000;
      15614: inst = 32'hc405140;
      15615: inst = 32'h8220000;
      15616: inst = 32'h10408000;
      15617: inst = 32'hc405141;
      15618: inst = 32'h8220000;
      15619: inst = 32'h10408000;
      15620: inst = 32'hc405146;
      15621: inst = 32'h8220000;
      15622: inst = 32'h10408000;
      15623: inst = 32'hc405147;
      15624: inst = 32'h8220000;
      15625: inst = 32'h10408000;
      15626: inst = 32'hc405158;
      15627: inst = 32'h8220000;
      15628: inst = 32'h10408000;
      15629: inst = 32'hc405159;
      15630: inst = 32'h8220000;
      15631: inst = 32'h10408000;
      15632: inst = 32'hc40515e;
      15633: inst = 32'h8220000;
      15634: inst = 32'h10408000;
      15635: inst = 32'hc40515f;
      15636: inst = 32'h8220000;
      15637: inst = 32'h10408000;
      15638: inst = 32'hc405160;
      15639: inst = 32'h8220000;
      15640: inst = 32'h10408000;
      15641: inst = 32'hc40519f;
      15642: inst = 32'h8220000;
      15643: inst = 32'h10408000;
      15644: inst = 32'hc4051a0;
      15645: inst = 32'h8220000;
      15646: inst = 32'h10408000;
      15647: inst = 32'hc4051a6;
      15648: inst = 32'h8220000;
      15649: inst = 32'h10408000;
      15650: inst = 32'hc4051a7;
      15651: inst = 32'h8220000;
      15652: inst = 32'h10408000;
      15653: inst = 32'hc4051b8;
      15654: inst = 32'h8220000;
      15655: inst = 32'h10408000;
      15656: inst = 32'hc4051b9;
      15657: inst = 32'h8220000;
      15658: inst = 32'h10408000;
      15659: inst = 32'hc4051bf;
      15660: inst = 32'h8220000;
      15661: inst = 32'h10408000;
      15662: inst = 32'hc4051c0;
      15663: inst = 32'h8220000;
      15664: inst = 32'h10408000;
      15665: inst = 32'hc4051ff;
      15666: inst = 32'h8220000;
      15667: inst = 32'h10408000;
      15668: inst = 32'hc405200;
      15669: inst = 32'h8220000;
      15670: inst = 32'h10408000;
      15671: inst = 32'hc405206;
      15672: inst = 32'h8220000;
      15673: inst = 32'h10408000;
      15674: inst = 32'hc405207;
      15675: inst = 32'h8220000;
      15676: inst = 32'h10408000;
      15677: inst = 32'hc405218;
      15678: inst = 32'h8220000;
      15679: inst = 32'h10408000;
      15680: inst = 32'hc405219;
      15681: inst = 32'h8220000;
      15682: inst = 32'h10408000;
      15683: inst = 32'hc40521f;
      15684: inst = 32'h8220000;
      15685: inst = 32'h10408000;
      15686: inst = 32'hc405220;
      15687: inst = 32'h8220000;
      15688: inst = 32'h10408000;
      15689: inst = 32'hc40525f;
      15690: inst = 32'h8220000;
      15691: inst = 32'h10408000;
      15692: inst = 32'hc405260;
      15693: inst = 32'h8220000;
      15694: inst = 32'h10408000;
      15695: inst = 32'hc405266;
      15696: inst = 32'h8220000;
      15697: inst = 32'h10408000;
      15698: inst = 32'hc405267;
      15699: inst = 32'h8220000;
      15700: inst = 32'h10408000;
      15701: inst = 32'hc405278;
      15702: inst = 32'h8220000;
      15703: inst = 32'h10408000;
      15704: inst = 32'hc405279;
      15705: inst = 32'h8220000;
      15706: inst = 32'h10408000;
      15707: inst = 32'hc40527f;
      15708: inst = 32'h8220000;
      15709: inst = 32'h10408000;
      15710: inst = 32'hc405280;
      15711: inst = 32'h8220000;
      15712: inst = 32'h10408000;
      15713: inst = 32'hc4052bf;
      15714: inst = 32'h8220000;
      15715: inst = 32'h10408000;
      15716: inst = 32'hc4052c0;
      15717: inst = 32'h8220000;
      15718: inst = 32'h10408000;
      15719: inst = 32'hc4052c6;
      15720: inst = 32'h8220000;
      15721: inst = 32'h10408000;
      15722: inst = 32'hc4052c7;
      15723: inst = 32'h8220000;
      15724: inst = 32'h10408000;
      15725: inst = 32'hc4052d8;
      15726: inst = 32'h8220000;
      15727: inst = 32'h10408000;
      15728: inst = 32'hc4052d9;
      15729: inst = 32'h8220000;
      15730: inst = 32'h10408000;
      15731: inst = 32'hc4052df;
      15732: inst = 32'h8220000;
      15733: inst = 32'h10408000;
      15734: inst = 32'hc4052e0;
      15735: inst = 32'h8220000;
      15736: inst = 32'hc207bae;
      15737: inst = 32'h10408000;
      15738: inst = 32'hc404ea5;
      15739: inst = 32'h8220000;
      15740: inst = 32'h10408000;
      15741: inst = 32'hc404eba;
      15742: inst = 32'h8220000;
      15743: inst = 32'hc20c5b4;
      15744: inst = 32'h10408000;
      15745: inst = 32'hc404ea6;
      15746: inst = 32'h8220000;
      15747: inst = 32'h10408000;
      15748: inst = 32'hc404eb9;
      15749: inst = 32'h8220000;
      15750: inst = 32'hc20d5f4;
      15751: inst = 32'h10408000;
      15752: inst = 32'hc404ea7;
      15753: inst = 32'h8220000;
      15754: inst = 32'h10408000;
      15755: inst = 32'hc404eb8;
      15756: inst = 32'h8220000;
      15757: inst = 32'hc20a4b1;
      15758: inst = 32'h10408000;
      15759: inst = 32'hc404eff;
      15760: inst = 32'h8220000;
      15761: inst = 32'h10408000;
      15762: inst = 32'hc404f20;
      15763: inst = 32'h8220000;
      15764: inst = 32'h10408000;
      15765: inst = 32'hc404fbf;
      15766: inst = 32'h8220000;
      15767: inst = 32'h10408000;
      15768: inst = 32'hc404fe0;
      15769: inst = 32'h8220000;
      15770: inst = 32'hc2062ed;
      15771: inst = 32'h10408000;
      15772: inst = 32'hc404f06;
      15773: inst = 32'h8220000;
      15774: inst = 32'h10408000;
      15775: inst = 32'hc404f19;
      15776: inst = 32'h8220000;
      15777: inst = 32'hc209450;
      15778: inst = 32'h10408000;
      15779: inst = 32'hc404f07;
      15780: inst = 32'h8220000;
      15781: inst = 32'h10408000;
      15782: inst = 32'hc404f18;
      15783: inst = 32'h8220000;
      15784: inst = 32'h10408000;
      15785: inst = 32'hc405209;
      15786: inst = 32'h8220000;
      15787: inst = 32'h10408000;
      15788: inst = 32'hc405216;
      15789: inst = 32'h8220000;
      15790: inst = 32'hc20a4d1;
      15791: inst = 32'h10408000;
      15792: inst = 32'hc404f5f;
      15793: inst = 32'h8220000;
      15794: inst = 32'h10408000;
      15795: inst = 32'hc404f80;
      15796: inst = 32'h8220000;
      15797: inst = 32'hc204a49;
      15798: inst = 32'h10408000;
      15799: inst = 32'hc404fa8;
      15800: inst = 32'h8220000;
      15801: inst = 32'h10408000;
      15802: inst = 32'hc404fac;
      15803: inst = 32'h8220000;
      15804: inst = 32'h10408000;
      15805: inst = 32'hc405008;
      15806: inst = 32'h8220000;
      15807: inst = 32'h10408000;
      15808: inst = 32'hc40500c;
      15809: inst = 32'h8220000;
      15810: inst = 32'hc205acb;
      15811: inst = 32'h10408000;
      15812: inst = 32'hc404fc5;
      15813: inst = 32'h8220000;
      15814: inst = 32'h10408000;
      15815: inst = 32'hc404fda;
      15816: inst = 32'h8220000;
      15817: inst = 32'h10408000;
      15818: inst = 32'hc405336;
      15819: inst = 32'h8220000;
      15820: inst = 32'h10408000;
      15821: inst = 32'hc405380;
      15822: inst = 32'h8220000;
      15823: inst = 32'h10408000;
      15824: inst = 32'hc40539f;
      15825: inst = 32'h8220000;
      15826: inst = 32'h10408000;
      15827: inst = 32'hc4053dd;
      15828: inst = 32'h8220000;
      15829: inst = 32'h10408000;
      15830: inst = 32'hc405402;
      15831: inst = 32'h8220000;
      15832: inst = 32'hc20630d;
      15833: inst = 32'h10408000;
      15834: inst = 32'hc40501f;
      15835: inst = 32'h8220000;
      15836: inst = 32'h10408000;
      15837: inst = 32'hc405040;
      15838: inst = 32'h8220000;
      15839: inst = 32'hc205aec;
      15840: inst = 32'h10408000;
      15841: inst = 32'hc405024;
      15842: inst = 32'h8220000;
      15843: inst = 32'h10408000;
      15844: inst = 32'hc40503b;
      15845: inst = 32'h8220000;
      15846: inst = 32'h10408000;
      15847: inst = 32'hc405083;
      15848: inst = 32'h8220000;
      15849: inst = 32'h10408000;
      15850: inst = 32'hc40509c;
      15851: inst = 32'h8220000;
      15852: inst = 32'h10408000;
      15853: inst = 32'hc4051a1;
      15854: inst = 32'h8220000;
      15855: inst = 32'h10408000;
      15856: inst = 32'hc4051be;
      15857: inst = 32'h8220000;
      15858: inst = 32'h10408000;
      15859: inst = 32'hc405329;
      15860: inst = 32'h8220000;
      15861: inst = 32'h10408000;
      15862: inst = 32'hc405568;
      15863: inst = 32'h8220000;
      15864: inst = 32'h10408000;
      15865: inst = 32'hc405577;
      15866: inst = 32'h8220000;
      15867: inst = 32'h10408000;
      15868: inst = 32'hc4057a7;
      15869: inst = 32'h8220000;
      15870: inst = 32'h10408000;
      15871: inst = 32'hc4057b8;
      15872: inst = 32'h8220000;
      15873: inst = 32'hc205269;
      15874: inst = 32'h10408000;
      15875: inst = 32'hc405025;
      15876: inst = 32'h8220000;
      15877: inst = 32'h10408000;
      15878: inst = 32'hc40503a;
      15879: inst = 32'h8220000;
      15880: inst = 32'h10408000;
      15881: inst = 32'hc40537e;
      15882: inst = 32'h8220000;
      15883: inst = 32'h10408000;
      15884: inst = 32'hc4053a1;
      15885: inst = 32'h8220000;
      15886: inst = 32'h10408000;
      15887: inst = 32'hc40549c;
      15888: inst = 32'h8220000;
      15889: inst = 32'h10408000;
      15890: inst = 32'hc4054c3;
      15891: inst = 32'h8220000;
      15892: inst = 32'hc20528a;
      15893: inst = 32'h10408000;
      15894: inst = 32'hc405084;
      15895: inst = 32'h8220000;
      15896: inst = 32'h10408000;
      15897: inst = 32'hc40509b;
      15898: inst = 32'h8220000;
      15899: inst = 32'h10408000;
      15900: inst = 32'hc4050e3;
      15901: inst = 32'h8220000;
      15902: inst = 32'h10408000;
      15903: inst = 32'hc4050fc;
      15904: inst = 32'h8220000;
      15905: inst = 32'h10408000;
      15906: inst = 32'hc4052c5;
      15907: inst = 32'h8220000;
      15908: inst = 32'h10408000;
      15909: inst = 32'hc4052da;
      15910: inst = 32'h8220000;
      15911: inst = 32'h10408000;
      15912: inst = 32'hc4053e9;
      15913: inst = 32'h8220000;
      15914: inst = 32'h10408000;
      15915: inst = 32'hc4053f6;
      15916: inst = 32'h8220000;
      15917: inst = 32'h10408000;
      15918: inst = 32'hc405449;
      15919: inst = 32'h8220000;
      15920: inst = 32'h10408000;
      15921: inst = 32'hc405456;
      15922: inst = 32'h8220000;
      15923: inst = 32'h10408000;
      15924: inst = 32'hc4054a9;
      15925: inst = 32'h8220000;
      15926: inst = 32'h10408000;
      15927: inst = 32'hc4054b6;
      15928: inst = 32'h8220000;
      15929: inst = 32'h10408000;
      15930: inst = 32'hc405509;
      15931: inst = 32'h8220000;
      15932: inst = 32'h10408000;
      15933: inst = 32'hc405516;
      15934: inst = 32'h8220000;
      15935: inst = 32'h10408000;
      15936: inst = 32'hc40555e;
      15937: inst = 32'h8220000;
      15938: inst = 32'h10408000;
      15939: inst = 32'hc405569;
      15940: inst = 32'h8220000;
      15941: inst = 32'h10408000;
      15942: inst = 32'hc405576;
      15943: inst = 32'h8220000;
      15944: inst = 32'h10408000;
      15945: inst = 32'hc405581;
      15946: inst = 32'h8220000;
      15947: inst = 32'h10408000;
      15948: inst = 32'hc4055c9;
      15949: inst = 32'h8220000;
      15950: inst = 32'h10408000;
      15951: inst = 32'hc4055d6;
      15952: inst = 32'h8220000;
      15953: inst = 32'h10408000;
      15954: inst = 32'hc405628;
      15955: inst = 32'h8220000;
      15956: inst = 32'h10408000;
      15957: inst = 32'hc405629;
      15958: inst = 32'h8220000;
      15959: inst = 32'h10408000;
      15960: inst = 32'hc405636;
      15961: inst = 32'h8220000;
      15962: inst = 32'h10408000;
      15963: inst = 32'hc405637;
      15964: inst = 32'h8220000;
      15965: inst = 32'h10408000;
      15966: inst = 32'hc40567d;
      15967: inst = 32'h8220000;
      15968: inst = 32'h10408000;
      15969: inst = 32'hc405688;
      15970: inst = 32'h8220000;
      15971: inst = 32'h10408000;
      15972: inst = 32'hc405689;
      15973: inst = 32'h8220000;
      15974: inst = 32'h10408000;
      15975: inst = 32'hc405696;
      15976: inst = 32'h8220000;
      15977: inst = 32'h10408000;
      15978: inst = 32'hc405697;
      15979: inst = 32'h8220000;
      15980: inst = 32'h10408000;
      15981: inst = 32'hc4056a2;
      15982: inst = 32'h8220000;
      15983: inst = 32'h10408000;
      15984: inst = 32'hc4056e8;
      15985: inst = 32'h8220000;
      15986: inst = 32'h10408000;
      15987: inst = 32'hc4056e9;
      15988: inst = 32'h8220000;
      15989: inst = 32'h10408000;
      15990: inst = 32'hc4056f6;
      15991: inst = 32'h8220000;
      15992: inst = 32'h10408000;
      15993: inst = 32'hc4056f7;
      15994: inst = 32'h8220000;
      15995: inst = 32'h10408000;
      15996: inst = 32'hc405748;
      15997: inst = 32'h8220000;
      15998: inst = 32'h10408000;
      15999: inst = 32'hc405749;
      16000: inst = 32'h8220000;
      16001: inst = 32'h10408000;
      16002: inst = 32'hc405756;
      16003: inst = 32'h8220000;
      16004: inst = 32'h10408000;
      16005: inst = 32'hc405757;
      16006: inst = 32'h8220000;
      16007: inst = 32'h10408000;
      16008: inst = 32'hc4057a8;
      16009: inst = 32'h8220000;
      16010: inst = 32'h10408000;
      16011: inst = 32'hc4057a9;
      16012: inst = 32'h8220000;
      16013: inst = 32'h10408000;
      16014: inst = 32'hc4057b6;
      16015: inst = 32'h8220000;
      16016: inst = 32'h10408000;
      16017: inst = 32'hc4057b7;
      16018: inst = 32'h8220000;
      16019: inst = 32'hc205aab;
      16020: inst = 32'h10408000;
      16021: inst = 32'hc405142;
      16022: inst = 32'h8220000;
      16023: inst = 32'h10408000;
      16024: inst = 32'hc40515d;
      16025: inst = 32'h8220000;
      16026: inst = 32'hc20cdd4;
      16027: inst = 32'h10408000;
      16028: inst = 32'hc40519e;
      16029: inst = 32'h8220000;
      16030: inst = 32'h10408000;
      16031: inst = 32'hc4051c1;
      16032: inst = 32'h8220000;
      16033: inst = 32'hc209471;
      16034: inst = 32'h10408000;
      16035: inst = 32'hc4051b6;
      16036: inst = 32'h8220000;
      16037: inst = 32'hc20de55;
      16038: inst = 32'h10408000;
      16039: inst = 32'hc4051fd;
      16040: inst = 32'h8220000;
      16041: inst = 32'h10408000;
      16042: inst = 32'hc405222;
      16043: inst = 32'h8220000;
      16044: inst = 32'hc209492;
      16045: inst = 32'h10408000;
      16046: inst = 32'hc4051fe;
      16047: inst = 32'h8220000;
      16048: inst = 32'h10408000;
      16049: inst = 32'hc405221;
      16050: inst = 32'h8220000;
      16051: inst = 32'hc205acc;
      16052: inst = 32'h10408000;
      16053: inst = 32'hc405201;
      16054: inst = 32'h8220000;
      16055: inst = 32'h10408000;
      16056: inst = 32'hc40521e;
      16057: inst = 32'h8220000;
      16058: inst = 32'h10408000;
      16059: inst = 32'hc405261;
      16060: inst = 32'h8220000;
      16061: inst = 32'h10408000;
      16062: inst = 32'hc40527e;
      16063: inst = 32'h8220000;
      16064: inst = 32'h10408000;
      16065: inst = 32'hc4052c1;
      16066: inst = 32'h8220000;
      16067: inst = 32'h10408000;
      16068: inst = 32'hc4052de;
      16069: inst = 32'h8220000;
      16070: inst = 32'hc20e696;
      16071: inst = 32'h10408000;
      16072: inst = 32'hc40525c;
      16073: inst = 32'h8220000;
      16074: inst = 32'h10408000;
      16075: inst = 32'hc405283;
      16076: inst = 32'h8220000;
      16077: inst = 32'hc209cb2;
      16078: inst = 32'h10408000;
      16079: inst = 32'hc40525d;
      16080: inst = 32'h8220000;
      16081: inst = 32'h10408000;
      16082: inst = 32'hc405282;
      16083: inst = 32'h8220000;
      16084: inst = 32'hc208c2f;
      16085: inst = 32'h10408000;
      16086: inst = 32'hc405269;
      16087: inst = 32'h8220000;
      16088: inst = 32'h10408000;
      16089: inst = 32'hc405276;
      16090: inst = 32'h8220000;
      16091: inst = 32'hc20ad33;
      16092: inst = 32'h10408000;
      16093: inst = 32'hc4052bc;
      16094: inst = 32'h8220000;
      16095: inst = 32'h10408000;
      16096: inst = 32'hc4052e3;
      16097: inst = 32'h8220000;
      16098: inst = 32'hc2083ee;
      16099: inst = 32'h10408000;
      16100: inst = 32'hc4052c9;
      16101: inst = 32'h8220000;
      16102: inst = 32'h10408000;
      16103: inst = 32'hc4052d6;
      16104: inst = 32'h8220000;
      16105: inst = 32'hc206b50;
      16106: inst = 32'h10408000;
      16107: inst = 32'hc405300;
      16108: inst = 32'h8220000;
      16109: inst = 32'h10408000;
      16110: inst = 32'hc405301;
      16111: inst = 32'h8220000;
      16112: inst = 32'h10408000;
      16113: inst = 32'hc405302;
      16114: inst = 32'h8220000;
      16115: inst = 32'h10408000;
      16116: inst = 32'hc405303;
      16117: inst = 32'h8220000;
      16118: inst = 32'h10408000;
      16119: inst = 32'hc405304;
      16120: inst = 32'h8220000;
      16121: inst = 32'h10408000;
      16122: inst = 32'hc405305;
      16123: inst = 32'h8220000;
      16124: inst = 32'h10408000;
      16125: inst = 32'hc405306;
      16126: inst = 32'h8220000;
      16127: inst = 32'h10408000;
      16128: inst = 32'hc405307;
      16129: inst = 32'h8220000;
      16130: inst = 32'h10408000;
      16131: inst = 32'hc405308;
      16132: inst = 32'h8220000;
      16133: inst = 32'h10408000;
      16134: inst = 32'hc405309;
      16135: inst = 32'h8220000;
      16136: inst = 32'h10408000;
      16137: inst = 32'hc40530a;
      16138: inst = 32'h8220000;
      16139: inst = 32'h10408000;
      16140: inst = 32'hc40530b;
      16141: inst = 32'h8220000;
      16142: inst = 32'h10408000;
      16143: inst = 32'hc40530c;
      16144: inst = 32'h8220000;
      16145: inst = 32'h10408000;
      16146: inst = 32'hc40530d;
      16147: inst = 32'h8220000;
      16148: inst = 32'h10408000;
      16149: inst = 32'hc40530e;
      16150: inst = 32'h8220000;
      16151: inst = 32'h10408000;
      16152: inst = 32'hc40530f;
      16153: inst = 32'h8220000;
      16154: inst = 32'h10408000;
      16155: inst = 32'hc405310;
      16156: inst = 32'h8220000;
      16157: inst = 32'h10408000;
      16158: inst = 32'hc405311;
      16159: inst = 32'h8220000;
      16160: inst = 32'h10408000;
      16161: inst = 32'hc405312;
      16162: inst = 32'h8220000;
      16163: inst = 32'h10408000;
      16164: inst = 32'hc405313;
      16165: inst = 32'h8220000;
      16166: inst = 32'h10408000;
      16167: inst = 32'hc405314;
      16168: inst = 32'h8220000;
      16169: inst = 32'h10408000;
      16170: inst = 32'hc405315;
      16171: inst = 32'h8220000;
      16172: inst = 32'h10408000;
      16173: inst = 32'hc405316;
      16174: inst = 32'h8220000;
      16175: inst = 32'h10408000;
      16176: inst = 32'hc405317;
      16177: inst = 32'h8220000;
      16178: inst = 32'h10408000;
      16179: inst = 32'hc405318;
      16180: inst = 32'h8220000;
      16181: inst = 32'h10408000;
      16182: inst = 32'hc405319;
      16183: inst = 32'h8220000;
      16184: inst = 32'h10408000;
      16185: inst = 32'hc40531a;
      16186: inst = 32'h8220000;
      16187: inst = 32'h10408000;
      16188: inst = 32'hc40532a;
      16189: inst = 32'h8220000;
      16190: inst = 32'h10408000;
      16191: inst = 32'hc40532b;
      16192: inst = 32'h8220000;
      16193: inst = 32'h10408000;
      16194: inst = 32'hc40532c;
      16195: inst = 32'h8220000;
      16196: inst = 32'h10408000;
      16197: inst = 32'hc40532d;
      16198: inst = 32'h8220000;
      16199: inst = 32'h10408000;
      16200: inst = 32'hc40532e;
      16201: inst = 32'h8220000;
      16202: inst = 32'h10408000;
      16203: inst = 32'hc40532f;
      16204: inst = 32'h8220000;
      16205: inst = 32'h10408000;
      16206: inst = 32'hc405330;
      16207: inst = 32'h8220000;
      16208: inst = 32'h10408000;
      16209: inst = 32'hc405331;
      16210: inst = 32'h8220000;
      16211: inst = 32'h10408000;
      16212: inst = 32'hc405332;
      16213: inst = 32'h8220000;
      16214: inst = 32'h10408000;
      16215: inst = 32'hc405333;
      16216: inst = 32'h8220000;
      16217: inst = 32'h10408000;
      16218: inst = 32'hc405334;
      16219: inst = 32'h8220000;
      16220: inst = 32'h10408000;
      16221: inst = 32'hc405335;
      16222: inst = 32'h8220000;
      16223: inst = 32'h10408000;
      16224: inst = 32'hc405345;
      16225: inst = 32'h8220000;
      16226: inst = 32'h10408000;
      16227: inst = 32'hc405346;
      16228: inst = 32'h8220000;
      16229: inst = 32'h10408000;
      16230: inst = 32'hc405347;
      16231: inst = 32'h8220000;
      16232: inst = 32'h10408000;
      16233: inst = 32'hc405348;
      16234: inst = 32'h8220000;
      16235: inst = 32'h10408000;
      16236: inst = 32'hc405349;
      16237: inst = 32'h8220000;
      16238: inst = 32'h10408000;
      16239: inst = 32'hc40534a;
      16240: inst = 32'h8220000;
      16241: inst = 32'h10408000;
      16242: inst = 32'hc40534b;
      16243: inst = 32'h8220000;
      16244: inst = 32'h10408000;
      16245: inst = 32'hc40534c;
      16246: inst = 32'h8220000;
      16247: inst = 32'h10408000;
      16248: inst = 32'hc40534d;
      16249: inst = 32'h8220000;
      16250: inst = 32'h10408000;
      16251: inst = 32'hc40534e;
      16252: inst = 32'h8220000;
      16253: inst = 32'h10408000;
      16254: inst = 32'hc40534f;
      16255: inst = 32'h8220000;
      16256: inst = 32'h10408000;
      16257: inst = 32'hc405350;
      16258: inst = 32'h8220000;
      16259: inst = 32'h10408000;
      16260: inst = 32'hc405351;
      16261: inst = 32'h8220000;
      16262: inst = 32'h10408000;
      16263: inst = 32'hc405352;
      16264: inst = 32'h8220000;
      16265: inst = 32'h10408000;
      16266: inst = 32'hc405353;
      16267: inst = 32'h8220000;
      16268: inst = 32'h10408000;
      16269: inst = 32'hc405354;
      16270: inst = 32'h8220000;
      16271: inst = 32'h10408000;
      16272: inst = 32'hc405355;
      16273: inst = 32'h8220000;
      16274: inst = 32'h10408000;
      16275: inst = 32'hc405356;
      16276: inst = 32'h8220000;
      16277: inst = 32'h10408000;
      16278: inst = 32'hc405357;
      16279: inst = 32'h8220000;
      16280: inst = 32'h10408000;
      16281: inst = 32'hc405358;
      16282: inst = 32'h8220000;
      16283: inst = 32'h10408000;
      16284: inst = 32'hc405359;
      16285: inst = 32'h8220000;
      16286: inst = 32'h10408000;
      16287: inst = 32'hc40535a;
      16288: inst = 32'h8220000;
      16289: inst = 32'h10408000;
      16290: inst = 32'hc40535b;
      16291: inst = 32'h8220000;
      16292: inst = 32'h10408000;
      16293: inst = 32'hc40535c;
      16294: inst = 32'h8220000;
      16295: inst = 32'h10408000;
      16296: inst = 32'hc40535d;
      16297: inst = 32'h8220000;
      16298: inst = 32'h10408000;
      16299: inst = 32'hc40535e;
      16300: inst = 32'h8220000;
      16301: inst = 32'h10408000;
      16302: inst = 32'hc40535f;
      16303: inst = 32'h8220000;
      16304: inst = 32'h10408000;
      16305: inst = 32'hc405360;
      16306: inst = 32'h8220000;
      16307: inst = 32'h10408000;
      16308: inst = 32'hc405361;
      16309: inst = 32'h8220000;
      16310: inst = 32'h10408000;
      16311: inst = 32'hc405362;
      16312: inst = 32'h8220000;
      16313: inst = 32'h10408000;
      16314: inst = 32'hc405363;
      16315: inst = 32'h8220000;
      16316: inst = 32'h10408000;
      16317: inst = 32'hc405364;
      16318: inst = 32'h8220000;
      16319: inst = 32'h10408000;
      16320: inst = 32'hc405365;
      16321: inst = 32'h8220000;
      16322: inst = 32'h10408000;
      16323: inst = 32'hc405366;
      16324: inst = 32'h8220000;
      16325: inst = 32'h10408000;
      16326: inst = 32'hc405367;
      16327: inst = 32'h8220000;
      16328: inst = 32'h10408000;
      16329: inst = 32'hc405368;
      16330: inst = 32'h8220000;
      16331: inst = 32'h10408000;
      16332: inst = 32'hc405369;
      16333: inst = 32'h8220000;
      16334: inst = 32'h10408000;
      16335: inst = 32'hc40536a;
      16336: inst = 32'h8220000;
      16337: inst = 32'h10408000;
      16338: inst = 32'hc40536b;
      16339: inst = 32'h8220000;
      16340: inst = 32'h10408000;
      16341: inst = 32'hc40536c;
      16342: inst = 32'h8220000;
      16343: inst = 32'h10408000;
      16344: inst = 32'hc40536d;
      16345: inst = 32'h8220000;
      16346: inst = 32'h10408000;
      16347: inst = 32'hc40536e;
      16348: inst = 32'h8220000;
      16349: inst = 32'h10408000;
      16350: inst = 32'hc40536f;
      16351: inst = 32'h8220000;
      16352: inst = 32'h10408000;
      16353: inst = 32'hc405370;
      16354: inst = 32'h8220000;
      16355: inst = 32'h10408000;
      16356: inst = 32'hc405371;
      16357: inst = 32'h8220000;
      16358: inst = 32'h10408000;
      16359: inst = 32'hc405372;
      16360: inst = 32'h8220000;
      16361: inst = 32'h10408000;
      16362: inst = 32'hc405373;
      16363: inst = 32'h8220000;
      16364: inst = 32'h10408000;
      16365: inst = 32'hc405374;
      16366: inst = 32'h8220000;
      16367: inst = 32'h10408000;
      16368: inst = 32'hc405375;
      16369: inst = 32'h8220000;
      16370: inst = 32'h10408000;
      16371: inst = 32'hc405376;
      16372: inst = 32'h8220000;
      16373: inst = 32'h10408000;
      16374: inst = 32'hc405377;
      16375: inst = 32'h8220000;
      16376: inst = 32'h10408000;
      16377: inst = 32'hc405378;
      16378: inst = 32'h8220000;
      16379: inst = 32'h10408000;
      16380: inst = 32'hc405379;
      16381: inst = 32'h8220000;
      16382: inst = 32'h10408000;
      16383: inst = 32'hc40538a;
      16384: inst = 32'h8220000;
      16385: inst = 32'h10408000;
      16386: inst = 32'hc40538b;
      16387: inst = 32'h8220000;
      16388: inst = 32'h10408000;
      16389: inst = 32'hc40538c;
      16390: inst = 32'h8220000;
      16391: inst = 32'h10408000;
      16392: inst = 32'hc40538d;
      16393: inst = 32'h8220000;
      16394: inst = 32'h10408000;
      16395: inst = 32'hc40538e;
      16396: inst = 32'h8220000;
      16397: inst = 32'h10408000;
      16398: inst = 32'hc40538f;
      16399: inst = 32'h8220000;
      16400: inst = 32'h10408000;
      16401: inst = 32'hc405390;
      16402: inst = 32'h8220000;
      16403: inst = 32'h10408000;
      16404: inst = 32'hc405391;
      16405: inst = 32'h8220000;
      16406: inst = 32'h10408000;
      16407: inst = 32'hc405392;
      16408: inst = 32'h8220000;
      16409: inst = 32'h10408000;
      16410: inst = 32'hc405393;
      16411: inst = 32'h8220000;
      16412: inst = 32'h10408000;
      16413: inst = 32'hc405394;
      16414: inst = 32'h8220000;
      16415: inst = 32'h10408000;
      16416: inst = 32'hc405395;
      16417: inst = 32'h8220000;
      16418: inst = 32'h10408000;
      16419: inst = 32'hc4053a6;
      16420: inst = 32'h8220000;
      16421: inst = 32'h10408000;
      16422: inst = 32'hc4053a7;
      16423: inst = 32'h8220000;
      16424: inst = 32'h10408000;
      16425: inst = 32'hc4053a8;
      16426: inst = 32'h8220000;
      16427: inst = 32'h10408000;
      16428: inst = 32'hc4053a9;
      16429: inst = 32'h8220000;
      16430: inst = 32'h10408000;
      16431: inst = 32'hc4053aa;
      16432: inst = 32'h8220000;
      16433: inst = 32'h10408000;
      16434: inst = 32'hc4053ab;
      16435: inst = 32'h8220000;
      16436: inst = 32'h10408000;
      16437: inst = 32'hc4053ac;
      16438: inst = 32'h8220000;
      16439: inst = 32'h10408000;
      16440: inst = 32'hc4053ad;
      16441: inst = 32'h8220000;
      16442: inst = 32'h10408000;
      16443: inst = 32'hc4053ae;
      16444: inst = 32'h8220000;
      16445: inst = 32'h10408000;
      16446: inst = 32'hc4053af;
      16447: inst = 32'h8220000;
      16448: inst = 32'h10408000;
      16449: inst = 32'hc4053b0;
      16450: inst = 32'h8220000;
      16451: inst = 32'h10408000;
      16452: inst = 32'hc4053b1;
      16453: inst = 32'h8220000;
      16454: inst = 32'h10408000;
      16455: inst = 32'hc4053b2;
      16456: inst = 32'h8220000;
      16457: inst = 32'h10408000;
      16458: inst = 32'hc4053b3;
      16459: inst = 32'h8220000;
      16460: inst = 32'h10408000;
      16461: inst = 32'hc4053b4;
      16462: inst = 32'h8220000;
      16463: inst = 32'h10408000;
      16464: inst = 32'hc4053b5;
      16465: inst = 32'h8220000;
      16466: inst = 32'h10408000;
      16467: inst = 32'hc4053b6;
      16468: inst = 32'h8220000;
      16469: inst = 32'h10408000;
      16470: inst = 32'hc4053b7;
      16471: inst = 32'h8220000;
      16472: inst = 32'h10408000;
      16473: inst = 32'hc4053b8;
      16474: inst = 32'h8220000;
      16475: inst = 32'h10408000;
      16476: inst = 32'hc4053b9;
      16477: inst = 32'h8220000;
      16478: inst = 32'h10408000;
      16479: inst = 32'hc4053ba;
      16480: inst = 32'h8220000;
      16481: inst = 32'h10408000;
      16482: inst = 32'hc4053bb;
      16483: inst = 32'h8220000;
      16484: inst = 32'h10408000;
      16485: inst = 32'hc4053bc;
      16486: inst = 32'h8220000;
      16487: inst = 32'h10408000;
      16488: inst = 32'hc4053bd;
      16489: inst = 32'h8220000;
      16490: inst = 32'h10408000;
      16491: inst = 32'hc4053be;
      16492: inst = 32'h8220000;
      16493: inst = 32'h10408000;
      16494: inst = 32'hc4053bf;
      16495: inst = 32'h8220000;
      16496: inst = 32'h10408000;
      16497: inst = 32'hc4053c0;
      16498: inst = 32'h8220000;
      16499: inst = 32'h10408000;
      16500: inst = 32'hc4053c1;
      16501: inst = 32'h8220000;
      16502: inst = 32'h10408000;
      16503: inst = 32'hc4053c2;
      16504: inst = 32'h8220000;
      16505: inst = 32'h10408000;
      16506: inst = 32'hc4053c3;
      16507: inst = 32'h8220000;
      16508: inst = 32'h10408000;
      16509: inst = 32'hc4053c4;
      16510: inst = 32'h8220000;
      16511: inst = 32'h10408000;
      16512: inst = 32'hc4053c5;
      16513: inst = 32'h8220000;
      16514: inst = 32'h10408000;
      16515: inst = 32'hc4053c6;
      16516: inst = 32'h8220000;
      16517: inst = 32'h10408000;
      16518: inst = 32'hc4053c7;
      16519: inst = 32'h8220000;
      16520: inst = 32'h10408000;
      16521: inst = 32'hc4053c8;
      16522: inst = 32'h8220000;
      16523: inst = 32'h10408000;
      16524: inst = 32'hc4053c9;
      16525: inst = 32'h8220000;
      16526: inst = 32'h10408000;
      16527: inst = 32'hc4053ca;
      16528: inst = 32'h8220000;
      16529: inst = 32'h10408000;
      16530: inst = 32'hc4053cb;
      16531: inst = 32'h8220000;
      16532: inst = 32'h10408000;
      16533: inst = 32'hc4053cc;
      16534: inst = 32'h8220000;
      16535: inst = 32'h10408000;
      16536: inst = 32'hc4053cd;
      16537: inst = 32'h8220000;
      16538: inst = 32'h10408000;
      16539: inst = 32'hc4053ce;
      16540: inst = 32'h8220000;
      16541: inst = 32'h10408000;
      16542: inst = 32'hc4053cf;
      16543: inst = 32'h8220000;
      16544: inst = 32'h10408000;
      16545: inst = 32'hc4053d0;
      16546: inst = 32'h8220000;
      16547: inst = 32'h10408000;
      16548: inst = 32'hc4053d1;
      16549: inst = 32'h8220000;
      16550: inst = 32'h10408000;
      16551: inst = 32'hc4053d2;
      16552: inst = 32'h8220000;
      16553: inst = 32'h10408000;
      16554: inst = 32'hc4053d3;
      16555: inst = 32'h8220000;
      16556: inst = 32'h10408000;
      16557: inst = 32'hc4053d4;
      16558: inst = 32'h8220000;
      16559: inst = 32'h10408000;
      16560: inst = 32'hc4053d5;
      16561: inst = 32'h8220000;
      16562: inst = 32'h10408000;
      16563: inst = 32'hc4053d6;
      16564: inst = 32'h8220000;
      16565: inst = 32'h10408000;
      16566: inst = 32'hc4053d7;
      16567: inst = 32'h8220000;
      16568: inst = 32'h10408000;
      16569: inst = 32'hc4053d8;
      16570: inst = 32'h8220000;
      16571: inst = 32'h10408000;
      16572: inst = 32'hc4053ea;
      16573: inst = 32'h8220000;
      16574: inst = 32'h10408000;
      16575: inst = 32'hc4053eb;
      16576: inst = 32'h8220000;
      16577: inst = 32'h10408000;
      16578: inst = 32'hc4053ec;
      16579: inst = 32'h8220000;
      16580: inst = 32'h10408000;
      16581: inst = 32'hc4053ed;
      16582: inst = 32'h8220000;
      16583: inst = 32'h10408000;
      16584: inst = 32'hc4053ee;
      16585: inst = 32'h8220000;
      16586: inst = 32'h10408000;
      16587: inst = 32'hc4053ef;
      16588: inst = 32'h8220000;
      16589: inst = 32'h10408000;
      16590: inst = 32'hc4053f0;
      16591: inst = 32'h8220000;
      16592: inst = 32'h10408000;
      16593: inst = 32'hc4053f1;
      16594: inst = 32'h8220000;
      16595: inst = 32'h10408000;
      16596: inst = 32'hc4053f2;
      16597: inst = 32'h8220000;
      16598: inst = 32'h10408000;
      16599: inst = 32'hc4053f3;
      16600: inst = 32'h8220000;
      16601: inst = 32'h10408000;
      16602: inst = 32'hc4053f4;
      16603: inst = 32'h8220000;
      16604: inst = 32'h10408000;
      16605: inst = 32'hc4053f5;
      16606: inst = 32'h8220000;
      16607: inst = 32'h10408000;
      16608: inst = 32'hc405407;
      16609: inst = 32'h8220000;
      16610: inst = 32'h10408000;
      16611: inst = 32'hc405408;
      16612: inst = 32'h8220000;
      16613: inst = 32'h10408000;
      16614: inst = 32'hc405409;
      16615: inst = 32'h8220000;
      16616: inst = 32'h10408000;
      16617: inst = 32'hc40540a;
      16618: inst = 32'h8220000;
      16619: inst = 32'h10408000;
      16620: inst = 32'hc40540b;
      16621: inst = 32'h8220000;
      16622: inst = 32'h10408000;
      16623: inst = 32'hc40540c;
      16624: inst = 32'h8220000;
      16625: inst = 32'h10408000;
      16626: inst = 32'hc40540d;
      16627: inst = 32'h8220000;
      16628: inst = 32'h10408000;
      16629: inst = 32'hc40540e;
      16630: inst = 32'h8220000;
      16631: inst = 32'h10408000;
      16632: inst = 32'hc40540f;
      16633: inst = 32'h8220000;
      16634: inst = 32'h10408000;
      16635: inst = 32'hc405410;
      16636: inst = 32'h8220000;
      16637: inst = 32'h10408000;
      16638: inst = 32'hc405411;
      16639: inst = 32'h8220000;
      16640: inst = 32'h10408000;
      16641: inst = 32'hc405412;
      16642: inst = 32'h8220000;
      16643: inst = 32'h10408000;
      16644: inst = 32'hc405413;
      16645: inst = 32'h8220000;
      16646: inst = 32'h10408000;
      16647: inst = 32'hc405414;
      16648: inst = 32'h8220000;
      16649: inst = 32'h10408000;
      16650: inst = 32'hc405415;
      16651: inst = 32'h8220000;
      16652: inst = 32'h10408000;
      16653: inst = 32'hc405416;
      16654: inst = 32'h8220000;
      16655: inst = 32'h10408000;
      16656: inst = 32'hc405417;
      16657: inst = 32'h8220000;
      16658: inst = 32'h10408000;
      16659: inst = 32'hc405418;
      16660: inst = 32'h8220000;
      16661: inst = 32'h10408000;
      16662: inst = 32'hc405419;
      16663: inst = 32'h8220000;
      16664: inst = 32'h10408000;
      16665: inst = 32'hc40541a;
      16666: inst = 32'h8220000;
      16667: inst = 32'h10408000;
      16668: inst = 32'hc40541b;
      16669: inst = 32'h8220000;
      16670: inst = 32'h10408000;
      16671: inst = 32'hc40541c;
      16672: inst = 32'h8220000;
      16673: inst = 32'h10408000;
      16674: inst = 32'hc40541d;
      16675: inst = 32'h8220000;
      16676: inst = 32'h10408000;
      16677: inst = 32'hc40541e;
      16678: inst = 32'h8220000;
      16679: inst = 32'h10408000;
      16680: inst = 32'hc40541f;
      16681: inst = 32'h8220000;
      16682: inst = 32'h10408000;
      16683: inst = 32'hc405420;
      16684: inst = 32'h8220000;
      16685: inst = 32'h10408000;
      16686: inst = 32'hc405421;
      16687: inst = 32'h8220000;
      16688: inst = 32'h10408000;
      16689: inst = 32'hc405422;
      16690: inst = 32'h8220000;
      16691: inst = 32'h10408000;
      16692: inst = 32'hc405423;
      16693: inst = 32'h8220000;
      16694: inst = 32'h10408000;
      16695: inst = 32'hc405424;
      16696: inst = 32'h8220000;
      16697: inst = 32'h10408000;
      16698: inst = 32'hc405425;
      16699: inst = 32'h8220000;
      16700: inst = 32'h10408000;
      16701: inst = 32'hc405426;
      16702: inst = 32'h8220000;
      16703: inst = 32'h10408000;
      16704: inst = 32'hc405427;
      16705: inst = 32'h8220000;
      16706: inst = 32'h10408000;
      16707: inst = 32'hc405428;
      16708: inst = 32'h8220000;
      16709: inst = 32'h10408000;
      16710: inst = 32'hc405429;
      16711: inst = 32'h8220000;
      16712: inst = 32'h10408000;
      16713: inst = 32'hc40542a;
      16714: inst = 32'h8220000;
      16715: inst = 32'h10408000;
      16716: inst = 32'hc40542b;
      16717: inst = 32'h8220000;
      16718: inst = 32'h10408000;
      16719: inst = 32'hc40542c;
      16720: inst = 32'h8220000;
      16721: inst = 32'h10408000;
      16722: inst = 32'hc40542d;
      16723: inst = 32'h8220000;
      16724: inst = 32'h10408000;
      16725: inst = 32'hc40542e;
      16726: inst = 32'h8220000;
      16727: inst = 32'h10408000;
      16728: inst = 32'hc40542f;
      16729: inst = 32'h8220000;
      16730: inst = 32'h10408000;
      16731: inst = 32'hc405430;
      16732: inst = 32'h8220000;
      16733: inst = 32'h10408000;
      16734: inst = 32'hc405431;
      16735: inst = 32'h8220000;
      16736: inst = 32'h10408000;
      16737: inst = 32'hc405432;
      16738: inst = 32'h8220000;
      16739: inst = 32'h10408000;
      16740: inst = 32'hc405433;
      16741: inst = 32'h8220000;
      16742: inst = 32'h10408000;
      16743: inst = 32'hc405434;
      16744: inst = 32'h8220000;
      16745: inst = 32'h10408000;
      16746: inst = 32'hc405435;
      16747: inst = 32'h8220000;
      16748: inst = 32'h10408000;
      16749: inst = 32'hc405436;
      16750: inst = 32'h8220000;
      16751: inst = 32'h10408000;
      16752: inst = 32'hc405437;
      16753: inst = 32'h8220000;
      16754: inst = 32'h10408000;
      16755: inst = 32'hc405438;
      16756: inst = 32'h8220000;
      16757: inst = 32'h10408000;
      16758: inst = 32'hc40544a;
      16759: inst = 32'h8220000;
      16760: inst = 32'h10408000;
      16761: inst = 32'hc40544b;
      16762: inst = 32'h8220000;
      16763: inst = 32'h10408000;
      16764: inst = 32'hc40544c;
      16765: inst = 32'h8220000;
      16766: inst = 32'h10408000;
      16767: inst = 32'hc40544d;
      16768: inst = 32'h8220000;
      16769: inst = 32'h10408000;
      16770: inst = 32'hc40544e;
      16771: inst = 32'h8220000;
      16772: inst = 32'h10408000;
      16773: inst = 32'hc40544f;
      16774: inst = 32'h8220000;
      16775: inst = 32'h10408000;
      16776: inst = 32'hc405450;
      16777: inst = 32'h8220000;
      16778: inst = 32'h10408000;
      16779: inst = 32'hc405451;
      16780: inst = 32'h8220000;
      16781: inst = 32'h10408000;
      16782: inst = 32'hc405452;
      16783: inst = 32'h8220000;
      16784: inst = 32'h10408000;
      16785: inst = 32'hc405453;
      16786: inst = 32'h8220000;
      16787: inst = 32'h10408000;
      16788: inst = 32'hc405454;
      16789: inst = 32'h8220000;
      16790: inst = 32'h10408000;
      16791: inst = 32'hc405455;
      16792: inst = 32'h8220000;
      16793: inst = 32'h10408000;
      16794: inst = 32'hc405467;
      16795: inst = 32'h8220000;
      16796: inst = 32'h10408000;
      16797: inst = 32'hc405468;
      16798: inst = 32'h8220000;
      16799: inst = 32'h10408000;
      16800: inst = 32'hc405469;
      16801: inst = 32'h8220000;
      16802: inst = 32'h10408000;
      16803: inst = 32'hc40546a;
      16804: inst = 32'h8220000;
      16805: inst = 32'h10408000;
      16806: inst = 32'hc40546b;
      16807: inst = 32'h8220000;
      16808: inst = 32'h10408000;
      16809: inst = 32'hc40546c;
      16810: inst = 32'h8220000;
      16811: inst = 32'h10408000;
      16812: inst = 32'hc40546d;
      16813: inst = 32'h8220000;
      16814: inst = 32'h10408000;
      16815: inst = 32'hc40546e;
      16816: inst = 32'h8220000;
      16817: inst = 32'h10408000;
      16818: inst = 32'hc40546f;
      16819: inst = 32'h8220000;
      16820: inst = 32'h10408000;
      16821: inst = 32'hc405470;
      16822: inst = 32'h8220000;
      16823: inst = 32'h10408000;
      16824: inst = 32'hc405471;
      16825: inst = 32'h8220000;
      16826: inst = 32'h10408000;
      16827: inst = 32'hc405472;
      16828: inst = 32'h8220000;
      16829: inst = 32'h10408000;
      16830: inst = 32'hc405473;
      16831: inst = 32'h8220000;
      16832: inst = 32'h10408000;
      16833: inst = 32'hc405474;
      16834: inst = 32'h8220000;
      16835: inst = 32'h10408000;
      16836: inst = 32'hc405475;
      16837: inst = 32'h8220000;
      16838: inst = 32'h10408000;
      16839: inst = 32'hc405476;
      16840: inst = 32'h8220000;
      16841: inst = 32'h10408000;
      16842: inst = 32'hc405477;
      16843: inst = 32'h8220000;
      16844: inst = 32'h10408000;
      16845: inst = 32'hc405478;
      16846: inst = 32'h8220000;
      16847: inst = 32'h10408000;
      16848: inst = 32'hc405479;
      16849: inst = 32'h8220000;
      16850: inst = 32'h10408000;
      16851: inst = 32'hc40547a;
      16852: inst = 32'h8220000;
      16853: inst = 32'h10408000;
      16854: inst = 32'hc40547b;
      16855: inst = 32'h8220000;
      16856: inst = 32'h10408000;
      16857: inst = 32'hc40547c;
      16858: inst = 32'h8220000;
      16859: inst = 32'h10408000;
      16860: inst = 32'hc40547d;
      16861: inst = 32'h8220000;
      16862: inst = 32'h10408000;
      16863: inst = 32'hc40547e;
      16864: inst = 32'h8220000;
      16865: inst = 32'h10408000;
      16866: inst = 32'hc40547f;
      16867: inst = 32'h8220000;
      16868: inst = 32'h10408000;
      16869: inst = 32'hc405480;
      16870: inst = 32'h8220000;
      16871: inst = 32'h10408000;
      16872: inst = 32'hc405481;
      16873: inst = 32'h8220000;
      16874: inst = 32'h10408000;
      16875: inst = 32'hc405482;
      16876: inst = 32'h8220000;
      16877: inst = 32'h10408000;
      16878: inst = 32'hc405483;
      16879: inst = 32'h8220000;
      16880: inst = 32'h10408000;
      16881: inst = 32'hc405484;
      16882: inst = 32'h8220000;
      16883: inst = 32'h10408000;
      16884: inst = 32'hc405485;
      16885: inst = 32'h8220000;
      16886: inst = 32'h10408000;
      16887: inst = 32'hc405486;
      16888: inst = 32'h8220000;
      16889: inst = 32'h10408000;
      16890: inst = 32'hc405487;
      16891: inst = 32'h8220000;
      16892: inst = 32'h10408000;
      16893: inst = 32'hc405488;
      16894: inst = 32'h8220000;
      16895: inst = 32'h10408000;
      16896: inst = 32'hc405489;
      16897: inst = 32'h8220000;
      16898: inst = 32'h10408000;
      16899: inst = 32'hc40548a;
      16900: inst = 32'h8220000;
      16901: inst = 32'h10408000;
      16902: inst = 32'hc40548b;
      16903: inst = 32'h8220000;
      16904: inst = 32'h10408000;
      16905: inst = 32'hc40548c;
      16906: inst = 32'h8220000;
      16907: inst = 32'h10408000;
      16908: inst = 32'hc40548d;
      16909: inst = 32'h8220000;
      16910: inst = 32'h10408000;
      16911: inst = 32'hc40548e;
      16912: inst = 32'h8220000;
      16913: inst = 32'h10408000;
      16914: inst = 32'hc40548f;
      16915: inst = 32'h8220000;
      16916: inst = 32'h10408000;
      16917: inst = 32'hc405490;
      16918: inst = 32'h8220000;
      16919: inst = 32'h10408000;
      16920: inst = 32'hc405491;
      16921: inst = 32'h8220000;
      16922: inst = 32'h10408000;
      16923: inst = 32'hc405492;
      16924: inst = 32'h8220000;
      16925: inst = 32'h10408000;
      16926: inst = 32'hc405493;
      16927: inst = 32'h8220000;
      16928: inst = 32'h10408000;
      16929: inst = 32'hc405494;
      16930: inst = 32'h8220000;
      16931: inst = 32'h10408000;
      16932: inst = 32'hc405495;
      16933: inst = 32'h8220000;
      16934: inst = 32'h10408000;
      16935: inst = 32'hc405496;
      16936: inst = 32'h8220000;
      16937: inst = 32'h10408000;
      16938: inst = 32'hc405497;
      16939: inst = 32'h8220000;
      16940: inst = 32'h10408000;
      16941: inst = 32'hc4054aa;
      16942: inst = 32'h8220000;
      16943: inst = 32'h10408000;
      16944: inst = 32'hc4054ab;
      16945: inst = 32'h8220000;
      16946: inst = 32'h10408000;
      16947: inst = 32'hc4054ac;
      16948: inst = 32'h8220000;
      16949: inst = 32'h10408000;
      16950: inst = 32'hc4054ad;
      16951: inst = 32'h8220000;
      16952: inst = 32'h10408000;
      16953: inst = 32'hc4054ae;
      16954: inst = 32'h8220000;
      16955: inst = 32'h10408000;
      16956: inst = 32'hc4054af;
      16957: inst = 32'h8220000;
      16958: inst = 32'h10408000;
      16959: inst = 32'hc4054b0;
      16960: inst = 32'h8220000;
      16961: inst = 32'h10408000;
      16962: inst = 32'hc4054b1;
      16963: inst = 32'h8220000;
      16964: inst = 32'h10408000;
      16965: inst = 32'hc4054b2;
      16966: inst = 32'h8220000;
      16967: inst = 32'h10408000;
      16968: inst = 32'hc4054b3;
      16969: inst = 32'h8220000;
      16970: inst = 32'h10408000;
      16971: inst = 32'hc4054b4;
      16972: inst = 32'h8220000;
      16973: inst = 32'h10408000;
      16974: inst = 32'hc4054b5;
      16975: inst = 32'h8220000;
      16976: inst = 32'h10408000;
      16977: inst = 32'hc4054c8;
      16978: inst = 32'h8220000;
      16979: inst = 32'h10408000;
      16980: inst = 32'hc4054c9;
      16981: inst = 32'h8220000;
      16982: inst = 32'h10408000;
      16983: inst = 32'hc4054ca;
      16984: inst = 32'h8220000;
      16985: inst = 32'h10408000;
      16986: inst = 32'hc4054cb;
      16987: inst = 32'h8220000;
      16988: inst = 32'h10408000;
      16989: inst = 32'hc4054cc;
      16990: inst = 32'h8220000;
      16991: inst = 32'h10408000;
      16992: inst = 32'hc4054cd;
      16993: inst = 32'h8220000;
      16994: inst = 32'h10408000;
      16995: inst = 32'hc4054ce;
      16996: inst = 32'h8220000;
      16997: inst = 32'h10408000;
      16998: inst = 32'hc4054cf;
      16999: inst = 32'h8220000;
      17000: inst = 32'h10408000;
      17001: inst = 32'hc4054d0;
      17002: inst = 32'h8220000;
      17003: inst = 32'h10408000;
      17004: inst = 32'hc4054d1;
      17005: inst = 32'h8220000;
      17006: inst = 32'h10408000;
      17007: inst = 32'hc4054d2;
      17008: inst = 32'h8220000;
      17009: inst = 32'h10408000;
      17010: inst = 32'hc4054d3;
      17011: inst = 32'h8220000;
      17012: inst = 32'h10408000;
      17013: inst = 32'hc4054d4;
      17014: inst = 32'h8220000;
      17015: inst = 32'h10408000;
      17016: inst = 32'hc4054d5;
      17017: inst = 32'h8220000;
      17018: inst = 32'h10408000;
      17019: inst = 32'hc4054d6;
      17020: inst = 32'h8220000;
      17021: inst = 32'h10408000;
      17022: inst = 32'hc4054d7;
      17023: inst = 32'h8220000;
      17024: inst = 32'h10408000;
      17025: inst = 32'hc4054d8;
      17026: inst = 32'h8220000;
      17027: inst = 32'h10408000;
      17028: inst = 32'hc4054d9;
      17029: inst = 32'h8220000;
      17030: inst = 32'h10408000;
      17031: inst = 32'hc4054da;
      17032: inst = 32'h8220000;
      17033: inst = 32'h10408000;
      17034: inst = 32'hc4054db;
      17035: inst = 32'h8220000;
      17036: inst = 32'h10408000;
      17037: inst = 32'hc4054dc;
      17038: inst = 32'h8220000;
      17039: inst = 32'h10408000;
      17040: inst = 32'hc4054dd;
      17041: inst = 32'h8220000;
      17042: inst = 32'h10408000;
      17043: inst = 32'hc4054de;
      17044: inst = 32'h8220000;
      17045: inst = 32'h10408000;
      17046: inst = 32'hc4054df;
      17047: inst = 32'h8220000;
      17048: inst = 32'h10408000;
      17049: inst = 32'hc4054e0;
      17050: inst = 32'h8220000;
      17051: inst = 32'h10408000;
      17052: inst = 32'hc4054e1;
      17053: inst = 32'h8220000;
      17054: inst = 32'h10408000;
      17055: inst = 32'hc4054e2;
      17056: inst = 32'h8220000;
      17057: inst = 32'h10408000;
      17058: inst = 32'hc4054e3;
      17059: inst = 32'h8220000;
      17060: inst = 32'h10408000;
      17061: inst = 32'hc4054e4;
      17062: inst = 32'h8220000;
      17063: inst = 32'h10408000;
      17064: inst = 32'hc4054e5;
      17065: inst = 32'h8220000;
      17066: inst = 32'h10408000;
      17067: inst = 32'hc4054e6;
      17068: inst = 32'h8220000;
      17069: inst = 32'h10408000;
      17070: inst = 32'hc4054e7;
      17071: inst = 32'h8220000;
      17072: inst = 32'h10408000;
      17073: inst = 32'hc4054e8;
      17074: inst = 32'h8220000;
      17075: inst = 32'h10408000;
      17076: inst = 32'hc4054e9;
      17077: inst = 32'h8220000;
      17078: inst = 32'h10408000;
      17079: inst = 32'hc4054ea;
      17080: inst = 32'h8220000;
      17081: inst = 32'h10408000;
      17082: inst = 32'hc4054eb;
      17083: inst = 32'h8220000;
      17084: inst = 32'h10408000;
      17085: inst = 32'hc4054ec;
      17086: inst = 32'h8220000;
      17087: inst = 32'h10408000;
      17088: inst = 32'hc4054ed;
      17089: inst = 32'h8220000;
      17090: inst = 32'h10408000;
      17091: inst = 32'hc4054ee;
      17092: inst = 32'h8220000;
      17093: inst = 32'h10408000;
      17094: inst = 32'hc4054ef;
      17095: inst = 32'h8220000;
      17096: inst = 32'h10408000;
      17097: inst = 32'hc4054f0;
      17098: inst = 32'h8220000;
      17099: inst = 32'h10408000;
      17100: inst = 32'hc4054f1;
      17101: inst = 32'h8220000;
      17102: inst = 32'h10408000;
      17103: inst = 32'hc4054f2;
      17104: inst = 32'h8220000;
      17105: inst = 32'h10408000;
      17106: inst = 32'hc4054f3;
      17107: inst = 32'h8220000;
      17108: inst = 32'h10408000;
      17109: inst = 32'hc4054f4;
      17110: inst = 32'h8220000;
      17111: inst = 32'h10408000;
      17112: inst = 32'hc4054f5;
      17113: inst = 32'h8220000;
      17114: inst = 32'h10408000;
      17115: inst = 32'hc4054f6;
      17116: inst = 32'h8220000;
      17117: inst = 32'h10408000;
      17118: inst = 32'hc40550a;
      17119: inst = 32'h8220000;
      17120: inst = 32'h10408000;
      17121: inst = 32'hc40550b;
      17122: inst = 32'h8220000;
      17123: inst = 32'h10408000;
      17124: inst = 32'hc40550c;
      17125: inst = 32'h8220000;
      17126: inst = 32'h10408000;
      17127: inst = 32'hc40550d;
      17128: inst = 32'h8220000;
      17129: inst = 32'h10408000;
      17130: inst = 32'hc40550e;
      17131: inst = 32'h8220000;
      17132: inst = 32'h10408000;
      17133: inst = 32'hc40550f;
      17134: inst = 32'h8220000;
      17135: inst = 32'h10408000;
      17136: inst = 32'hc405510;
      17137: inst = 32'h8220000;
      17138: inst = 32'h10408000;
      17139: inst = 32'hc405511;
      17140: inst = 32'h8220000;
      17141: inst = 32'h10408000;
      17142: inst = 32'hc405512;
      17143: inst = 32'h8220000;
      17144: inst = 32'h10408000;
      17145: inst = 32'hc405513;
      17146: inst = 32'h8220000;
      17147: inst = 32'h10408000;
      17148: inst = 32'hc405514;
      17149: inst = 32'h8220000;
      17150: inst = 32'h10408000;
      17151: inst = 32'hc405515;
      17152: inst = 32'h8220000;
      17153: inst = 32'h10408000;
      17154: inst = 32'hc405529;
      17155: inst = 32'h8220000;
      17156: inst = 32'h10408000;
      17157: inst = 32'hc40552a;
      17158: inst = 32'h8220000;
      17159: inst = 32'h10408000;
      17160: inst = 32'hc40552b;
      17161: inst = 32'h8220000;
      17162: inst = 32'h10408000;
      17163: inst = 32'hc40552c;
      17164: inst = 32'h8220000;
      17165: inst = 32'h10408000;
      17166: inst = 32'hc40552d;
      17167: inst = 32'h8220000;
      17168: inst = 32'h10408000;
      17169: inst = 32'hc40552e;
      17170: inst = 32'h8220000;
      17171: inst = 32'h10408000;
      17172: inst = 32'hc40552f;
      17173: inst = 32'h8220000;
      17174: inst = 32'h10408000;
      17175: inst = 32'hc405530;
      17176: inst = 32'h8220000;
      17177: inst = 32'h10408000;
      17178: inst = 32'hc405531;
      17179: inst = 32'h8220000;
      17180: inst = 32'h10408000;
      17181: inst = 32'hc405532;
      17182: inst = 32'h8220000;
      17183: inst = 32'h10408000;
      17184: inst = 32'hc405533;
      17185: inst = 32'h8220000;
      17186: inst = 32'h10408000;
      17187: inst = 32'hc405534;
      17188: inst = 32'h8220000;
      17189: inst = 32'h10408000;
      17190: inst = 32'hc405535;
      17191: inst = 32'h8220000;
      17192: inst = 32'h10408000;
      17193: inst = 32'hc405536;
      17194: inst = 32'h8220000;
      17195: inst = 32'h10408000;
      17196: inst = 32'hc405537;
      17197: inst = 32'h8220000;
      17198: inst = 32'h10408000;
      17199: inst = 32'hc405538;
      17200: inst = 32'h8220000;
      17201: inst = 32'h10408000;
      17202: inst = 32'hc405539;
      17203: inst = 32'h8220000;
      17204: inst = 32'h10408000;
      17205: inst = 32'hc40553a;
      17206: inst = 32'h8220000;
      17207: inst = 32'h10408000;
      17208: inst = 32'hc40553b;
      17209: inst = 32'h8220000;
      17210: inst = 32'h10408000;
      17211: inst = 32'hc40553c;
      17212: inst = 32'h8220000;
      17213: inst = 32'h10408000;
      17214: inst = 32'hc40553d;
      17215: inst = 32'h8220000;
      17216: inst = 32'h10408000;
      17217: inst = 32'hc40553e;
      17218: inst = 32'h8220000;
      17219: inst = 32'h10408000;
      17220: inst = 32'hc40553f;
      17221: inst = 32'h8220000;
      17222: inst = 32'h10408000;
      17223: inst = 32'hc405540;
      17224: inst = 32'h8220000;
      17225: inst = 32'h10408000;
      17226: inst = 32'hc405541;
      17227: inst = 32'h8220000;
      17228: inst = 32'h10408000;
      17229: inst = 32'hc405542;
      17230: inst = 32'h8220000;
      17231: inst = 32'h10408000;
      17232: inst = 32'hc405543;
      17233: inst = 32'h8220000;
      17234: inst = 32'h10408000;
      17235: inst = 32'hc405544;
      17236: inst = 32'h8220000;
      17237: inst = 32'h10408000;
      17238: inst = 32'hc405545;
      17239: inst = 32'h8220000;
      17240: inst = 32'h10408000;
      17241: inst = 32'hc405546;
      17242: inst = 32'h8220000;
      17243: inst = 32'h10408000;
      17244: inst = 32'hc405547;
      17245: inst = 32'h8220000;
      17246: inst = 32'h10408000;
      17247: inst = 32'hc405548;
      17248: inst = 32'h8220000;
      17249: inst = 32'h10408000;
      17250: inst = 32'hc405549;
      17251: inst = 32'h8220000;
      17252: inst = 32'h10408000;
      17253: inst = 32'hc40554a;
      17254: inst = 32'h8220000;
      17255: inst = 32'h10408000;
      17256: inst = 32'hc40554b;
      17257: inst = 32'h8220000;
      17258: inst = 32'h10408000;
      17259: inst = 32'hc40554c;
      17260: inst = 32'h8220000;
      17261: inst = 32'h10408000;
      17262: inst = 32'hc40554d;
      17263: inst = 32'h8220000;
      17264: inst = 32'h10408000;
      17265: inst = 32'hc40554e;
      17266: inst = 32'h8220000;
      17267: inst = 32'h10408000;
      17268: inst = 32'hc40554f;
      17269: inst = 32'h8220000;
      17270: inst = 32'h10408000;
      17271: inst = 32'hc405550;
      17272: inst = 32'h8220000;
      17273: inst = 32'h10408000;
      17274: inst = 32'hc405551;
      17275: inst = 32'h8220000;
      17276: inst = 32'h10408000;
      17277: inst = 32'hc405552;
      17278: inst = 32'h8220000;
      17279: inst = 32'h10408000;
      17280: inst = 32'hc405553;
      17281: inst = 32'h8220000;
      17282: inst = 32'h10408000;
      17283: inst = 32'hc405554;
      17284: inst = 32'h8220000;
      17285: inst = 32'h10408000;
      17286: inst = 32'hc405555;
      17287: inst = 32'h8220000;
      17288: inst = 32'h10408000;
      17289: inst = 32'hc40556a;
      17290: inst = 32'h8220000;
      17291: inst = 32'h10408000;
      17292: inst = 32'hc40556b;
      17293: inst = 32'h8220000;
      17294: inst = 32'h10408000;
      17295: inst = 32'hc40556c;
      17296: inst = 32'h8220000;
      17297: inst = 32'h10408000;
      17298: inst = 32'hc40556d;
      17299: inst = 32'h8220000;
      17300: inst = 32'h10408000;
      17301: inst = 32'hc40556e;
      17302: inst = 32'h8220000;
      17303: inst = 32'h10408000;
      17304: inst = 32'hc40556f;
      17305: inst = 32'h8220000;
      17306: inst = 32'h10408000;
      17307: inst = 32'hc405570;
      17308: inst = 32'h8220000;
      17309: inst = 32'h10408000;
      17310: inst = 32'hc405571;
      17311: inst = 32'h8220000;
      17312: inst = 32'h10408000;
      17313: inst = 32'hc405572;
      17314: inst = 32'h8220000;
      17315: inst = 32'h10408000;
      17316: inst = 32'hc405573;
      17317: inst = 32'h8220000;
      17318: inst = 32'h10408000;
      17319: inst = 32'hc405574;
      17320: inst = 32'h8220000;
      17321: inst = 32'h10408000;
      17322: inst = 32'hc405575;
      17323: inst = 32'h8220000;
      17324: inst = 32'h10408000;
      17325: inst = 32'hc40558a;
      17326: inst = 32'h8220000;
      17327: inst = 32'h10408000;
      17328: inst = 32'hc40558b;
      17329: inst = 32'h8220000;
      17330: inst = 32'h10408000;
      17331: inst = 32'hc40558c;
      17332: inst = 32'h8220000;
      17333: inst = 32'h10408000;
      17334: inst = 32'hc40558d;
      17335: inst = 32'h8220000;
      17336: inst = 32'h10408000;
      17337: inst = 32'hc40558e;
      17338: inst = 32'h8220000;
      17339: inst = 32'h10408000;
      17340: inst = 32'hc40558f;
      17341: inst = 32'h8220000;
      17342: inst = 32'h10408000;
      17343: inst = 32'hc405590;
      17344: inst = 32'h8220000;
      17345: inst = 32'h10408000;
      17346: inst = 32'hc405591;
      17347: inst = 32'h8220000;
      17348: inst = 32'h10408000;
      17349: inst = 32'hc405592;
      17350: inst = 32'h8220000;
      17351: inst = 32'h10408000;
      17352: inst = 32'hc405593;
      17353: inst = 32'h8220000;
      17354: inst = 32'h10408000;
      17355: inst = 32'hc405594;
      17356: inst = 32'h8220000;
      17357: inst = 32'h10408000;
      17358: inst = 32'hc405595;
      17359: inst = 32'h8220000;
      17360: inst = 32'h10408000;
      17361: inst = 32'hc405596;
      17362: inst = 32'h8220000;
      17363: inst = 32'h10408000;
      17364: inst = 32'hc405597;
      17365: inst = 32'h8220000;
      17366: inst = 32'h10408000;
      17367: inst = 32'hc405598;
      17368: inst = 32'h8220000;
      17369: inst = 32'h10408000;
      17370: inst = 32'hc405599;
      17371: inst = 32'h8220000;
      17372: inst = 32'h10408000;
      17373: inst = 32'hc40559a;
      17374: inst = 32'h8220000;
      17375: inst = 32'h10408000;
      17376: inst = 32'hc40559b;
      17377: inst = 32'h8220000;
      17378: inst = 32'h10408000;
      17379: inst = 32'hc40559c;
      17380: inst = 32'h8220000;
      17381: inst = 32'h10408000;
      17382: inst = 32'hc40559d;
      17383: inst = 32'h8220000;
      17384: inst = 32'h10408000;
      17385: inst = 32'hc40559e;
      17386: inst = 32'h8220000;
      17387: inst = 32'h10408000;
      17388: inst = 32'hc40559f;
      17389: inst = 32'h8220000;
      17390: inst = 32'h10408000;
      17391: inst = 32'hc4055a0;
      17392: inst = 32'h8220000;
      17393: inst = 32'h10408000;
      17394: inst = 32'hc4055a1;
      17395: inst = 32'h8220000;
      17396: inst = 32'h10408000;
      17397: inst = 32'hc4055a2;
      17398: inst = 32'h8220000;
      17399: inst = 32'h10408000;
      17400: inst = 32'hc4055a3;
      17401: inst = 32'h8220000;
      17402: inst = 32'h10408000;
      17403: inst = 32'hc4055a4;
      17404: inst = 32'h8220000;
      17405: inst = 32'h10408000;
      17406: inst = 32'hc4055a5;
      17407: inst = 32'h8220000;
      17408: inst = 32'h10408000;
      17409: inst = 32'hc4055a6;
      17410: inst = 32'h8220000;
      17411: inst = 32'h10408000;
      17412: inst = 32'hc4055a7;
      17413: inst = 32'h8220000;
      17414: inst = 32'h10408000;
      17415: inst = 32'hc4055a8;
      17416: inst = 32'h8220000;
      17417: inst = 32'h10408000;
      17418: inst = 32'hc4055a9;
      17419: inst = 32'h8220000;
      17420: inst = 32'h10408000;
      17421: inst = 32'hc4055aa;
      17422: inst = 32'h8220000;
      17423: inst = 32'h10408000;
      17424: inst = 32'hc4055ab;
      17425: inst = 32'h8220000;
      17426: inst = 32'h10408000;
      17427: inst = 32'hc4055ac;
      17428: inst = 32'h8220000;
      17429: inst = 32'h10408000;
      17430: inst = 32'hc4055ad;
      17431: inst = 32'h8220000;
      17432: inst = 32'h10408000;
      17433: inst = 32'hc4055ae;
      17434: inst = 32'h8220000;
      17435: inst = 32'h10408000;
      17436: inst = 32'hc4055af;
      17437: inst = 32'h8220000;
      17438: inst = 32'h10408000;
      17439: inst = 32'hc4055b0;
      17440: inst = 32'h8220000;
      17441: inst = 32'h10408000;
      17442: inst = 32'hc4055b1;
      17443: inst = 32'h8220000;
      17444: inst = 32'h10408000;
      17445: inst = 32'hc4055b2;
      17446: inst = 32'h8220000;
      17447: inst = 32'h10408000;
      17448: inst = 32'hc4055b3;
      17449: inst = 32'h8220000;
      17450: inst = 32'h10408000;
      17451: inst = 32'hc4055b4;
      17452: inst = 32'h8220000;
      17453: inst = 32'h10408000;
      17454: inst = 32'hc4055ca;
      17455: inst = 32'h8220000;
      17456: inst = 32'h10408000;
      17457: inst = 32'hc4055cb;
      17458: inst = 32'h8220000;
      17459: inst = 32'h10408000;
      17460: inst = 32'hc4055cc;
      17461: inst = 32'h8220000;
      17462: inst = 32'h10408000;
      17463: inst = 32'hc4055cd;
      17464: inst = 32'h8220000;
      17465: inst = 32'h10408000;
      17466: inst = 32'hc4055ce;
      17467: inst = 32'h8220000;
      17468: inst = 32'h10408000;
      17469: inst = 32'hc4055cf;
      17470: inst = 32'h8220000;
      17471: inst = 32'h10408000;
      17472: inst = 32'hc4055d0;
      17473: inst = 32'h8220000;
      17474: inst = 32'h10408000;
      17475: inst = 32'hc4055d1;
      17476: inst = 32'h8220000;
      17477: inst = 32'h10408000;
      17478: inst = 32'hc4055d2;
      17479: inst = 32'h8220000;
      17480: inst = 32'h10408000;
      17481: inst = 32'hc4055d3;
      17482: inst = 32'h8220000;
      17483: inst = 32'h10408000;
      17484: inst = 32'hc4055d4;
      17485: inst = 32'h8220000;
      17486: inst = 32'h10408000;
      17487: inst = 32'hc4055d5;
      17488: inst = 32'h8220000;
      17489: inst = 32'h10408000;
      17490: inst = 32'hc4055eb;
      17491: inst = 32'h8220000;
      17492: inst = 32'h10408000;
      17493: inst = 32'hc4055ec;
      17494: inst = 32'h8220000;
      17495: inst = 32'h10408000;
      17496: inst = 32'hc4055ed;
      17497: inst = 32'h8220000;
      17498: inst = 32'h10408000;
      17499: inst = 32'hc4055ee;
      17500: inst = 32'h8220000;
      17501: inst = 32'h10408000;
      17502: inst = 32'hc4055ef;
      17503: inst = 32'h8220000;
      17504: inst = 32'h10408000;
      17505: inst = 32'hc4055f0;
      17506: inst = 32'h8220000;
      17507: inst = 32'h10408000;
      17508: inst = 32'hc4055f1;
      17509: inst = 32'h8220000;
      17510: inst = 32'h10408000;
      17511: inst = 32'hc4055f2;
      17512: inst = 32'h8220000;
      17513: inst = 32'h10408000;
      17514: inst = 32'hc4055f3;
      17515: inst = 32'h8220000;
      17516: inst = 32'h10408000;
      17517: inst = 32'hc4055f4;
      17518: inst = 32'h8220000;
      17519: inst = 32'h10408000;
      17520: inst = 32'hc4055f5;
      17521: inst = 32'h8220000;
      17522: inst = 32'h10408000;
      17523: inst = 32'hc4055f6;
      17524: inst = 32'h8220000;
      17525: inst = 32'h10408000;
      17526: inst = 32'hc4055f7;
      17527: inst = 32'h8220000;
      17528: inst = 32'h10408000;
      17529: inst = 32'hc4055f8;
      17530: inst = 32'h8220000;
      17531: inst = 32'h10408000;
      17532: inst = 32'hc4055f9;
      17533: inst = 32'h8220000;
      17534: inst = 32'h10408000;
      17535: inst = 32'hc4055fa;
      17536: inst = 32'h8220000;
      17537: inst = 32'h10408000;
      17538: inst = 32'hc4055fb;
      17539: inst = 32'h8220000;
      17540: inst = 32'h10408000;
      17541: inst = 32'hc4055fc;
      17542: inst = 32'h8220000;
      17543: inst = 32'h10408000;
      17544: inst = 32'hc4055fd;
      17545: inst = 32'h8220000;
      17546: inst = 32'h10408000;
      17547: inst = 32'hc4055fe;
      17548: inst = 32'h8220000;
      17549: inst = 32'h10408000;
      17550: inst = 32'hc4055ff;
      17551: inst = 32'h8220000;
      17552: inst = 32'h10408000;
      17553: inst = 32'hc405600;
      17554: inst = 32'h8220000;
      17555: inst = 32'h10408000;
      17556: inst = 32'hc405601;
      17557: inst = 32'h8220000;
      17558: inst = 32'h10408000;
      17559: inst = 32'hc405602;
      17560: inst = 32'h8220000;
      17561: inst = 32'h10408000;
      17562: inst = 32'hc405603;
      17563: inst = 32'h8220000;
      17564: inst = 32'h10408000;
      17565: inst = 32'hc405604;
      17566: inst = 32'h8220000;
      17567: inst = 32'h10408000;
      17568: inst = 32'hc405605;
      17569: inst = 32'h8220000;
      17570: inst = 32'h10408000;
      17571: inst = 32'hc405606;
      17572: inst = 32'h8220000;
      17573: inst = 32'h10408000;
      17574: inst = 32'hc405607;
      17575: inst = 32'h8220000;
      17576: inst = 32'h10408000;
      17577: inst = 32'hc405608;
      17578: inst = 32'h8220000;
      17579: inst = 32'h10408000;
      17580: inst = 32'hc405609;
      17581: inst = 32'h8220000;
      17582: inst = 32'h10408000;
      17583: inst = 32'hc40560a;
      17584: inst = 32'h8220000;
      17585: inst = 32'h10408000;
      17586: inst = 32'hc40560b;
      17587: inst = 32'h8220000;
      17588: inst = 32'h10408000;
      17589: inst = 32'hc40560c;
      17590: inst = 32'h8220000;
      17591: inst = 32'h10408000;
      17592: inst = 32'hc40560d;
      17593: inst = 32'h8220000;
      17594: inst = 32'h10408000;
      17595: inst = 32'hc40560e;
      17596: inst = 32'h8220000;
      17597: inst = 32'h10408000;
      17598: inst = 32'hc40560f;
      17599: inst = 32'h8220000;
      17600: inst = 32'h10408000;
      17601: inst = 32'hc405610;
      17602: inst = 32'h8220000;
      17603: inst = 32'h10408000;
      17604: inst = 32'hc405611;
      17605: inst = 32'h8220000;
      17606: inst = 32'h10408000;
      17607: inst = 32'hc405612;
      17608: inst = 32'h8220000;
      17609: inst = 32'h10408000;
      17610: inst = 32'hc405613;
      17611: inst = 32'h8220000;
      17612: inst = 32'h10408000;
      17613: inst = 32'hc405614;
      17614: inst = 32'h8220000;
      17615: inst = 32'h10408000;
      17616: inst = 32'hc40562a;
      17617: inst = 32'h8220000;
      17618: inst = 32'h10408000;
      17619: inst = 32'hc40562b;
      17620: inst = 32'h8220000;
      17621: inst = 32'h10408000;
      17622: inst = 32'hc40562c;
      17623: inst = 32'h8220000;
      17624: inst = 32'h10408000;
      17625: inst = 32'hc40562d;
      17626: inst = 32'h8220000;
      17627: inst = 32'h10408000;
      17628: inst = 32'hc40562e;
      17629: inst = 32'h8220000;
      17630: inst = 32'h10408000;
      17631: inst = 32'hc40562f;
      17632: inst = 32'h8220000;
      17633: inst = 32'h10408000;
      17634: inst = 32'hc405630;
      17635: inst = 32'h8220000;
      17636: inst = 32'h10408000;
      17637: inst = 32'hc405631;
      17638: inst = 32'h8220000;
      17639: inst = 32'h10408000;
      17640: inst = 32'hc405632;
      17641: inst = 32'h8220000;
      17642: inst = 32'h10408000;
      17643: inst = 32'hc405633;
      17644: inst = 32'h8220000;
      17645: inst = 32'h10408000;
      17646: inst = 32'hc405634;
      17647: inst = 32'h8220000;
      17648: inst = 32'h10408000;
      17649: inst = 32'hc405635;
      17650: inst = 32'h8220000;
      17651: inst = 32'h10408000;
      17652: inst = 32'hc40564b;
      17653: inst = 32'h8220000;
      17654: inst = 32'h10408000;
      17655: inst = 32'hc40564c;
      17656: inst = 32'h8220000;
      17657: inst = 32'h10408000;
      17658: inst = 32'hc40564d;
      17659: inst = 32'h8220000;
      17660: inst = 32'h10408000;
      17661: inst = 32'hc40564e;
      17662: inst = 32'h8220000;
      17663: inst = 32'h10408000;
      17664: inst = 32'hc40564f;
      17665: inst = 32'h8220000;
      17666: inst = 32'h10408000;
      17667: inst = 32'hc405650;
      17668: inst = 32'h8220000;
      17669: inst = 32'h10408000;
      17670: inst = 32'hc405651;
      17671: inst = 32'h8220000;
      17672: inst = 32'h10408000;
      17673: inst = 32'hc405652;
      17674: inst = 32'h8220000;
      17675: inst = 32'h10408000;
      17676: inst = 32'hc405653;
      17677: inst = 32'h8220000;
      17678: inst = 32'h10408000;
      17679: inst = 32'hc405654;
      17680: inst = 32'h8220000;
      17681: inst = 32'h10408000;
      17682: inst = 32'hc405655;
      17683: inst = 32'h8220000;
      17684: inst = 32'h10408000;
      17685: inst = 32'hc405656;
      17686: inst = 32'h8220000;
      17687: inst = 32'h10408000;
      17688: inst = 32'hc405657;
      17689: inst = 32'h8220000;
      17690: inst = 32'h10408000;
      17691: inst = 32'hc405658;
      17692: inst = 32'h8220000;
      17693: inst = 32'h10408000;
      17694: inst = 32'hc405659;
      17695: inst = 32'h8220000;
      17696: inst = 32'h10408000;
      17697: inst = 32'hc40565a;
      17698: inst = 32'h8220000;
      17699: inst = 32'h10408000;
      17700: inst = 32'hc40565b;
      17701: inst = 32'h8220000;
      17702: inst = 32'h10408000;
      17703: inst = 32'hc40565c;
      17704: inst = 32'h8220000;
      17705: inst = 32'h10408000;
      17706: inst = 32'hc40565d;
      17707: inst = 32'h8220000;
      17708: inst = 32'h10408000;
      17709: inst = 32'hc40565e;
      17710: inst = 32'h8220000;
      17711: inst = 32'h10408000;
      17712: inst = 32'hc40565f;
      17713: inst = 32'h8220000;
      17714: inst = 32'h10408000;
      17715: inst = 32'hc405660;
      17716: inst = 32'h8220000;
      17717: inst = 32'h10408000;
      17718: inst = 32'hc405661;
      17719: inst = 32'h8220000;
      17720: inst = 32'h10408000;
      17721: inst = 32'hc405662;
      17722: inst = 32'h8220000;
      17723: inst = 32'h10408000;
      17724: inst = 32'hc405663;
      17725: inst = 32'h8220000;
      17726: inst = 32'h10408000;
      17727: inst = 32'hc405664;
      17728: inst = 32'h8220000;
      17729: inst = 32'h10408000;
      17730: inst = 32'hc405665;
      17731: inst = 32'h8220000;
      17732: inst = 32'h10408000;
      17733: inst = 32'hc405666;
      17734: inst = 32'h8220000;
      17735: inst = 32'h10408000;
      17736: inst = 32'hc405667;
      17737: inst = 32'h8220000;
      17738: inst = 32'h10408000;
      17739: inst = 32'hc405668;
      17740: inst = 32'h8220000;
      17741: inst = 32'h10408000;
      17742: inst = 32'hc405669;
      17743: inst = 32'h8220000;
      17744: inst = 32'h10408000;
      17745: inst = 32'hc40566a;
      17746: inst = 32'h8220000;
      17747: inst = 32'h10408000;
      17748: inst = 32'hc40566b;
      17749: inst = 32'h8220000;
      17750: inst = 32'h10408000;
      17751: inst = 32'hc40566c;
      17752: inst = 32'h8220000;
      17753: inst = 32'h10408000;
      17754: inst = 32'hc40566d;
      17755: inst = 32'h8220000;
      17756: inst = 32'h10408000;
      17757: inst = 32'hc40566e;
      17758: inst = 32'h8220000;
      17759: inst = 32'h10408000;
      17760: inst = 32'hc40566f;
      17761: inst = 32'h8220000;
      17762: inst = 32'h10408000;
      17763: inst = 32'hc405670;
      17764: inst = 32'h8220000;
      17765: inst = 32'h10408000;
      17766: inst = 32'hc405671;
      17767: inst = 32'h8220000;
      17768: inst = 32'h10408000;
      17769: inst = 32'hc405672;
      17770: inst = 32'h8220000;
      17771: inst = 32'h10408000;
      17772: inst = 32'hc405673;
      17773: inst = 32'h8220000;
      17774: inst = 32'h10408000;
      17775: inst = 32'hc40568a;
      17776: inst = 32'h8220000;
      17777: inst = 32'h10408000;
      17778: inst = 32'hc40568b;
      17779: inst = 32'h8220000;
      17780: inst = 32'h10408000;
      17781: inst = 32'hc40568c;
      17782: inst = 32'h8220000;
      17783: inst = 32'h10408000;
      17784: inst = 32'hc40568d;
      17785: inst = 32'h8220000;
      17786: inst = 32'h10408000;
      17787: inst = 32'hc40568e;
      17788: inst = 32'h8220000;
      17789: inst = 32'h10408000;
      17790: inst = 32'hc40568f;
      17791: inst = 32'h8220000;
      17792: inst = 32'h10408000;
      17793: inst = 32'hc405690;
      17794: inst = 32'h8220000;
      17795: inst = 32'h10408000;
      17796: inst = 32'hc405691;
      17797: inst = 32'h8220000;
      17798: inst = 32'h10408000;
      17799: inst = 32'hc405692;
      17800: inst = 32'h8220000;
      17801: inst = 32'h10408000;
      17802: inst = 32'hc405693;
      17803: inst = 32'h8220000;
      17804: inst = 32'h10408000;
      17805: inst = 32'hc405694;
      17806: inst = 32'h8220000;
      17807: inst = 32'h10408000;
      17808: inst = 32'hc405695;
      17809: inst = 32'h8220000;
      17810: inst = 32'h10408000;
      17811: inst = 32'hc4056ac;
      17812: inst = 32'h8220000;
      17813: inst = 32'h10408000;
      17814: inst = 32'hc4056ad;
      17815: inst = 32'h8220000;
      17816: inst = 32'h10408000;
      17817: inst = 32'hc4056ae;
      17818: inst = 32'h8220000;
      17819: inst = 32'h10408000;
      17820: inst = 32'hc4056af;
      17821: inst = 32'h8220000;
      17822: inst = 32'h10408000;
      17823: inst = 32'hc4056b0;
      17824: inst = 32'h8220000;
      17825: inst = 32'h10408000;
      17826: inst = 32'hc4056b1;
      17827: inst = 32'h8220000;
      17828: inst = 32'h10408000;
      17829: inst = 32'hc4056b2;
      17830: inst = 32'h8220000;
      17831: inst = 32'h10408000;
      17832: inst = 32'hc4056b3;
      17833: inst = 32'h8220000;
      17834: inst = 32'h10408000;
      17835: inst = 32'hc4056b4;
      17836: inst = 32'h8220000;
      17837: inst = 32'h10408000;
      17838: inst = 32'hc4056b5;
      17839: inst = 32'h8220000;
      17840: inst = 32'h10408000;
      17841: inst = 32'hc4056b6;
      17842: inst = 32'h8220000;
      17843: inst = 32'h10408000;
      17844: inst = 32'hc4056b7;
      17845: inst = 32'h8220000;
      17846: inst = 32'h10408000;
      17847: inst = 32'hc4056b8;
      17848: inst = 32'h8220000;
      17849: inst = 32'h10408000;
      17850: inst = 32'hc4056b9;
      17851: inst = 32'h8220000;
      17852: inst = 32'h10408000;
      17853: inst = 32'hc4056ba;
      17854: inst = 32'h8220000;
      17855: inst = 32'h10408000;
      17856: inst = 32'hc4056bb;
      17857: inst = 32'h8220000;
      17858: inst = 32'h10408000;
      17859: inst = 32'hc4056bc;
      17860: inst = 32'h8220000;
      17861: inst = 32'h10408000;
      17862: inst = 32'hc4056bd;
      17863: inst = 32'h8220000;
      17864: inst = 32'h10408000;
      17865: inst = 32'hc4056be;
      17866: inst = 32'h8220000;
      17867: inst = 32'h10408000;
      17868: inst = 32'hc4056bf;
      17869: inst = 32'h8220000;
      17870: inst = 32'h10408000;
      17871: inst = 32'hc4056c0;
      17872: inst = 32'h8220000;
      17873: inst = 32'h10408000;
      17874: inst = 32'hc4056c1;
      17875: inst = 32'h8220000;
      17876: inst = 32'h10408000;
      17877: inst = 32'hc4056c2;
      17878: inst = 32'h8220000;
      17879: inst = 32'h10408000;
      17880: inst = 32'hc4056c3;
      17881: inst = 32'h8220000;
      17882: inst = 32'h10408000;
      17883: inst = 32'hc4056c4;
      17884: inst = 32'h8220000;
      17885: inst = 32'h10408000;
      17886: inst = 32'hc4056c5;
      17887: inst = 32'h8220000;
      17888: inst = 32'h10408000;
      17889: inst = 32'hc4056c6;
      17890: inst = 32'h8220000;
      17891: inst = 32'h10408000;
      17892: inst = 32'hc4056c7;
      17893: inst = 32'h8220000;
      17894: inst = 32'h10408000;
      17895: inst = 32'hc4056c8;
      17896: inst = 32'h8220000;
      17897: inst = 32'h10408000;
      17898: inst = 32'hc4056c9;
      17899: inst = 32'h8220000;
      17900: inst = 32'h10408000;
      17901: inst = 32'hc4056ca;
      17902: inst = 32'h8220000;
      17903: inst = 32'h10408000;
      17904: inst = 32'hc4056cb;
      17905: inst = 32'h8220000;
      17906: inst = 32'h10408000;
      17907: inst = 32'hc4056cc;
      17908: inst = 32'h8220000;
      17909: inst = 32'h10408000;
      17910: inst = 32'hc4056cd;
      17911: inst = 32'h8220000;
      17912: inst = 32'h10408000;
      17913: inst = 32'hc4056ce;
      17914: inst = 32'h8220000;
      17915: inst = 32'h10408000;
      17916: inst = 32'hc4056cf;
      17917: inst = 32'h8220000;
      17918: inst = 32'h10408000;
      17919: inst = 32'hc4056d0;
      17920: inst = 32'h8220000;
      17921: inst = 32'h10408000;
      17922: inst = 32'hc4056d1;
      17923: inst = 32'h8220000;
      17924: inst = 32'h10408000;
      17925: inst = 32'hc4056d2;
      17926: inst = 32'h8220000;
      17927: inst = 32'h10408000;
      17928: inst = 32'hc4056ea;
      17929: inst = 32'h8220000;
      17930: inst = 32'h10408000;
      17931: inst = 32'hc4056eb;
      17932: inst = 32'h8220000;
      17933: inst = 32'h10408000;
      17934: inst = 32'hc4056ec;
      17935: inst = 32'h8220000;
      17936: inst = 32'h10408000;
      17937: inst = 32'hc4056ed;
      17938: inst = 32'h8220000;
      17939: inst = 32'h10408000;
      17940: inst = 32'hc4056ee;
      17941: inst = 32'h8220000;
      17942: inst = 32'h10408000;
      17943: inst = 32'hc4056ef;
      17944: inst = 32'h8220000;
      17945: inst = 32'h10408000;
      17946: inst = 32'hc4056f0;
      17947: inst = 32'h8220000;
      17948: inst = 32'h10408000;
      17949: inst = 32'hc4056f1;
      17950: inst = 32'h8220000;
      17951: inst = 32'h10408000;
      17952: inst = 32'hc4056f2;
      17953: inst = 32'h8220000;
      17954: inst = 32'h10408000;
      17955: inst = 32'hc4056f3;
      17956: inst = 32'h8220000;
      17957: inst = 32'h10408000;
      17958: inst = 32'hc4056f4;
      17959: inst = 32'h8220000;
      17960: inst = 32'h10408000;
      17961: inst = 32'hc4056f5;
      17962: inst = 32'h8220000;
      17963: inst = 32'h10408000;
      17964: inst = 32'hc40570d;
      17965: inst = 32'h8220000;
      17966: inst = 32'h10408000;
      17967: inst = 32'hc40570e;
      17968: inst = 32'h8220000;
      17969: inst = 32'h10408000;
      17970: inst = 32'hc40570f;
      17971: inst = 32'h8220000;
      17972: inst = 32'h10408000;
      17973: inst = 32'hc405710;
      17974: inst = 32'h8220000;
      17975: inst = 32'h10408000;
      17976: inst = 32'hc405711;
      17977: inst = 32'h8220000;
      17978: inst = 32'h10408000;
      17979: inst = 32'hc405712;
      17980: inst = 32'h8220000;
      17981: inst = 32'h10408000;
      17982: inst = 32'hc405713;
      17983: inst = 32'h8220000;
      17984: inst = 32'h10408000;
      17985: inst = 32'hc405714;
      17986: inst = 32'h8220000;
      17987: inst = 32'h10408000;
      17988: inst = 32'hc405715;
      17989: inst = 32'h8220000;
      17990: inst = 32'h10408000;
      17991: inst = 32'hc405716;
      17992: inst = 32'h8220000;
      17993: inst = 32'h10408000;
      17994: inst = 32'hc405717;
      17995: inst = 32'h8220000;
      17996: inst = 32'h10408000;
      17997: inst = 32'hc405718;
      17998: inst = 32'h8220000;
      17999: inst = 32'h10408000;
      18000: inst = 32'hc405719;
      18001: inst = 32'h8220000;
      18002: inst = 32'h10408000;
      18003: inst = 32'hc40571a;
      18004: inst = 32'h8220000;
      18005: inst = 32'h10408000;
      18006: inst = 32'hc40571b;
      18007: inst = 32'h8220000;
      18008: inst = 32'h10408000;
      18009: inst = 32'hc40571c;
      18010: inst = 32'h8220000;
      18011: inst = 32'h10408000;
      18012: inst = 32'hc40571d;
      18013: inst = 32'h8220000;
      18014: inst = 32'h10408000;
      18015: inst = 32'hc40571e;
      18016: inst = 32'h8220000;
      18017: inst = 32'h10408000;
      18018: inst = 32'hc40571f;
      18019: inst = 32'h8220000;
      18020: inst = 32'h10408000;
      18021: inst = 32'hc405720;
      18022: inst = 32'h8220000;
      18023: inst = 32'h10408000;
      18024: inst = 32'hc405721;
      18025: inst = 32'h8220000;
      18026: inst = 32'h10408000;
      18027: inst = 32'hc405722;
      18028: inst = 32'h8220000;
      18029: inst = 32'h10408000;
      18030: inst = 32'hc405723;
      18031: inst = 32'h8220000;
      18032: inst = 32'h10408000;
      18033: inst = 32'hc405724;
      18034: inst = 32'h8220000;
      18035: inst = 32'h10408000;
      18036: inst = 32'hc405725;
      18037: inst = 32'h8220000;
      18038: inst = 32'h10408000;
      18039: inst = 32'hc405726;
      18040: inst = 32'h8220000;
      18041: inst = 32'h10408000;
      18042: inst = 32'hc405727;
      18043: inst = 32'h8220000;
      18044: inst = 32'h10408000;
      18045: inst = 32'hc405728;
      18046: inst = 32'h8220000;
      18047: inst = 32'h10408000;
      18048: inst = 32'hc405729;
      18049: inst = 32'h8220000;
      18050: inst = 32'h10408000;
      18051: inst = 32'hc40572a;
      18052: inst = 32'h8220000;
      18053: inst = 32'h10408000;
      18054: inst = 32'hc40572b;
      18055: inst = 32'h8220000;
      18056: inst = 32'h10408000;
      18057: inst = 32'hc40572c;
      18058: inst = 32'h8220000;
      18059: inst = 32'h10408000;
      18060: inst = 32'hc40572d;
      18061: inst = 32'h8220000;
      18062: inst = 32'h10408000;
      18063: inst = 32'hc40572e;
      18064: inst = 32'h8220000;
      18065: inst = 32'h10408000;
      18066: inst = 32'hc40572f;
      18067: inst = 32'h8220000;
      18068: inst = 32'h10408000;
      18069: inst = 32'hc405730;
      18070: inst = 32'h8220000;
      18071: inst = 32'h10408000;
      18072: inst = 32'hc405731;
      18073: inst = 32'h8220000;
      18074: inst = 32'h10408000;
      18075: inst = 32'hc40574a;
      18076: inst = 32'h8220000;
      18077: inst = 32'h10408000;
      18078: inst = 32'hc40574b;
      18079: inst = 32'h8220000;
      18080: inst = 32'h10408000;
      18081: inst = 32'hc40574c;
      18082: inst = 32'h8220000;
      18083: inst = 32'h10408000;
      18084: inst = 32'hc40574d;
      18085: inst = 32'h8220000;
      18086: inst = 32'h10408000;
      18087: inst = 32'hc40574e;
      18088: inst = 32'h8220000;
      18089: inst = 32'h10408000;
      18090: inst = 32'hc40574f;
      18091: inst = 32'h8220000;
      18092: inst = 32'h10408000;
      18093: inst = 32'hc405750;
      18094: inst = 32'h8220000;
      18095: inst = 32'h10408000;
      18096: inst = 32'hc405751;
      18097: inst = 32'h8220000;
      18098: inst = 32'h10408000;
      18099: inst = 32'hc405752;
      18100: inst = 32'h8220000;
      18101: inst = 32'h10408000;
      18102: inst = 32'hc405753;
      18103: inst = 32'h8220000;
      18104: inst = 32'h10408000;
      18105: inst = 32'hc405754;
      18106: inst = 32'h8220000;
      18107: inst = 32'h10408000;
      18108: inst = 32'hc405755;
      18109: inst = 32'h8220000;
      18110: inst = 32'h10408000;
      18111: inst = 32'hc40576e;
      18112: inst = 32'h8220000;
      18113: inst = 32'h10408000;
      18114: inst = 32'hc40576f;
      18115: inst = 32'h8220000;
      18116: inst = 32'h10408000;
      18117: inst = 32'hc405770;
      18118: inst = 32'h8220000;
      18119: inst = 32'h10408000;
      18120: inst = 32'hc405771;
      18121: inst = 32'h8220000;
      18122: inst = 32'h10408000;
      18123: inst = 32'hc405772;
      18124: inst = 32'h8220000;
      18125: inst = 32'h10408000;
      18126: inst = 32'hc405773;
      18127: inst = 32'h8220000;
      18128: inst = 32'h10408000;
      18129: inst = 32'hc405774;
      18130: inst = 32'h8220000;
      18131: inst = 32'h10408000;
      18132: inst = 32'hc405775;
      18133: inst = 32'h8220000;
      18134: inst = 32'h10408000;
      18135: inst = 32'hc405776;
      18136: inst = 32'h8220000;
      18137: inst = 32'h10408000;
      18138: inst = 32'hc405777;
      18139: inst = 32'h8220000;
      18140: inst = 32'h10408000;
      18141: inst = 32'hc405778;
      18142: inst = 32'h8220000;
      18143: inst = 32'h10408000;
      18144: inst = 32'hc405779;
      18145: inst = 32'h8220000;
      18146: inst = 32'h10408000;
      18147: inst = 32'hc40577a;
      18148: inst = 32'h8220000;
      18149: inst = 32'h10408000;
      18150: inst = 32'hc40577b;
      18151: inst = 32'h8220000;
      18152: inst = 32'h10408000;
      18153: inst = 32'hc40577c;
      18154: inst = 32'h8220000;
      18155: inst = 32'h10408000;
      18156: inst = 32'hc40577d;
      18157: inst = 32'h8220000;
      18158: inst = 32'h10408000;
      18159: inst = 32'hc40577e;
      18160: inst = 32'h8220000;
      18161: inst = 32'h10408000;
      18162: inst = 32'hc40577f;
      18163: inst = 32'h8220000;
      18164: inst = 32'h10408000;
      18165: inst = 32'hc405780;
      18166: inst = 32'h8220000;
      18167: inst = 32'h10408000;
      18168: inst = 32'hc405781;
      18169: inst = 32'h8220000;
      18170: inst = 32'h10408000;
      18171: inst = 32'hc405782;
      18172: inst = 32'h8220000;
      18173: inst = 32'h10408000;
      18174: inst = 32'hc405783;
      18175: inst = 32'h8220000;
      18176: inst = 32'h10408000;
      18177: inst = 32'hc405784;
      18178: inst = 32'h8220000;
      18179: inst = 32'h10408000;
      18180: inst = 32'hc405785;
      18181: inst = 32'h8220000;
      18182: inst = 32'h10408000;
      18183: inst = 32'hc405786;
      18184: inst = 32'h8220000;
      18185: inst = 32'h10408000;
      18186: inst = 32'hc405787;
      18187: inst = 32'h8220000;
      18188: inst = 32'h10408000;
      18189: inst = 32'hc405788;
      18190: inst = 32'h8220000;
      18191: inst = 32'h10408000;
      18192: inst = 32'hc405789;
      18193: inst = 32'h8220000;
      18194: inst = 32'h10408000;
      18195: inst = 32'hc40578a;
      18196: inst = 32'h8220000;
      18197: inst = 32'h10408000;
      18198: inst = 32'hc40578b;
      18199: inst = 32'h8220000;
      18200: inst = 32'h10408000;
      18201: inst = 32'hc40578c;
      18202: inst = 32'h8220000;
      18203: inst = 32'h10408000;
      18204: inst = 32'hc40578d;
      18205: inst = 32'h8220000;
      18206: inst = 32'h10408000;
      18207: inst = 32'hc40578e;
      18208: inst = 32'h8220000;
      18209: inst = 32'h10408000;
      18210: inst = 32'hc40578f;
      18211: inst = 32'h8220000;
      18212: inst = 32'h10408000;
      18213: inst = 32'hc405790;
      18214: inst = 32'h8220000;
      18215: inst = 32'h10408000;
      18216: inst = 32'hc405791;
      18217: inst = 32'h8220000;
      18218: inst = 32'h10408000;
      18219: inst = 32'hc4057aa;
      18220: inst = 32'h8220000;
      18221: inst = 32'h10408000;
      18222: inst = 32'hc4057ab;
      18223: inst = 32'h8220000;
      18224: inst = 32'h10408000;
      18225: inst = 32'hc4057ac;
      18226: inst = 32'h8220000;
      18227: inst = 32'h10408000;
      18228: inst = 32'hc4057ad;
      18229: inst = 32'h8220000;
      18230: inst = 32'h10408000;
      18231: inst = 32'hc4057ae;
      18232: inst = 32'h8220000;
      18233: inst = 32'h10408000;
      18234: inst = 32'hc4057af;
      18235: inst = 32'h8220000;
      18236: inst = 32'h10408000;
      18237: inst = 32'hc4057b0;
      18238: inst = 32'h8220000;
      18239: inst = 32'h10408000;
      18240: inst = 32'hc4057b1;
      18241: inst = 32'h8220000;
      18242: inst = 32'h10408000;
      18243: inst = 32'hc4057b2;
      18244: inst = 32'h8220000;
      18245: inst = 32'h10408000;
      18246: inst = 32'hc4057b3;
      18247: inst = 32'h8220000;
      18248: inst = 32'h10408000;
      18249: inst = 32'hc4057b4;
      18250: inst = 32'h8220000;
      18251: inst = 32'h10408000;
      18252: inst = 32'hc4057b5;
      18253: inst = 32'h8220000;
      18254: inst = 32'h10408000;
      18255: inst = 32'hc4057ce;
      18256: inst = 32'h8220000;
      18257: inst = 32'h10408000;
      18258: inst = 32'hc4057cf;
      18259: inst = 32'h8220000;
      18260: inst = 32'h10408000;
      18261: inst = 32'hc4057d0;
      18262: inst = 32'h8220000;
      18263: inst = 32'h10408000;
      18264: inst = 32'hc4057d1;
      18265: inst = 32'h8220000;
      18266: inst = 32'h10408000;
      18267: inst = 32'hc4057d2;
      18268: inst = 32'h8220000;
      18269: inst = 32'h10408000;
      18270: inst = 32'hc4057d3;
      18271: inst = 32'h8220000;
      18272: inst = 32'h10408000;
      18273: inst = 32'hc4057d4;
      18274: inst = 32'h8220000;
      18275: inst = 32'h10408000;
      18276: inst = 32'hc4057d5;
      18277: inst = 32'h8220000;
      18278: inst = 32'h10408000;
      18279: inst = 32'hc4057d6;
      18280: inst = 32'h8220000;
      18281: inst = 32'h10408000;
      18282: inst = 32'hc4057d7;
      18283: inst = 32'h8220000;
      18284: inst = 32'h10408000;
      18285: inst = 32'hc4057d8;
      18286: inst = 32'h8220000;
      18287: inst = 32'h10408000;
      18288: inst = 32'hc4057d9;
      18289: inst = 32'h8220000;
      18290: inst = 32'h10408000;
      18291: inst = 32'hc4057da;
      18292: inst = 32'h8220000;
      18293: inst = 32'h10408000;
      18294: inst = 32'hc4057db;
      18295: inst = 32'h8220000;
      18296: inst = 32'h10408000;
      18297: inst = 32'hc4057dc;
      18298: inst = 32'h8220000;
      18299: inst = 32'h10408000;
      18300: inst = 32'hc4057dd;
      18301: inst = 32'h8220000;
      18302: inst = 32'h10408000;
      18303: inst = 32'hc4057de;
      18304: inst = 32'h8220000;
      18305: inst = 32'h10408000;
      18306: inst = 32'hc4057df;
      18307: inst = 32'h8220000;
      18308: inst = 32'hc207bd0;
      18309: inst = 32'h10408000;
      18310: inst = 32'hc40531b;
      18311: inst = 32'h8220000;
      18312: inst = 32'h10408000;
      18313: inst = 32'hc405344;
      18314: inst = 32'h8220000;
      18315: inst = 32'hc207bcf;
      18316: inst = 32'h10408000;
      18317: inst = 32'hc405321;
      18318: inst = 32'h8220000;
      18319: inst = 32'h10408000;
      18320: inst = 32'hc40533e;
      18321: inst = 32'h8220000;
      18322: inst = 32'h10408000;
      18323: inst = 32'hc405381;
      18324: inst = 32'h8220000;
      18325: inst = 32'h10408000;
      18326: inst = 32'hc40539e;
      18327: inst = 32'h8220000;
      18328: inst = 32'h10408000;
      18329: inst = 32'hc4053e1;
      18330: inst = 32'h8220000;
      18331: inst = 32'h10408000;
      18332: inst = 32'hc4053fe;
      18333: inst = 32'h8220000;
      18334: inst = 32'h10408000;
      18335: inst = 32'hc405441;
      18336: inst = 32'h8220000;
      18337: inst = 32'h10408000;
      18338: inst = 32'hc405448;
      18339: inst = 32'h8220000;
      18340: inst = 32'h10408000;
      18341: inst = 32'hc405457;
      18342: inst = 32'h8220000;
      18343: inst = 32'h10408000;
      18344: inst = 32'hc40545e;
      18345: inst = 32'h8220000;
      18346: inst = 32'h10408000;
      18347: inst = 32'hc405501;
      18348: inst = 32'h8220000;
      18349: inst = 32'h10408000;
      18350: inst = 32'hc40551e;
      18351: inst = 32'h8220000;
      18352: inst = 32'h10408000;
      18353: inst = 32'hc405561;
      18354: inst = 32'h8220000;
      18355: inst = 32'h10408000;
      18356: inst = 32'hc40557e;
      18357: inst = 32'h8220000;
      18358: inst = 32'h10408000;
      18359: inst = 32'hc4055b9;
      18360: inst = 32'h8220000;
      18361: inst = 32'h10408000;
      18362: inst = 32'hc4055c1;
      18363: inst = 32'h8220000;
      18364: inst = 32'h10408000;
      18365: inst = 32'hc4055de;
      18366: inst = 32'h8220000;
      18367: inst = 32'h10408000;
      18368: inst = 32'hc4055e6;
      18369: inst = 32'h8220000;
      18370: inst = 32'h10408000;
      18371: inst = 32'hc40561e;
      18372: inst = 32'h8220000;
      18373: inst = 32'h10408000;
      18374: inst = 32'hc405621;
      18375: inst = 32'h8220000;
      18376: inst = 32'h10408000;
      18377: inst = 32'hc40563e;
      18378: inst = 32'h8220000;
      18379: inst = 32'h10408000;
      18380: inst = 32'hc405641;
      18381: inst = 32'h8220000;
      18382: inst = 32'h10408000;
      18383: inst = 32'hc405681;
      18384: inst = 32'h8220000;
      18385: inst = 32'h10408000;
      18386: inst = 32'hc405698;
      18387: inst = 32'h8220000;
      18388: inst = 32'h10408000;
      18389: inst = 32'hc40569e;
      18390: inst = 32'h8220000;
      18391: inst = 32'h10408000;
      18392: inst = 32'hc4056e1;
      18393: inst = 32'h8220000;
      18394: inst = 32'h10408000;
      18395: inst = 32'hc4056fe;
      18396: inst = 32'h8220000;
      18397: inst = 32'hc207390;
      18398: inst = 32'h10408000;
      18399: inst = 32'hc40537a;
      18400: inst = 32'h8220000;
      18401: inst = 32'h10408000;
      18402: inst = 32'hc4053a5;
      18403: inst = 32'h8220000;
      18404: inst = 32'hc2052aa;
      18405: inst = 32'h10408000;
      18406: inst = 32'hc405389;
      18407: inst = 32'h8220000;
      18408: inst = 32'h10408000;
      18409: inst = 32'hc405396;
      18410: inst = 32'h8220000;
      18411: inst = 32'h10408000;
      18412: inst = 32'hc4054fb;
      18413: inst = 32'h8220000;
      18414: inst = 32'h10408000;
      18415: inst = 32'hc405503;
      18416: inst = 32'h8220000;
      18417: inst = 32'h10408000;
      18418: inst = 32'hc40551c;
      18419: inst = 32'h8220000;
      18420: inst = 32'h10408000;
      18421: inst = 32'hc405524;
      18422: inst = 32'h8220000;
      18423: inst = 32'h10408000;
      18424: inst = 32'hc4055c8;
      18425: inst = 32'h8220000;
      18426: inst = 32'h10408000;
      18427: inst = 32'hc4055d7;
      18428: inst = 32'h8220000;
      18429: inst = 32'h10408000;
      18430: inst = 32'hc405619;
      18431: inst = 32'h8220000;
      18432: inst = 32'h10408000;
      18433: inst = 32'hc405622;
      18434: inst = 32'h8220000;
      18435: inst = 32'h10408000;
      18436: inst = 32'hc40563d;
      18437: inst = 32'h8220000;
      18438: inst = 32'h10408000;
      18439: inst = 32'hc405646;
      18440: inst = 32'h8220000;
      18441: inst = 32'hc206b70;
      18442: inst = 32'h10408000;
      18443: inst = 32'hc4053d9;
      18444: inst = 32'h8220000;
      18445: inst = 32'h10408000;
      18446: inst = 32'hc405406;
      18447: inst = 32'h8220000;
      18448: inst = 32'h10408000;
      18449: inst = 32'hc405556;
      18450: inst = 32'h8220000;
      18451: inst = 32'h10408000;
      18452: inst = 32'hc405589;
      18453: inst = 32'h8220000;
      18454: inst = 32'h10408000;
      18455: inst = 32'hc4055b5;
      18456: inst = 32'h8220000;
      18457: inst = 32'h10408000;
      18458: inst = 32'hc4055ea;
      18459: inst = 32'h8220000;
      18460: inst = 32'h10408000;
      18461: inst = 32'hc405732;
      18462: inst = 32'h8220000;
      18463: inst = 32'h10408000;
      18464: inst = 32'hc40576d;
      18465: inst = 32'h8220000;
      18466: inst = 32'hc20736e;
      18467: inst = 32'h10408000;
      18468: inst = 32'hc4053e0;
      18469: inst = 32'h8220000;
      18470: inst = 32'h10408000;
      18471: inst = 32'hc4053ff;
      18472: inst = 32'h8220000;
      18473: inst = 32'hc205aaa;
      18474: inst = 32'h10408000;
      18475: inst = 32'hc4053e4;
      18476: inst = 32'h8220000;
      18477: inst = 32'h10408000;
      18478: inst = 32'hc4053fb;
      18479: inst = 32'h8220000;
      18480: inst = 32'hc208431;
      18481: inst = 32'h10408000;
      18482: inst = 32'hc4053e8;
      18483: inst = 32'h8220000;
      18484: inst = 32'h10408000;
      18485: inst = 32'hc4053f7;
      18486: inst = 32'h8220000;
      18487: inst = 32'h10408000;
      18488: inst = 32'hc405439;
      18489: inst = 32'h8220000;
      18490: inst = 32'h10408000;
      18491: inst = 32'hc405466;
      18492: inst = 32'h8220000;
      18493: inst = 32'h10408000;
      18494: inst = 32'hc4055b6;
      18495: inst = 32'h8220000;
      18496: inst = 32'h10408000;
      18497: inst = 32'hc4055e9;
      18498: inst = 32'h8220000;
      18499: inst = 32'h10408000;
      18500: inst = 32'hc405733;
      18501: inst = 32'h8220000;
      18502: inst = 32'h10408000;
      18503: inst = 32'hc40576c;
      18504: inst = 32'h8220000;
      18505: inst = 32'hc206b4d;
      18506: inst = 32'h10408000;
      18507: inst = 32'hc40543c;
      18508: inst = 32'h8220000;
      18509: inst = 32'h10408000;
      18510: inst = 32'hc405444;
      18511: inst = 32'h8220000;
      18512: inst = 32'h10408000;
      18513: inst = 32'hc40545b;
      18514: inst = 32'h8220000;
      18515: inst = 32'h10408000;
      18516: inst = 32'hc405463;
      18517: inst = 32'h8220000;
      18518: inst = 32'h10408000;
      18519: inst = 32'hc405563;
      18520: inst = 32'h8220000;
      18521: inst = 32'h10408000;
      18522: inst = 32'hc40557c;
      18523: inst = 32'h8220000;
      18524: inst = 32'h10408000;
      18525: inst = 32'hc405682;
      18526: inst = 32'h8220000;
      18527: inst = 32'h10408000;
      18528: inst = 32'hc40569d;
      18529: inst = 32'h8220000;
      18530: inst = 32'hc208430;
      18531: inst = 32'h10408000;
      18532: inst = 32'hc405440;
      18533: inst = 32'h8220000;
      18534: inst = 32'h10408000;
      18535: inst = 32'hc40545f;
      18536: inst = 32'h8220000;
      18537: inst = 32'hc207bf1;
      18538: inst = 32'h10408000;
      18539: inst = 32'hc405498;
      18540: inst = 32'h8220000;
      18541: inst = 32'h10408000;
      18542: inst = 32'hc4054c7;
      18543: inst = 32'h8220000;
      18544: inst = 32'h10408000;
      18545: inst = 32'hc405615;
      18546: inst = 32'h8220000;
      18547: inst = 32'h10408000;
      18548: inst = 32'hc40564a;
      18549: inst = 32'h8220000;
      18550: inst = 32'hc207bef;
      18551: inst = 32'h10408000;
      18552: inst = 32'hc40549b;
      18553: inst = 32'h8220000;
      18554: inst = 32'h10408000;
      18555: inst = 32'hc4054c4;
      18556: inst = 32'h8220000;
      18557: inst = 32'h10408000;
      18558: inst = 32'hc405687;
      18559: inst = 32'h8220000;
      18560: inst = 32'h10408000;
      18561: inst = 32'hc4056e2;
      18562: inst = 32'h8220000;
      18563: inst = 32'h10408000;
      18564: inst = 32'hc4056fd;
      18565: inst = 32'h8220000;
      18566: inst = 32'hc205aeb;
      18567: inst = 32'h10408000;
      18568: inst = 32'hc40549f;
      18569: inst = 32'h8220000;
      18570: inst = 32'h10408000;
      18571: inst = 32'hc4054c0;
      18572: inst = 32'h8220000;
      18573: inst = 32'hc206b6e;
      18574: inst = 32'h10408000;
      18575: inst = 32'hc4054a8;
      18576: inst = 32'h8220000;
      18577: inst = 32'h10408000;
      18578: inst = 32'hc4054b7;
      18579: inst = 32'h8220000;
      18580: inst = 32'h10408000;
      18581: inst = 32'hc4056e7;
      18582: inst = 32'h8220000;
      18583: inst = 32'h10408000;
      18584: inst = 32'hc4056f8;
      18585: inst = 32'h8220000;
      18586: inst = 32'hc2073b0;
      18587: inst = 32'h10408000;
      18588: inst = 32'hc4054f7;
      18589: inst = 32'h8220000;
      18590: inst = 32'h10408000;
      18591: inst = 32'hc405528;
      18592: inst = 32'h8220000;
      18593: inst = 32'h10408000;
      18594: inst = 32'hc405674;
      18595: inst = 32'h8220000;
      18596: inst = 32'h10408000;
      18597: inst = 32'hc4056ab;
      18598: inst = 32'h8220000;
      18599: inst = 32'hc2073ae;
      18600: inst = 32'h10408000;
      18601: inst = 32'hc4054ff;
      18602: inst = 32'h8220000;
      18603: inst = 32'h10408000;
      18604: inst = 32'hc405520;
      18605: inst = 32'h8220000;
      18606: inst = 32'hc20632d;
      18607: inst = 32'h10408000;
      18608: inst = 32'hc405508;
      18609: inst = 32'h8220000;
      18610: inst = 32'h10408000;
      18611: inst = 32'hc405517;
      18612: inst = 32'h8220000;
      18613: inst = 32'h10408000;
      18614: inst = 32'hc405747;
      18615: inst = 32'h8220000;
      18616: inst = 32'h10408000;
      18617: inst = 32'hc405758;
      18618: inst = 32'h8220000;
      18619: inst = 32'hc206b2d;
      18620: inst = 32'h10408000;
      18621: inst = 32'hc40555a;
      18622: inst = 32'h8220000;
      18623: inst = 32'h10408000;
      18624: inst = 32'hc405585;
      18625: inst = 32'h8220000;
      18626: inst = 32'hc20630c;
      18627: inst = 32'h10408000;
      18628: inst = 32'hc4055be;
      18629: inst = 32'h8220000;
      18630: inst = 32'h10408000;
      18631: inst = 32'hc4055e1;
      18632: inst = 32'h8220000;
      18633: inst = 32'h10408000;
      18634: inst = 32'hc405678;
      18635: inst = 32'h8220000;
      18636: inst = 32'hc20632c;
      18637: inst = 32'h10408000;
      18638: inst = 32'hc4056a7;
      18639: inst = 32'h8220000;
      18640: inst = 32'hc206b90;
      18641: inst = 32'h10408000;
      18642: inst = 32'hc4056d3;
      18643: inst = 32'h8220000;
      18644: inst = 32'h10408000;
      18645: inst = 32'hc40570c;
      18646: inst = 32'h8220000;
      18647: inst = 32'hc207c11;
      18648: inst = 32'h10408000;
      18649: inst = 32'hc405792;
      18650: inst = 32'h8220000;
      18651: inst = 32'h10408000;
      18652: inst = 32'hc4057cd;
      18653: inst = 32'h8220000;
      18654: inst = 32'h58000000;
      18655: inst = 32'hc20ea25;
      18656: inst = 32'h10408000;
      18657: inst = 32'hc40464d;
      18658: inst = 32'h8220000;
      18659: inst = 32'h10408000;
      18660: inst = 32'hc40464e;
      18661: inst = 32'h8220000;
      18662: inst = 32'h10408000;
      18663: inst = 32'hc40464f;
      18664: inst = 32'h8220000;
      18665: inst = 32'h10408000;
      18666: inst = 32'hc404650;
      18667: inst = 32'h8220000;
      18668: inst = 32'h10408000;
      18669: inst = 32'hc404651;
      18670: inst = 32'h8220000;
      18671: inst = 32'h10408000;
      18672: inst = 32'hc404652;
      18673: inst = 32'h8220000;
      18674: inst = 32'h10408000;
      18675: inst = 32'hc404653;
      18676: inst = 32'h8220000;
      18677: inst = 32'h10408000;
      18678: inst = 32'hc404654;
      18679: inst = 32'h8220000;
      18680: inst = 32'h10408000;
      18681: inst = 32'hc404655;
      18682: inst = 32'h8220000;
      18683: inst = 32'h10408000;
      18684: inst = 32'hc404659;
      18685: inst = 32'h8220000;
      18686: inst = 32'h10408000;
      18687: inst = 32'hc40465a;
      18688: inst = 32'h8220000;
      18689: inst = 32'h10408000;
      18690: inst = 32'hc40465b;
      18691: inst = 32'h8220000;
      18692: inst = 32'h10408000;
      18693: inst = 32'hc40465c;
      18694: inst = 32'h8220000;
      18695: inst = 32'h10408000;
      18696: inst = 32'hc40465d;
      18697: inst = 32'h8220000;
      18698: inst = 32'h10408000;
      18699: inst = 32'hc40465e;
      18700: inst = 32'h8220000;
      18701: inst = 32'h10408000;
      18702: inst = 32'hc40465f;
      18703: inst = 32'h8220000;
      18704: inst = 32'h10408000;
      18705: inst = 32'hc404660;
      18706: inst = 32'h8220000;
      18707: inst = 32'h10408000;
      18708: inst = 32'hc404661;
      18709: inst = 32'h8220000;
      18710: inst = 32'h10408000;
      18711: inst = 32'hc404663;
      18712: inst = 32'h8220000;
      18713: inst = 32'h10408000;
      18714: inst = 32'hc404664;
      18715: inst = 32'h8220000;
      18716: inst = 32'h10408000;
      18717: inst = 32'hc404665;
      18718: inst = 32'h8220000;
      18719: inst = 32'h10408000;
      18720: inst = 32'hc404666;
      18721: inst = 32'h8220000;
      18722: inst = 32'h10408000;
      18723: inst = 32'hc404667;
      18724: inst = 32'h8220000;
      18725: inst = 32'h10408000;
      18726: inst = 32'hc404668;
      18727: inst = 32'h8220000;
      18728: inst = 32'h10408000;
      18729: inst = 32'hc404669;
      18730: inst = 32'h8220000;
      18731: inst = 32'h10408000;
      18732: inst = 32'hc40466a;
      18733: inst = 32'h8220000;
      18734: inst = 32'h10408000;
      18735: inst = 32'hc40466b;
      18736: inst = 32'h8220000;
      18737: inst = 32'h10408000;
      18738: inst = 32'hc404671;
      18739: inst = 32'h8220000;
      18740: inst = 32'h10408000;
      18741: inst = 32'hc404672;
      18742: inst = 32'h8220000;
      18743: inst = 32'h10408000;
      18744: inst = 32'hc404673;
      18745: inst = 32'h8220000;
      18746: inst = 32'h10408000;
      18747: inst = 32'hc404674;
      18748: inst = 32'h8220000;
      18749: inst = 32'h10408000;
      18750: inst = 32'hc404675;
      18751: inst = 32'h8220000;
      18752: inst = 32'h10408000;
      18753: inst = 32'hc404676;
      18754: inst = 32'h8220000;
      18755: inst = 32'h10408000;
      18756: inst = 32'hc404677;
      18757: inst = 32'h8220000;
      18758: inst = 32'h10408000;
      18759: inst = 32'hc404678;
      18760: inst = 32'h8220000;
      18761: inst = 32'h10408000;
      18762: inst = 32'hc404679;
      18763: inst = 32'h8220000;
      18764: inst = 32'h10408000;
      18765: inst = 32'hc40467c;
      18766: inst = 32'h8220000;
      18767: inst = 32'h10408000;
      18768: inst = 32'hc40467d;
      18769: inst = 32'h8220000;
      18770: inst = 32'h10408000;
      18771: inst = 32'hc40467e;
      18772: inst = 32'h8220000;
      18773: inst = 32'h10408000;
      18774: inst = 32'hc40467f;
      18775: inst = 32'h8220000;
      18776: inst = 32'h10408000;
      18777: inst = 32'hc404680;
      18778: inst = 32'h8220000;
      18779: inst = 32'h10408000;
      18780: inst = 32'hc404681;
      18781: inst = 32'h8220000;
      18782: inst = 32'h10408000;
      18783: inst = 32'hc404682;
      18784: inst = 32'h8220000;
      18785: inst = 32'h10408000;
      18786: inst = 32'hc404683;
      18787: inst = 32'h8220000;
      18788: inst = 32'h10408000;
      18789: inst = 32'hc404684;
      18790: inst = 32'h8220000;
      18791: inst = 32'h10408000;
      18792: inst = 32'hc404685;
      18793: inst = 32'h8220000;
      18794: inst = 32'h10408000;
      18795: inst = 32'hc40468b;
      18796: inst = 32'h8220000;
      18797: inst = 32'h10408000;
      18798: inst = 32'hc40468c;
      18799: inst = 32'h8220000;
      18800: inst = 32'h10408000;
      18801: inst = 32'hc40468d;
      18802: inst = 32'h8220000;
      18803: inst = 32'h10408000;
      18804: inst = 32'hc40468e;
      18805: inst = 32'h8220000;
      18806: inst = 32'h10408000;
      18807: inst = 32'hc40468f;
      18808: inst = 32'h8220000;
      18809: inst = 32'h10408000;
      18810: inst = 32'hc404690;
      18811: inst = 32'h8220000;
      18812: inst = 32'h10408000;
      18813: inst = 32'hc404691;
      18814: inst = 32'h8220000;
      18815: inst = 32'h10408000;
      18816: inst = 32'hc404692;
      18817: inst = 32'h8220000;
      18818: inst = 32'h10408000;
      18819: inst = 32'hc404693;
      18820: inst = 32'h8220000;
      18821: inst = 32'h10408000;
      18822: inst = 32'hc4046ac;
      18823: inst = 32'h8220000;
      18824: inst = 32'h10408000;
      18825: inst = 32'hc4046ad;
      18826: inst = 32'h8220000;
      18827: inst = 32'h10408000;
      18828: inst = 32'hc4046ae;
      18829: inst = 32'h8220000;
      18830: inst = 32'h10408000;
      18831: inst = 32'hc4046af;
      18832: inst = 32'h8220000;
      18833: inst = 32'h10408000;
      18834: inst = 32'hc4046b0;
      18835: inst = 32'h8220000;
      18836: inst = 32'h10408000;
      18837: inst = 32'hc4046b1;
      18838: inst = 32'h8220000;
      18839: inst = 32'h10408000;
      18840: inst = 32'hc4046b2;
      18841: inst = 32'h8220000;
      18842: inst = 32'h10408000;
      18843: inst = 32'hc4046b3;
      18844: inst = 32'h8220000;
      18845: inst = 32'h10408000;
      18846: inst = 32'hc4046b4;
      18847: inst = 32'h8220000;
      18848: inst = 32'h10408000;
      18849: inst = 32'hc4046b5;
      18850: inst = 32'h8220000;
      18851: inst = 32'h10408000;
      18852: inst = 32'hc4046b8;
      18853: inst = 32'h8220000;
      18854: inst = 32'h10408000;
      18855: inst = 32'hc4046b9;
      18856: inst = 32'h8220000;
      18857: inst = 32'h10408000;
      18858: inst = 32'hc4046ba;
      18859: inst = 32'h8220000;
      18860: inst = 32'h10408000;
      18861: inst = 32'hc4046bb;
      18862: inst = 32'h8220000;
      18863: inst = 32'h10408000;
      18864: inst = 32'hc4046bc;
      18865: inst = 32'h8220000;
      18866: inst = 32'h10408000;
      18867: inst = 32'hc4046bd;
      18868: inst = 32'h8220000;
      18869: inst = 32'h10408000;
      18870: inst = 32'hc4046be;
      18871: inst = 32'h8220000;
      18872: inst = 32'h10408000;
      18873: inst = 32'hc4046bf;
      18874: inst = 32'h8220000;
      18875: inst = 32'h10408000;
      18876: inst = 32'hc4046c0;
      18877: inst = 32'h8220000;
      18878: inst = 32'h10408000;
      18879: inst = 32'hc4046c1;
      18880: inst = 32'h8220000;
      18881: inst = 32'h10408000;
      18882: inst = 32'hc4046c3;
      18883: inst = 32'h8220000;
      18884: inst = 32'h10408000;
      18885: inst = 32'hc4046c4;
      18886: inst = 32'h8220000;
      18887: inst = 32'h10408000;
      18888: inst = 32'hc4046c5;
      18889: inst = 32'h8220000;
      18890: inst = 32'h10408000;
      18891: inst = 32'hc4046c6;
      18892: inst = 32'h8220000;
      18893: inst = 32'h10408000;
      18894: inst = 32'hc4046c7;
      18895: inst = 32'h8220000;
      18896: inst = 32'h10408000;
      18897: inst = 32'hc4046c8;
      18898: inst = 32'h8220000;
      18899: inst = 32'h10408000;
      18900: inst = 32'hc4046c9;
      18901: inst = 32'h8220000;
      18902: inst = 32'h10408000;
      18903: inst = 32'hc4046ca;
      18904: inst = 32'h8220000;
      18905: inst = 32'h10408000;
      18906: inst = 32'hc4046cb;
      18907: inst = 32'h8220000;
      18908: inst = 32'h10408000;
      18909: inst = 32'hc4046d0;
      18910: inst = 32'h8220000;
      18911: inst = 32'h10408000;
      18912: inst = 32'hc4046d1;
      18913: inst = 32'h8220000;
      18914: inst = 32'h10408000;
      18915: inst = 32'hc4046d2;
      18916: inst = 32'h8220000;
      18917: inst = 32'h10408000;
      18918: inst = 32'hc4046d3;
      18919: inst = 32'h8220000;
      18920: inst = 32'h10408000;
      18921: inst = 32'hc4046d4;
      18922: inst = 32'h8220000;
      18923: inst = 32'h10408000;
      18924: inst = 32'hc4046d5;
      18925: inst = 32'h8220000;
      18926: inst = 32'h10408000;
      18927: inst = 32'hc4046d6;
      18928: inst = 32'h8220000;
      18929: inst = 32'h10408000;
      18930: inst = 32'hc4046d7;
      18931: inst = 32'h8220000;
      18932: inst = 32'h10408000;
      18933: inst = 32'hc4046d8;
      18934: inst = 32'h8220000;
      18935: inst = 32'h10408000;
      18936: inst = 32'hc4046da;
      18937: inst = 32'h8220000;
      18938: inst = 32'h10408000;
      18939: inst = 32'hc4046dc;
      18940: inst = 32'h8220000;
      18941: inst = 32'h10408000;
      18942: inst = 32'hc4046dd;
      18943: inst = 32'h8220000;
      18944: inst = 32'h10408000;
      18945: inst = 32'hc4046de;
      18946: inst = 32'h8220000;
      18947: inst = 32'h10408000;
      18948: inst = 32'hc4046df;
      18949: inst = 32'h8220000;
      18950: inst = 32'h10408000;
      18951: inst = 32'hc4046e0;
      18952: inst = 32'h8220000;
      18953: inst = 32'h10408000;
      18954: inst = 32'hc4046e1;
      18955: inst = 32'h8220000;
      18956: inst = 32'h10408000;
      18957: inst = 32'hc4046e2;
      18958: inst = 32'h8220000;
      18959: inst = 32'h10408000;
      18960: inst = 32'hc4046e3;
      18961: inst = 32'h8220000;
      18962: inst = 32'h10408000;
      18963: inst = 32'hc4046e4;
      18964: inst = 32'h8220000;
      18965: inst = 32'h10408000;
      18966: inst = 32'hc4046e5;
      18967: inst = 32'h8220000;
      18968: inst = 32'h10408000;
      18969: inst = 32'hc4046ea;
      18970: inst = 32'h8220000;
      18971: inst = 32'h10408000;
      18972: inst = 32'hc4046eb;
      18973: inst = 32'h8220000;
      18974: inst = 32'h10408000;
      18975: inst = 32'hc4046ec;
      18976: inst = 32'h8220000;
      18977: inst = 32'h10408000;
      18978: inst = 32'hc4046ed;
      18979: inst = 32'h8220000;
      18980: inst = 32'h10408000;
      18981: inst = 32'hc4046ee;
      18982: inst = 32'h8220000;
      18983: inst = 32'h10408000;
      18984: inst = 32'hc4046ef;
      18985: inst = 32'h8220000;
      18986: inst = 32'h10408000;
      18987: inst = 32'hc4046f0;
      18988: inst = 32'h8220000;
      18989: inst = 32'h10408000;
      18990: inst = 32'hc4046f1;
      18991: inst = 32'h8220000;
      18992: inst = 32'h10408000;
      18993: inst = 32'hc4046f2;
      18994: inst = 32'h8220000;
      18995: inst = 32'h10408000;
      18996: inst = 32'hc4046f3;
      18997: inst = 32'h8220000;
      18998: inst = 32'h10408000;
      18999: inst = 32'hc40470b;
      19000: inst = 32'h8220000;
      19001: inst = 32'h10408000;
      19002: inst = 32'hc40470c;
      19003: inst = 32'h8220000;
      19004: inst = 32'h10408000;
      19005: inst = 32'hc40470d;
      19006: inst = 32'h8220000;
      19007: inst = 32'h10408000;
      19008: inst = 32'hc404717;
      19009: inst = 32'h8220000;
      19010: inst = 32'h10408000;
      19011: inst = 32'hc404718;
      19012: inst = 32'h8220000;
      19013: inst = 32'h10408000;
      19014: inst = 32'hc404719;
      19015: inst = 32'h8220000;
      19016: inst = 32'h10408000;
      19017: inst = 32'hc404728;
      19018: inst = 32'h8220000;
      19019: inst = 32'h10408000;
      19020: inst = 32'hc404729;
      19021: inst = 32'h8220000;
      19022: inst = 32'h10408000;
      19023: inst = 32'hc40472a;
      19024: inst = 32'h8220000;
      19025: inst = 32'h10408000;
      19026: inst = 32'hc40472b;
      19027: inst = 32'h8220000;
      19028: inst = 32'h10408000;
      19029: inst = 32'hc404730;
      19030: inst = 32'h8220000;
      19031: inst = 32'h10408000;
      19032: inst = 32'hc404731;
      19033: inst = 32'h8220000;
      19034: inst = 32'h10408000;
      19035: inst = 32'hc404735;
      19036: inst = 32'h8220000;
      19037: inst = 32'h10408000;
      19038: inst = 32'hc404736;
      19039: inst = 32'h8220000;
      19040: inst = 32'h10408000;
      19041: inst = 32'hc404737;
      19042: inst = 32'h8220000;
      19043: inst = 32'h10408000;
      19044: inst = 32'hc404739;
      19045: inst = 32'h8220000;
      19046: inst = 32'h10408000;
      19047: inst = 32'hc40473a;
      19048: inst = 32'h8220000;
      19049: inst = 32'h10408000;
      19050: inst = 32'hc404742;
      19051: inst = 32'h8220000;
      19052: inst = 32'h10408000;
      19053: inst = 32'hc404743;
      19054: inst = 32'h8220000;
      19055: inst = 32'h10408000;
      19056: inst = 32'hc404744;
      19057: inst = 32'h8220000;
      19058: inst = 32'h10408000;
      19059: inst = 32'hc404745;
      19060: inst = 32'h8220000;
      19061: inst = 32'h10408000;
      19062: inst = 32'hc404749;
      19063: inst = 32'h8220000;
      19064: inst = 32'h10408000;
      19065: inst = 32'hc40474a;
      19066: inst = 32'h8220000;
      19067: inst = 32'h10408000;
      19068: inst = 32'hc40474b;
      19069: inst = 32'h8220000;
      19070: inst = 32'h10408000;
      19071: inst = 32'hc40476b;
      19072: inst = 32'h8220000;
      19073: inst = 32'h10408000;
      19074: inst = 32'hc40476c;
      19075: inst = 32'h8220000;
      19076: inst = 32'h10408000;
      19077: inst = 32'hc404777;
      19078: inst = 32'h8220000;
      19079: inst = 32'h10408000;
      19080: inst = 32'hc404778;
      19081: inst = 32'h8220000;
      19082: inst = 32'h10408000;
      19083: inst = 32'hc404788;
      19084: inst = 32'h8220000;
      19085: inst = 32'h10408000;
      19086: inst = 32'hc404789;
      19087: inst = 32'h8220000;
      19088: inst = 32'h10408000;
      19089: inst = 32'hc40478a;
      19090: inst = 32'h8220000;
      19091: inst = 32'h10408000;
      19092: inst = 32'hc404790;
      19093: inst = 32'h8220000;
      19094: inst = 32'h10408000;
      19095: inst = 32'hc404791;
      19096: inst = 32'h8220000;
      19097: inst = 32'h10408000;
      19098: inst = 32'hc404795;
      19099: inst = 32'h8220000;
      19100: inst = 32'h10408000;
      19101: inst = 32'hc404799;
      19102: inst = 32'h8220000;
      19103: inst = 32'h10408000;
      19104: inst = 32'hc40479a;
      19105: inst = 32'h8220000;
      19106: inst = 32'h10408000;
      19107: inst = 32'hc4047a2;
      19108: inst = 32'h8220000;
      19109: inst = 32'h10408000;
      19110: inst = 32'hc4047a3;
      19111: inst = 32'h8220000;
      19112: inst = 32'h10408000;
      19113: inst = 32'hc4047a4;
      19114: inst = 32'h8220000;
      19115: inst = 32'h10408000;
      19116: inst = 32'hc4047a9;
      19117: inst = 32'h8220000;
      19118: inst = 32'h10408000;
      19119: inst = 32'hc4047aa;
      19120: inst = 32'h8220000;
      19121: inst = 32'h10408000;
      19122: inst = 32'hc4047cb;
      19123: inst = 32'h8220000;
      19124: inst = 32'h10408000;
      19125: inst = 32'hc4047cc;
      19126: inst = 32'h8220000;
      19127: inst = 32'h10408000;
      19128: inst = 32'hc4047ce;
      19129: inst = 32'h8220000;
      19130: inst = 32'h10408000;
      19131: inst = 32'hc4047cf;
      19132: inst = 32'h8220000;
      19133: inst = 32'h10408000;
      19134: inst = 32'hc4047d0;
      19135: inst = 32'h8220000;
      19136: inst = 32'h10408000;
      19137: inst = 32'hc4047d1;
      19138: inst = 32'h8220000;
      19139: inst = 32'h10408000;
      19140: inst = 32'hc4047d2;
      19141: inst = 32'h8220000;
      19142: inst = 32'h10408000;
      19143: inst = 32'hc4047d7;
      19144: inst = 32'h8220000;
      19145: inst = 32'h10408000;
      19146: inst = 32'hc4047d8;
      19147: inst = 32'h8220000;
      19148: inst = 32'h10408000;
      19149: inst = 32'hc4047da;
      19150: inst = 32'h8220000;
      19151: inst = 32'h10408000;
      19152: inst = 32'hc4047db;
      19153: inst = 32'h8220000;
      19154: inst = 32'h10408000;
      19155: inst = 32'hc4047dc;
      19156: inst = 32'h8220000;
      19157: inst = 32'h10408000;
      19158: inst = 32'hc4047dd;
      19159: inst = 32'h8220000;
      19160: inst = 32'h10408000;
      19161: inst = 32'hc4047de;
      19162: inst = 32'h8220000;
      19163: inst = 32'h10408000;
      19164: inst = 32'hc4047e7;
      19165: inst = 32'h8220000;
      19166: inst = 32'h10408000;
      19167: inst = 32'hc4047e8;
      19168: inst = 32'h8220000;
      19169: inst = 32'h10408000;
      19170: inst = 32'hc4047e9;
      19171: inst = 32'h8220000;
      19172: inst = 32'h10408000;
      19173: inst = 32'hc4047f0;
      19174: inst = 32'h8220000;
      19175: inst = 32'h10408000;
      19176: inst = 32'hc4047f1;
      19177: inst = 32'h8220000;
      19178: inst = 32'h10408000;
      19179: inst = 32'hc4047f9;
      19180: inst = 32'h8220000;
      19181: inst = 32'h10408000;
      19182: inst = 32'hc4047fa;
      19183: inst = 32'h8220000;
      19184: inst = 32'h10408000;
      19185: inst = 32'hc404800;
      19186: inst = 32'h8220000;
      19187: inst = 32'h10408000;
      19188: inst = 32'hc404801;
      19189: inst = 32'h8220000;
      19190: inst = 32'h10408000;
      19191: inst = 32'hc404802;
      19192: inst = 32'h8220000;
      19193: inst = 32'h10408000;
      19194: inst = 32'hc404803;
      19195: inst = 32'h8220000;
      19196: inst = 32'h10408000;
      19197: inst = 32'hc404809;
      19198: inst = 32'h8220000;
      19199: inst = 32'h10408000;
      19200: inst = 32'hc40480a;
      19201: inst = 32'h8220000;
      19202: inst = 32'h10408000;
      19203: inst = 32'hc40480c;
      19204: inst = 32'h8220000;
      19205: inst = 32'h10408000;
      19206: inst = 32'hc40480d;
      19207: inst = 32'h8220000;
      19208: inst = 32'h10408000;
      19209: inst = 32'hc40480e;
      19210: inst = 32'h8220000;
      19211: inst = 32'h10408000;
      19212: inst = 32'hc40480f;
      19213: inst = 32'h8220000;
      19214: inst = 32'h10408000;
      19215: inst = 32'hc404810;
      19216: inst = 32'h8220000;
      19217: inst = 32'h10408000;
      19218: inst = 32'hc404811;
      19219: inst = 32'h8220000;
      19220: inst = 32'h10408000;
      19221: inst = 32'hc40482b;
      19222: inst = 32'h8220000;
      19223: inst = 32'h10408000;
      19224: inst = 32'hc40482c;
      19225: inst = 32'h8220000;
      19226: inst = 32'h10408000;
      19227: inst = 32'hc40482e;
      19228: inst = 32'h8220000;
      19229: inst = 32'h10408000;
      19230: inst = 32'hc40482f;
      19231: inst = 32'h8220000;
      19232: inst = 32'h10408000;
      19233: inst = 32'hc404830;
      19234: inst = 32'h8220000;
      19235: inst = 32'h10408000;
      19236: inst = 32'hc404831;
      19237: inst = 32'h8220000;
      19238: inst = 32'h10408000;
      19239: inst = 32'hc404832;
      19240: inst = 32'h8220000;
      19241: inst = 32'h10408000;
      19242: inst = 32'hc404837;
      19243: inst = 32'h8220000;
      19244: inst = 32'h10408000;
      19245: inst = 32'hc404838;
      19246: inst = 32'h8220000;
      19247: inst = 32'h10408000;
      19248: inst = 32'hc40483a;
      19249: inst = 32'h8220000;
      19250: inst = 32'h10408000;
      19251: inst = 32'hc40483b;
      19252: inst = 32'h8220000;
      19253: inst = 32'h10408000;
      19254: inst = 32'hc40483c;
      19255: inst = 32'h8220000;
      19256: inst = 32'h10408000;
      19257: inst = 32'hc40483d;
      19258: inst = 32'h8220000;
      19259: inst = 32'h10408000;
      19260: inst = 32'hc40483e;
      19261: inst = 32'h8220000;
      19262: inst = 32'h10408000;
      19263: inst = 32'hc404846;
      19264: inst = 32'h8220000;
      19265: inst = 32'h10408000;
      19266: inst = 32'hc404847;
      19267: inst = 32'h8220000;
      19268: inst = 32'h10408000;
      19269: inst = 32'hc404848;
      19270: inst = 32'h8220000;
      19271: inst = 32'h10408000;
      19272: inst = 32'hc404850;
      19273: inst = 32'h8220000;
      19274: inst = 32'h10408000;
      19275: inst = 32'hc404851;
      19276: inst = 32'h8220000;
      19277: inst = 32'h10408000;
      19278: inst = 32'hc404859;
      19279: inst = 32'h8220000;
      19280: inst = 32'h10408000;
      19281: inst = 32'hc40485a;
      19282: inst = 32'h8220000;
      19283: inst = 32'h10408000;
      19284: inst = 32'hc40485f;
      19285: inst = 32'h8220000;
      19286: inst = 32'h10408000;
      19287: inst = 32'hc404860;
      19288: inst = 32'h8220000;
      19289: inst = 32'h10408000;
      19290: inst = 32'hc404861;
      19291: inst = 32'h8220000;
      19292: inst = 32'h10408000;
      19293: inst = 32'hc404862;
      19294: inst = 32'h8220000;
      19295: inst = 32'h10408000;
      19296: inst = 32'hc404869;
      19297: inst = 32'h8220000;
      19298: inst = 32'h10408000;
      19299: inst = 32'hc40486a;
      19300: inst = 32'h8220000;
      19301: inst = 32'h10408000;
      19302: inst = 32'hc40486c;
      19303: inst = 32'h8220000;
      19304: inst = 32'h10408000;
      19305: inst = 32'hc40486d;
      19306: inst = 32'h8220000;
      19307: inst = 32'h10408000;
      19308: inst = 32'hc40486e;
      19309: inst = 32'h8220000;
      19310: inst = 32'h10408000;
      19311: inst = 32'hc40486f;
      19312: inst = 32'h8220000;
      19313: inst = 32'h10408000;
      19314: inst = 32'hc404870;
      19315: inst = 32'h8220000;
      19316: inst = 32'h10408000;
      19317: inst = 32'hc404871;
      19318: inst = 32'h8220000;
      19319: inst = 32'h10408000;
      19320: inst = 32'hc404872;
      19321: inst = 32'h8220000;
      19322: inst = 32'h10408000;
      19323: inst = 32'hc40488b;
      19324: inst = 32'h8220000;
      19325: inst = 32'h10408000;
      19326: inst = 32'hc40488c;
      19327: inst = 32'h8220000;
      19328: inst = 32'h10408000;
      19329: inst = 32'hc404897;
      19330: inst = 32'h8220000;
      19331: inst = 32'h10408000;
      19332: inst = 32'hc404898;
      19333: inst = 32'h8220000;
      19334: inst = 32'h10408000;
      19335: inst = 32'hc4048a6;
      19336: inst = 32'h8220000;
      19337: inst = 32'h10408000;
      19338: inst = 32'hc4048b0;
      19339: inst = 32'h8220000;
      19340: inst = 32'h10408000;
      19341: inst = 32'hc4048b1;
      19342: inst = 32'h8220000;
      19343: inst = 32'h10408000;
      19344: inst = 32'hc4048b4;
      19345: inst = 32'h8220000;
      19346: inst = 32'h10408000;
      19347: inst = 32'hc4048b5;
      19348: inst = 32'h8220000;
      19349: inst = 32'h10408000;
      19350: inst = 32'hc4048b9;
      19351: inst = 32'h8220000;
      19352: inst = 32'h10408000;
      19353: inst = 32'hc4048ba;
      19354: inst = 32'h8220000;
      19355: inst = 32'h10408000;
      19356: inst = 32'hc4048bf;
      19357: inst = 32'h8220000;
      19358: inst = 32'h10408000;
      19359: inst = 32'hc4048c9;
      19360: inst = 32'h8220000;
      19361: inst = 32'h10408000;
      19362: inst = 32'hc4048ca;
      19363: inst = 32'h8220000;
      19364: inst = 32'h10408000;
      19365: inst = 32'hc4048d1;
      19366: inst = 32'h8220000;
      19367: inst = 32'h10408000;
      19368: inst = 32'hc4048d2;
      19369: inst = 32'h8220000;
      19370: inst = 32'h10408000;
      19371: inst = 32'hc4048d3;
      19372: inst = 32'h8220000;
      19373: inst = 32'h10408000;
      19374: inst = 32'hc4048eb;
      19375: inst = 32'h8220000;
      19376: inst = 32'h10408000;
      19377: inst = 32'hc4048ec;
      19378: inst = 32'h8220000;
      19379: inst = 32'h10408000;
      19380: inst = 32'hc4048ed;
      19381: inst = 32'h8220000;
      19382: inst = 32'h10408000;
      19383: inst = 32'hc4048ee;
      19384: inst = 32'h8220000;
      19385: inst = 32'h10408000;
      19386: inst = 32'hc4048ef;
      19387: inst = 32'h8220000;
      19388: inst = 32'h10408000;
      19389: inst = 32'hc4048f0;
      19390: inst = 32'h8220000;
      19391: inst = 32'h10408000;
      19392: inst = 32'hc4048f1;
      19393: inst = 32'h8220000;
      19394: inst = 32'h10408000;
      19395: inst = 32'hc4048f2;
      19396: inst = 32'h8220000;
      19397: inst = 32'h10408000;
      19398: inst = 32'hc4048f3;
      19399: inst = 32'h8220000;
      19400: inst = 32'h10408000;
      19401: inst = 32'hc4048f4;
      19402: inst = 32'h8220000;
      19403: inst = 32'h10408000;
      19404: inst = 32'hc4048f5;
      19405: inst = 32'h8220000;
      19406: inst = 32'h10408000;
      19407: inst = 32'hc4048f7;
      19408: inst = 32'h8220000;
      19409: inst = 32'h10408000;
      19410: inst = 32'hc4048f8;
      19411: inst = 32'h8220000;
      19412: inst = 32'h10408000;
      19413: inst = 32'hc4048f9;
      19414: inst = 32'h8220000;
      19415: inst = 32'h10408000;
      19416: inst = 32'hc4048fa;
      19417: inst = 32'h8220000;
      19418: inst = 32'h10408000;
      19419: inst = 32'hc4048fb;
      19420: inst = 32'h8220000;
      19421: inst = 32'h10408000;
      19422: inst = 32'hc4048fc;
      19423: inst = 32'h8220000;
      19424: inst = 32'h10408000;
      19425: inst = 32'hc4048fd;
      19426: inst = 32'h8220000;
      19427: inst = 32'h10408000;
      19428: inst = 32'hc4048fe;
      19429: inst = 32'h8220000;
      19430: inst = 32'h10408000;
      19431: inst = 32'hc4048ff;
      19432: inst = 32'h8220000;
      19433: inst = 32'h10408000;
      19434: inst = 32'hc404900;
      19435: inst = 32'h8220000;
      19436: inst = 32'h10408000;
      19437: inst = 32'hc404901;
      19438: inst = 32'h8220000;
      19439: inst = 32'h10408000;
      19440: inst = 32'hc404904;
      19441: inst = 32'h8220000;
      19442: inst = 32'h10408000;
      19443: inst = 32'hc404905;
      19444: inst = 32'h8220000;
      19445: inst = 32'h10408000;
      19446: inst = 32'hc404906;
      19447: inst = 32'h8220000;
      19448: inst = 32'h10408000;
      19449: inst = 32'hc404907;
      19450: inst = 32'h8220000;
      19451: inst = 32'h10408000;
      19452: inst = 32'hc404908;
      19453: inst = 32'h8220000;
      19454: inst = 32'h10408000;
      19455: inst = 32'hc404909;
      19456: inst = 32'h8220000;
      19457: inst = 32'h10408000;
      19458: inst = 32'hc40490a;
      19459: inst = 32'h8220000;
      19460: inst = 32'h10408000;
      19461: inst = 32'hc40490b;
      19462: inst = 32'h8220000;
      19463: inst = 32'h10408000;
      19464: inst = 32'hc40490c;
      19465: inst = 32'h8220000;
      19466: inst = 32'h10408000;
      19467: inst = 32'hc40490d;
      19468: inst = 32'h8220000;
      19469: inst = 32'h10408000;
      19470: inst = 32'hc404910;
      19471: inst = 32'h8220000;
      19472: inst = 32'h10408000;
      19473: inst = 32'hc404911;
      19474: inst = 32'h8220000;
      19475: inst = 32'h10408000;
      19476: inst = 32'hc404912;
      19477: inst = 32'h8220000;
      19478: inst = 32'h10408000;
      19479: inst = 32'hc404913;
      19480: inst = 32'h8220000;
      19481: inst = 32'h10408000;
      19482: inst = 32'hc404914;
      19483: inst = 32'h8220000;
      19484: inst = 32'h10408000;
      19485: inst = 32'hc404915;
      19486: inst = 32'h8220000;
      19487: inst = 32'h10408000;
      19488: inst = 32'hc404916;
      19489: inst = 32'h8220000;
      19490: inst = 32'h10408000;
      19491: inst = 32'hc404917;
      19492: inst = 32'h8220000;
      19493: inst = 32'h10408000;
      19494: inst = 32'hc404918;
      19495: inst = 32'h8220000;
      19496: inst = 32'h10408000;
      19497: inst = 32'hc404919;
      19498: inst = 32'h8220000;
      19499: inst = 32'h10408000;
      19500: inst = 32'hc40491a;
      19501: inst = 32'h8220000;
      19502: inst = 32'h10408000;
      19503: inst = 32'hc40491e;
      19504: inst = 32'h8220000;
      19505: inst = 32'h10408000;
      19506: inst = 32'hc40491f;
      19507: inst = 32'h8220000;
      19508: inst = 32'h10408000;
      19509: inst = 32'hc404920;
      19510: inst = 32'h8220000;
      19511: inst = 32'h10408000;
      19512: inst = 32'hc404921;
      19513: inst = 32'h8220000;
      19514: inst = 32'h10408000;
      19515: inst = 32'hc404922;
      19516: inst = 32'h8220000;
      19517: inst = 32'h10408000;
      19518: inst = 32'hc404923;
      19519: inst = 32'h8220000;
      19520: inst = 32'h10408000;
      19521: inst = 32'hc404924;
      19522: inst = 32'h8220000;
      19523: inst = 32'h10408000;
      19524: inst = 32'hc404925;
      19525: inst = 32'h8220000;
      19526: inst = 32'h10408000;
      19527: inst = 32'hc404926;
      19528: inst = 32'h8220000;
      19529: inst = 32'h10408000;
      19530: inst = 32'hc404927;
      19531: inst = 32'h8220000;
      19532: inst = 32'h10408000;
      19533: inst = 32'hc404929;
      19534: inst = 32'h8220000;
      19535: inst = 32'h10408000;
      19536: inst = 32'hc40492a;
      19537: inst = 32'h8220000;
      19538: inst = 32'h10408000;
      19539: inst = 32'hc40492b;
      19540: inst = 32'h8220000;
      19541: inst = 32'h10408000;
      19542: inst = 32'hc40492c;
      19543: inst = 32'h8220000;
      19544: inst = 32'h10408000;
      19545: inst = 32'hc40492d;
      19546: inst = 32'h8220000;
      19547: inst = 32'h10408000;
      19548: inst = 32'hc40492e;
      19549: inst = 32'h8220000;
      19550: inst = 32'h10408000;
      19551: inst = 32'hc40492f;
      19552: inst = 32'h8220000;
      19553: inst = 32'h10408000;
      19554: inst = 32'hc404930;
      19555: inst = 32'h8220000;
      19556: inst = 32'h10408000;
      19557: inst = 32'hc404931;
      19558: inst = 32'h8220000;
      19559: inst = 32'h10408000;
      19560: inst = 32'hc404932;
      19561: inst = 32'h8220000;
      19562: inst = 32'h10408000;
      19563: inst = 32'hc404933;
      19564: inst = 32'h8220000;
      19565: inst = 32'h10408000;
      19566: inst = 32'hc40494b;
      19567: inst = 32'h8220000;
      19568: inst = 32'h10408000;
      19569: inst = 32'hc40494c;
      19570: inst = 32'h8220000;
      19571: inst = 32'h10408000;
      19572: inst = 32'hc40494d;
      19573: inst = 32'h8220000;
      19574: inst = 32'h10408000;
      19575: inst = 32'hc40494e;
      19576: inst = 32'h8220000;
      19577: inst = 32'h10408000;
      19578: inst = 32'hc40494f;
      19579: inst = 32'h8220000;
      19580: inst = 32'h10408000;
      19581: inst = 32'hc404950;
      19582: inst = 32'h8220000;
      19583: inst = 32'h10408000;
      19584: inst = 32'hc404951;
      19585: inst = 32'h8220000;
      19586: inst = 32'h10408000;
      19587: inst = 32'hc404952;
      19588: inst = 32'h8220000;
      19589: inst = 32'h10408000;
      19590: inst = 32'hc404953;
      19591: inst = 32'h8220000;
      19592: inst = 32'h10408000;
      19593: inst = 32'hc404954;
      19594: inst = 32'h8220000;
      19595: inst = 32'h10408000;
      19596: inst = 32'hc404957;
      19597: inst = 32'h8220000;
      19598: inst = 32'h10408000;
      19599: inst = 32'hc404958;
      19600: inst = 32'h8220000;
      19601: inst = 32'h10408000;
      19602: inst = 32'hc404959;
      19603: inst = 32'h8220000;
      19604: inst = 32'h10408000;
      19605: inst = 32'hc40495a;
      19606: inst = 32'h8220000;
      19607: inst = 32'h10408000;
      19608: inst = 32'hc40495b;
      19609: inst = 32'h8220000;
      19610: inst = 32'h10408000;
      19611: inst = 32'hc40495c;
      19612: inst = 32'h8220000;
      19613: inst = 32'h10408000;
      19614: inst = 32'hc40495d;
      19615: inst = 32'h8220000;
      19616: inst = 32'h10408000;
      19617: inst = 32'hc40495e;
      19618: inst = 32'h8220000;
      19619: inst = 32'h10408000;
      19620: inst = 32'hc40495f;
      19621: inst = 32'h8220000;
      19622: inst = 32'h10408000;
      19623: inst = 32'hc404960;
      19624: inst = 32'h8220000;
      19625: inst = 32'h10408000;
      19626: inst = 32'hc404961;
      19627: inst = 32'h8220000;
      19628: inst = 32'h10408000;
      19629: inst = 32'hc404963;
      19630: inst = 32'h8220000;
      19631: inst = 32'h10408000;
      19632: inst = 32'hc404964;
      19633: inst = 32'h8220000;
      19634: inst = 32'h10408000;
      19635: inst = 32'hc404965;
      19636: inst = 32'h8220000;
      19637: inst = 32'h10408000;
      19638: inst = 32'hc404966;
      19639: inst = 32'h8220000;
      19640: inst = 32'h10408000;
      19641: inst = 32'hc404967;
      19642: inst = 32'h8220000;
      19643: inst = 32'h10408000;
      19644: inst = 32'hc404968;
      19645: inst = 32'h8220000;
      19646: inst = 32'h10408000;
      19647: inst = 32'hc404969;
      19648: inst = 32'h8220000;
      19649: inst = 32'h10408000;
      19650: inst = 32'hc40496a;
      19651: inst = 32'h8220000;
      19652: inst = 32'h10408000;
      19653: inst = 32'hc40496b;
      19654: inst = 32'h8220000;
      19655: inst = 32'h10408000;
      19656: inst = 32'hc40496c;
      19657: inst = 32'h8220000;
      19658: inst = 32'h10408000;
      19659: inst = 32'hc40496d;
      19660: inst = 32'h8220000;
      19661: inst = 32'h10408000;
      19662: inst = 32'hc404970;
      19663: inst = 32'h8220000;
      19664: inst = 32'h10408000;
      19665: inst = 32'hc404971;
      19666: inst = 32'h8220000;
      19667: inst = 32'h10408000;
      19668: inst = 32'hc404972;
      19669: inst = 32'h8220000;
      19670: inst = 32'h10408000;
      19671: inst = 32'hc404973;
      19672: inst = 32'h8220000;
      19673: inst = 32'h10408000;
      19674: inst = 32'hc404974;
      19675: inst = 32'h8220000;
      19676: inst = 32'h10408000;
      19677: inst = 32'hc404975;
      19678: inst = 32'h8220000;
      19679: inst = 32'h10408000;
      19680: inst = 32'hc404976;
      19681: inst = 32'h8220000;
      19682: inst = 32'h10408000;
      19683: inst = 32'hc404977;
      19684: inst = 32'h8220000;
      19685: inst = 32'h10408000;
      19686: inst = 32'hc404978;
      19687: inst = 32'h8220000;
      19688: inst = 32'h10408000;
      19689: inst = 32'hc404979;
      19690: inst = 32'h8220000;
      19691: inst = 32'h10408000;
      19692: inst = 32'hc40497d;
      19693: inst = 32'h8220000;
      19694: inst = 32'h10408000;
      19695: inst = 32'hc40497e;
      19696: inst = 32'h8220000;
      19697: inst = 32'h10408000;
      19698: inst = 32'hc40497f;
      19699: inst = 32'h8220000;
      19700: inst = 32'h10408000;
      19701: inst = 32'hc404980;
      19702: inst = 32'h8220000;
      19703: inst = 32'h10408000;
      19704: inst = 32'hc404981;
      19705: inst = 32'h8220000;
      19706: inst = 32'h10408000;
      19707: inst = 32'hc404982;
      19708: inst = 32'h8220000;
      19709: inst = 32'h10408000;
      19710: inst = 32'hc404983;
      19711: inst = 32'h8220000;
      19712: inst = 32'h10408000;
      19713: inst = 32'hc404984;
      19714: inst = 32'h8220000;
      19715: inst = 32'h10408000;
      19716: inst = 32'hc404985;
      19717: inst = 32'h8220000;
      19718: inst = 32'h10408000;
      19719: inst = 32'hc404986;
      19720: inst = 32'h8220000;
      19721: inst = 32'h10408000;
      19722: inst = 32'hc404987;
      19723: inst = 32'h8220000;
      19724: inst = 32'h10408000;
      19725: inst = 32'hc404989;
      19726: inst = 32'h8220000;
      19727: inst = 32'h10408000;
      19728: inst = 32'hc40498a;
      19729: inst = 32'h8220000;
      19730: inst = 32'h10408000;
      19731: inst = 32'hc40498b;
      19732: inst = 32'h8220000;
      19733: inst = 32'h10408000;
      19734: inst = 32'hc40498c;
      19735: inst = 32'h8220000;
      19736: inst = 32'h10408000;
      19737: inst = 32'hc40498d;
      19738: inst = 32'h8220000;
      19739: inst = 32'h10408000;
      19740: inst = 32'hc40498e;
      19741: inst = 32'h8220000;
      19742: inst = 32'h10408000;
      19743: inst = 32'hc40498f;
      19744: inst = 32'h8220000;
      19745: inst = 32'h10408000;
      19746: inst = 32'hc404990;
      19747: inst = 32'h8220000;
      19748: inst = 32'h10408000;
      19749: inst = 32'hc404991;
      19750: inst = 32'h8220000;
      19751: inst = 32'h10408000;
      19752: inst = 32'hc404992;
      19753: inst = 32'h8220000;
      19754: inst = 32'h10408000;
      19755: inst = 32'hc404993;
      19756: inst = 32'h8220000;
      19757: inst = 32'h10408000;
      19758: inst = 32'hc404dcd;
      19759: inst = 32'h8220000;
      19760: inst = 32'h10408000;
      19761: inst = 32'hc404dce;
      19762: inst = 32'h8220000;
      19763: inst = 32'h10408000;
      19764: inst = 32'hc404dcf;
      19765: inst = 32'h8220000;
      19766: inst = 32'h10408000;
      19767: inst = 32'hc404dd0;
      19768: inst = 32'h8220000;
      19769: inst = 32'h10408000;
      19770: inst = 32'hc404dd1;
      19771: inst = 32'h8220000;
      19772: inst = 32'h10408000;
      19773: inst = 32'hc404dd2;
      19774: inst = 32'h8220000;
      19775: inst = 32'h10408000;
      19776: inst = 32'hc404dd3;
      19777: inst = 32'h8220000;
      19778: inst = 32'h10408000;
      19779: inst = 32'hc404dd4;
      19780: inst = 32'h8220000;
      19781: inst = 32'h10408000;
      19782: inst = 32'hc404dd5;
      19783: inst = 32'h8220000;
      19784: inst = 32'h10408000;
      19785: inst = 32'hc404dd7;
      19786: inst = 32'h8220000;
      19787: inst = 32'h10408000;
      19788: inst = 32'hc404dd8;
      19789: inst = 32'h8220000;
      19790: inst = 32'h10408000;
      19791: inst = 32'hc404dd9;
      19792: inst = 32'h8220000;
      19793: inst = 32'h10408000;
      19794: inst = 32'hc404dda;
      19795: inst = 32'h8220000;
      19796: inst = 32'h10408000;
      19797: inst = 32'hc404ddb;
      19798: inst = 32'h8220000;
      19799: inst = 32'h10408000;
      19800: inst = 32'hc404ddc;
      19801: inst = 32'h8220000;
      19802: inst = 32'h10408000;
      19803: inst = 32'hc404ddd;
      19804: inst = 32'h8220000;
      19805: inst = 32'h10408000;
      19806: inst = 32'hc404dde;
      19807: inst = 32'h8220000;
      19808: inst = 32'h10408000;
      19809: inst = 32'hc404ddf;
      19810: inst = 32'h8220000;
      19811: inst = 32'h10408000;
      19812: inst = 32'hc404de0;
      19813: inst = 32'h8220000;
      19814: inst = 32'h10408000;
      19815: inst = 32'hc404de1;
      19816: inst = 32'h8220000;
      19817: inst = 32'h10408000;
      19818: inst = 32'hc404de2;
      19819: inst = 32'h8220000;
      19820: inst = 32'h10408000;
      19821: inst = 32'hc404de4;
      19822: inst = 32'h8220000;
      19823: inst = 32'h10408000;
      19824: inst = 32'hc404de5;
      19825: inst = 32'h8220000;
      19826: inst = 32'h10408000;
      19827: inst = 32'hc404de6;
      19828: inst = 32'h8220000;
      19829: inst = 32'h10408000;
      19830: inst = 32'hc404de7;
      19831: inst = 32'h8220000;
      19832: inst = 32'h10408000;
      19833: inst = 32'hc404de8;
      19834: inst = 32'h8220000;
      19835: inst = 32'h10408000;
      19836: inst = 32'hc404de9;
      19837: inst = 32'h8220000;
      19838: inst = 32'h10408000;
      19839: inst = 32'hc404dea;
      19840: inst = 32'h8220000;
      19841: inst = 32'h10408000;
      19842: inst = 32'hc404deb;
      19843: inst = 32'h8220000;
      19844: inst = 32'h10408000;
      19845: inst = 32'hc404dec;
      19846: inst = 32'h8220000;
      19847: inst = 32'h10408000;
      19848: inst = 32'hc404ded;
      19849: inst = 32'h8220000;
      19850: inst = 32'h10408000;
      19851: inst = 32'hc404df0;
      19852: inst = 32'h8220000;
      19853: inst = 32'h10408000;
      19854: inst = 32'hc404df1;
      19855: inst = 32'h8220000;
      19856: inst = 32'h10408000;
      19857: inst = 32'hc404df2;
      19858: inst = 32'h8220000;
      19859: inst = 32'h10408000;
      19860: inst = 32'hc404dfc;
      19861: inst = 32'h8220000;
      19862: inst = 32'h10408000;
      19863: inst = 32'hc404dfd;
      19864: inst = 32'h8220000;
      19865: inst = 32'h10408000;
      19866: inst = 32'hc404dfe;
      19867: inst = 32'h8220000;
      19868: inst = 32'h10408000;
      19869: inst = 32'hc404dff;
      19870: inst = 32'h8220000;
      19871: inst = 32'h10408000;
      19872: inst = 32'hc404e00;
      19873: inst = 32'h8220000;
      19874: inst = 32'h10408000;
      19875: inst = 32'hc404e01;
      19876: inst = 32'h8220000;
      19877: inst = 32'h10408000;
      19878: inst = 32'hc404e02;
      19879: inst = 32'h8220000;
      19880: inst = 32'h10408000;
      19881: inst = 32'hc404e03;
      19882: inst = 32'h8220000;
      19883: inst = 32'h10408000;
      19884: inst = 32'hc404e04;
      19885: inst = 32'h8220000;
      19886: inst = 32'h10408000;
      19887: inst = 32'hc404e05;
      19888: inst = 32'h8220000;
      19889: inst = 32'h10408000;
      19890: inst = 32'hc404e06;
      19891: inst = 32'h8220000;
      19892: inst = 32'h10408000;
      19893: inst = 32'hc404e07;
      19894: inst = 32'h8220000;
      19895: inst = 32'h10408000;
      19896: inst = 32'hc404e0b;
      19897: inst = 32'h8220000;
      19898: inst = 32'h10408000;
      19899: inst = 32'hc404e0c;
      19900: inst = 32'h8220000;
      19901: inst = 32'h10408000;
      19902: inst = 32'hc404e0d;
      19903: inst = 32'h8220000;
      19904: inst = 32'h10408000;
      19905: inst = 32'hc404e0e;
      19906: inst = 32'h8220000;
      19907: inst = 32'h10408000;
      19908: inst = 32'hc404e0f;
      19909: inst = 32'h8220000;
      19910: inst = 32'h10408000;
      19911: inst = 32'hc404e10;
      19912: inst = 32'h8220000;
      19913: inst = 32'h10408000;
      19914: inst = 32'hc404e11;
      19915: inst = 32'h8220000;
      19916: inst = 32'h10408000;
      19917: inst = 32'hc404e12;
      19918: inst = 32'h8220000;
      19919: inst = 32'h10408000;
      19920: inst = 32'hc404e13;
      19921: inst = 32'h8220000;
      19922: inst = 32'h10408000;
      19923: inst = 32'hc404e2c;
      19924: inst = 32'h8220000;
      19925: inst = 32'h10408000;
      19926: inst = 32'hc404e2d;
      19927: inst = 32'h8220000;
      19928: inst = 32'h10408000;
      19929: inst = 32'hc404e2e;
      19930: inst = 32'h8220000;
      19931: inst = 32'h10408000;
      19932: inst = 32'hc404e2f;
      19933: inst = 32'h8220000;
      19934: inst = 32'h10408000;
      19935: inst = 32'hc404e30;
      19936: inst = 32'h8220000;
      19937: inst = 32'h10408000;
      19938: inst = 32'hc404e31;
      19939: inst = 32'h8220000;
      19940: inst = 32'h10408000;
      19941: inst = 32'hc404e32;
      19942: inst = 32'h8220000;
      19943: inst = 32'h10408000;
      19944: inst = 32'hc404e33;
      19945: inst = 32'h8220000;
      19946: inst = 32'h10408000;
      19947: inst = 32'hc404e34;
      19948: inst = 32'h8220000;
      19949: inst = 32'h10408000;
      19950: inst = 32'hc404e35;
      19951: inst = 32'h8220000;
      19952: inst = 32'h10408000;
      19953: inst = 32'hc404e38;
      19954: inst = 32'h8220000;
      19955: inst = 32'h10408000;
      19956: inst = 32'hc404e39;
      19957: inst = 32'h8220000;
      19958: inst = 32'h10408000;
      19959: inst = 32'hc404e3a;
      19960: inst = 32'h8220000;
      19961: inst = 32'h10408000;
      19962: inst = 32'hc404e3b;
      19963: inst = 32'h8220000;
      19964: inst = 32'h10408000;
      19965: inst = 32'hc404e3c;
      19966: inst = 32'h8220000;
      19967: inst = 32'h10408000;
      19968: inst = 32'hc404e3d;
      19969: inst = 32'h8220000;
      19970: inst = 32'h10408000;
      19971: inst = 32'hc404e3e;
      19972: inst = 32'h8220000;
      19973: inst = 32'h10408000;
      19974: inst = 32'hc404e3f;
      19975: inst = 32'h8220000;
      19976: inst = 32'h10408000;
      19977: inst = 32'hc404e40;
      19978: inst = 32'h8220000;
      19979: inst = 32'h10408000;
      19980: inst = 32'hc404e41;
      19981: inst = 32'h8220000;
      19982: inst = 32'h10408000;
      19983: inst = 32'hc404e42;
      19984: inst = 32'h8220000;
      19985: inst = 32'h10408000;
      19986: inst = 32'hc404e44;
      19987: inst = 32'h8220000;
      19988: inst = 32'h10408000;
      19989: inst = 32'hc404e45;
      19990: inst = 32'h8220000;
      19991: inst = 32'h10408000;
      19992: inst = 32'hc404e46;
      19993: inst = 32'h8220000;
      19994: inst = 32'h10408000;
      19995: inst = 32'hc404e47;
      19996: inst = 32'h8220000;
      19997: inst = 32'h10408000;
      19998: inst = 32'hc404e48;
      19999: inst = 32'h8220000;
      20000: inst = 32'h10408000;
      20001: inst = 32'hc404e49;
      20002: inst = 32'h8220000;
      20003: inst = 32'h10408000;
      20004: inst = 32'hc404e4a;
      20005: inst = 32'h8220000;
      20006: inst = 32'h10408000;
      20007: inst = 32'hc404e4b;
      20008: inst = 32'h8220000;
      20009: inst = 32'h10408000;
      20010: inst = 32'hc404e4c;
      20011: inst = 32'h8220000;
      20012: inst = 32'h10408000;
      20013: inst = 32'hc404e4d;
      20014: inst = 32'h8220000;
      20015: inst = 32'h10408000;
      20016: inst = 32'hc404e50;
      20017: inst = 32'h8220000;
      20018: inst = 32'h10408000;
      20019: inst = 32'hc404e51;
      20020: inst = 32'h8220000;
      20021: inst = 32'h10408000;
      20022: inst = 32'hc404e52;
      20023: inst = 32'h8220000;
      20024: inst = 32'h10408000;
      20025: inst = 32'hc404e53;
      20026: inst = 32'h8220000;
      20027: inst = 32'h10408000;
      20028: inst = 32'hc404e5c;
      20029: inst = 32'h8220000;
      20030: inst = 32'h10408000;
      20031: inst = 32'hc404e5d;
      20032: inst = 32'h8220000;
      20033: inst = 32'h10408000;
      20034: inst = 32'hc404e5e;
      20035: inst = 32'h8220000;
      20036: inst = 32'h10408000;
      20037: inst = 32'hc404e5f;
      20038: inst = 32'h8220000;
      20039: inst = 32'h10408000;
      20040: inst = 32'hc404e60;
      20041: inst = 32'h8220000;
      20042: inst = 32'h10408000;
      20043: inst = 32'hc404e61;
      20044: inst = 32'h8220000;
      20045: inst = 32'h10408000;
      20046: inst = 32'hc404e62;
      20047: inst = 32'h8220000;
      20048: inst = 32'h10408000;
      20049: inst = 32'hc404e63;
      20050: inst = 32'h8220000;
      20051: inst = 32'h10408000;
      20052: inst = 32'hc404e64;
      20053: inst = 32'h8220000;
      20054: inst = 32'h10408000;
      20055: inst = 32'hc404e65;
      20056: inst = 32'h8220000;
      20057: inst = 32'h10408000;
      20058: inst = 32'hc404e66;
      20059: inst = 32'h8220000;
      20060: inst = 32'h10408000;
      20061: inst = 32'hc404e6a;
      20062: inst = 32'h8220000;
      20063: inst = 32'h10408000;
      20064: inst = 32'hc404e6b;
      20065: inst = 32'h8220000;
      20066: inst = 32'h10408000;
      20067: inst = 32'hc404e6c;
      20068: inst = 32'h8220000;
      20069: inst = 32'h10408000;
      20070: inst = 32'hc404e6d;
      20071: inst = 32'h8220000;
      20072: inst = 32'h10408000;
      20073: inst = 32'hc404e6e;
      20074: inst = 32'h8220000;
      20075: inst = 32'h10408000;
      20076: inst = 32'hc404e6f;
      20077: inst = 32'h8220000;
      20078: inst = 32'h10408000;
      20079: inst = 32'hc404e70;
      20080: inst = 32'h8220000;
      20081: inst = 32'h10408000;
      20082: inst = 32'hc404e71;
      20083: inst = 32'h8220000;
      20084: inst = 32'h10408000;
      20085: inst = 32'hc404e72;
      20086: inst = 32'h8220000;
      20087: inst = 32'h10408000;
      20088: inst = 32'hc404e73;
      20089: inst = 32'h8220000;
      20090: inst = 32'h10408000;
      20091: inst = 32'hc404e8b;
      20092: inst = 32'h8220000;
      20093: inst = 32'h10408000;
      20094: inst = 32'hc404e8c;
      20095: inst = 32'h8220000;
      20096: inst = 32'h10408000;
      20097: inst = 32'hc404e8d;
      20098: inst = 32'h8220000;
      20099: inst = 32'h10408000;
      20100: inst = 32'hc404e99;
      20101: inst = 32'h8220000;
      20102: inst = 32'h10408000;
      20103: inst = 32'hc404e9a;
      20104: inst = 32'h8220000;
      20105: inst = 32'h10408000;
      20106: inst = 32'hc404e9b;
      20107: inst = 32'h8220000;
      20108: inst = 32'h10408000;
      20109: inst = 32'hc404e9c;
      20110: inst = 32'h8220000;
      20111: inst = 32'h10408000;
      20112: inst = 32'hc404ea4;
      20113: inst = 32'h8220000;
      20114: inst = 32'h10408000;
      20115: inst = 32'hc404ea5;
      20116: inst = 32'h8220000;
      20117: inst = 32'h10408000;
      20118: inst = 32'hc404eac;
      20119: inst = 32'h8220000;
      20120: inst = 32'h10408000;
      20121: inst = 32'hc404ead;
      20122: inst = 32'h8220000;
      20123: inst = 32'h10408000;
      20124: inst = 32'hc404eb0;
      20125: inst = 32'h8220000;
      20126: inst = 32'h10408000;
      20127: inst = 32'hc404eb1;
      20128: inst = 32'h8220000;
      20129: inst = 32'h10408000;
      20130: inst = 32'hc404eb2;
      20131: inst = 32'h8220000;
      20132: inst = 32'h10408000;
      20133: inst = 32'hc404eb3;
      20134: inst = 32'h8220000;
      20135: inst = 32'h10408000;
      20136: inst = 32'hc404eb4;
      20137: inst = 32'h8220000;
      20138: inst = 32'h10408000;
      20139: inst = 32'hc404ebc;
      20140: inst = 32'h8220000;
      20141: inst = 32'h10408000;
      20142: inst = 32'hc404ebd;
      20143: inst = 32'h8220000;
      20144: inst = 32'h10408000;
      20145: inst = 32'hc404ec2;
      20146: inst = 32'h8220000;
      20147: inst = 32'h10408000;
      20148: inst = 32'hc404ec3;
      20149: inst = 32'h8220000;
      20150: inst = 32'h10408000;
      20151: inst = 32'hc404ec4;
      20152: inst = 32'h8220000;
      20153: inst = 32'h10408000;
      20154: inst = 32'hc404ec5;
      20155: inst = 32'h8220000;
      20156: inst = 32'h10408000;
      20157: inst = 32'hc404ec9;
      20158: inst = 32'h8220000;
      20159: inst = 32'h10408000;
      20160: inst = 32'hc404eca;
      20161: inst = 32'h8220000;
      20162: inst = 32'h10408000;
      20163: inst = 32'hc404eeb;
      20164: inst = 32'h8220000;
      20165: inst = 32'h10408000;
      20166: inst = 32'hc404eec;
      20167: inst = 32'h8220000;
      20168: inst = 32'h10408000;
      20169: inst = 32'hc404efa;
      20170: inst = 32'h8220000;
      20171: inst = 32'h10408000;
      20172: inst = 32'hc404efb;
      20173: inst = 32'h8220000;
      20174: inst = 32'h10408000;
      20175: inst = 32'hc404efc;
      20176: inst = 32'h8220000;
      20177: inst = 32'h10408000;
      20178: inst = 32'hc404f04;
      20179: inst = 32'h8220000;
      20180: inst = 32'h10408000;
      20181: inst = 32'hc404f05;
      20182: inst = 32'h8220000;
      20183: inst = 32'h10408000;
      20184: inst = 32'hc404f0c;
      20185: inst = 32'h8220000;
      20186: inst = 32'h10408000;
      20187: inst = 32'hc404f0d;
      20188: inst = 32'h8220000;
      20189: inst = 32'h10408000;
      20190: inst = 32'hc404f10;
      20191: inst = 32'h8220000;
      20192: inst = 32'h10408000;
      20193: inst = 32'hc404f12;
      20194: inst = 32'h8220000;
      20195: inst = 32'h10408000;
      20196: inst = 32'hc404f13;
      20197: inst = 32'h8220000;
      20198: inst = 32'h10408000;
      20199: inst = 32'hc404f14;
      20200: inst = 32'h8220000;
      20201: inst = 32'h10408000;
      20202: inst = 32'hc404f15;
      20203: inst = 32'h8220000;
      20204: inst = 32'h10408000;
      20205: inst = 32'hc404f1c;
      20206: inst = 32'h8220000;
      20207: inst = 32'h10408000;
      20208: inst = 32'hc404f1d;
      20209: inst = 32'h8220000;
      20210: inst = 32'h10408000;
      20211: inst = 32'hc404f22;
      20212: inst = 32'h8220000;
      20213: inst = 32'h10408000;
      20214: inst = 32'hc404f23;
      20215: inst = 32'h8220000;
      20216: inst = 32'h10408000;
      20217: inst = 32'hc404f24;
      20218: inst = 32'h8220000;
      20219: inst = 32'h10408000;
      20220: inst = 32'hc404f29;
      20221: inst = 32'h8220000;
      20222: inst = 32'h10408000;
      20223: inst = 32'hc404f2a;
      20224: inst = 32'h8220000;
      20225: inst = 32'h10408000;
      20226: inst = 32'hc404f4b;
      20227: inst = 32'h8220000;
      20228: inst = 32'h10408000;
      20229: inst = 32'hc404f4c;
      20230: inst = 32'h8220000;
      20231: inst = 32'h10408000;
      20232: inst = 32'hc404f4e;
      20233: inst = 32'h8220000;
      20234: inst = 32'h10408000;
      20235: inst = 32'hc404f4f;
      20236: inst = 32'h8220000;
      20237: inst = 32'h10408000;
      20238: inst = 32'hc404f50;
      20239: inst = 32'h8220000;
      20240: inst = 32'h10408000;
      20241: inst = 32'hc404f51;
      20242: inst = 32'h8220000;
      20243: inst = 32'h10408000;
      20244: inst = 32'hc404f52;
      20245: inst = 32'h8220000;
      20246: inst = 32'h10408000;
      20247: inst = 32'hc404f5b;
      20248: inst = 32'h8220000;
      20249: inst = 32'h10408000;
      20250: inst = 32'hc404f5c;
      20251: inst = 32'h8220000;
      20252: inst = 32'h10408000;
      20253: inst = 32'hc404f5d;
      20254: inst = 32'h8220000;
      20255: inst = 32'h10408000;
      20256: inst = 32'hc404f64;
      20257: inst = 32'h8220000;
      20258: inst = 32'h10408000;
      20259: inst = 32'hc404f65;
      20260: inst = 32'h8220000;
      20261: inst = 32'h10408000;
      20262: inst = 32'hc404f6c;
      20263: inst = 32'h8220000;
      20264: inst = 32'h10408000;
      20265: inst = 32'hc404f70;
      20266: inst = 32'h8220000;
      20267: inst = 32'h10408000;
      20268: inst = 32'hc404f71;
      20269: inst = 32'h8220000;
      20270: inst = 32'h10408000;
      20271: inst = 32'hc404f72;
      20272: inst = 32'h8220000;
      20273: inst = 32'h10408000;
      20274: inst = 32'hc404f73;
      20275: inst = 32'h8220000;
      20276: inst = 32'h10408000;
      20277: inst = 32'hc404f74;
      20278: inst = 32'h8220000;
      20279: inst = 32'h10408000;
      20280: inst = 32'hc404f75;
      20281: inst = 32'h8220000;
      20282: inst = 32'h10408000;
      20283: inst = 32'hc404f76;
      20284: inst = 32'h8220000;
      20285: inst = 32'h10408000;
      20286: inst = 32'hc404f7c;
      20287: inst = 32'h8220000;
      20288: inst = 32'h10408000;
      20289: inst = 32'hc404f7d;
      20290: inst = 32'h8220000;
      20291: inst = 32'h10408000;
      20292: inst = 32'hc404f7f;
      20293: inst = 32'h8220000;
      20294: inst = 32'h10408000;
      20295: inst = 32'hc404f80;
      20296: inst = 32'h8220000;
      20297: inst = 32'h10408000;
      20298: inst = 32'hc404f81;
      20299: inst = 32'h8220000;
      20300: inst = 32'h10408000;
      20301: inst = 32'hc404f82;
      20302: inst = 32'h8220000;
      20303: inst = 32'h10408000;
      20304: inst = 32'hc404f83;
      20305: inst = 32'h8220000;
      20306: inst = 32'h10408000;
      20307: inst = 32'hc404f89;
      20308: inst = 32'h8220000;
      20309: inst = 32'h10408000;
      20310: inst = 32'hc404f8a;
      20311: inst = 32'h8220000;
      20312: inst = 32'h10408000;
      20313: inst = 32'hc404f8c;
      20314: inst = 32'h8220000;
      20315: inst = 32'h10408000;
      20316: inst = 32'hc404f8d;
      20317: inst = 32'h8220000;
      20318: inst = 32'h10408000;
      20319: inst = 32'hc404f8e;
      20320: inst = 32'h8220000;
      20321: inst = 32'h10408000;
      20322: inst = 32'hc404f8f;
      20323: inst = 32'h8220000;
      20324: inst = 32'h10408000;
      20325: inst = 32'hc404f90;
      20326: inst = 32'h8220000;
      20327: inst = 32'h10408000;
      20328: inst = 32'hc404fab;
      20329: inst = 32'h8220000;
      20330: inst = 32'h10408000;
      20331: inst = 32'hc404fac;
      20332: inst = 32'h8220000;
      20333: inst = 32'h10408000;
      20334: inst = 32'hc404fae;
      20335: inst = 32'h8220000;
      20336: inst = 32'h10408000;
      20337: inst = 32'hc404faf;
      20338: inst = 32'h8220000;
      20339: inst = 32'h10408000;
      20340: inst = 32'hc404fb0;
      20341: inst = 32'h8220000;
      20342: inst = 32'h10408000;
      20343: inst = 32'hc404fb1;
      20344: inst = 32'h8220000;
      20345: inst = 32'h10408000;
      20346: inst = 32'hc404fb2;
      20347: inst = 32'h8220000;
      20348: inst = 32'h10408000;
      20349: inst = 32'hc404fbc;
      20350: inst = 32'h8220000;
      20351: inst = 32'h10408000;
      20352: inst = 32'hc404fbd;
      20353: inst = 32'h8220000;
      20354: inst = 32'h10408000;
      20355: inst = 32'hc404fbe;
      20356: inst = 32'h8220000;
      20357: inst = 32'h10408000;
      20358: inst = 32'hc404fc4;
      20359: inst = 32'h8220000;
      20360: inst = 32'h10408000;
      20361: inst = 32'hc404fc5;
      20362: inst = 32'h8220000;
      20363: inst = 32'h10408000;
      20364: inst = 32'hc404fd0;
      20365: inst = 32'h8220000;
      20366: inst = 32'h10408000;
      20367: inst = 32'hc404fd1;
      20368: inst = 32'h8220000;
      20369: inst = 32'h10408000;
      20370: inst = 32'hc404fd2;
      20371: inst = 32'h8220000;
      20372: inst = 32'h10408000;
      20373: inst = 32'hc404fd4;
      20374: inst = 32'h8220000;
      20375: inst = 32'h10408000;
      20376: inst = 32'hc404fd5;
      20377: inst = 32'h8220000;
      20378: inst = 32'h10408000;
      20379: inst = 32'hc404fd6;
      20380: inst = 32'h8220000;
      20381: inst = 32'h10408000;
      20382: inst = 32'hc404fd7;
      20383: inst = 32'h8220000;
      20384: inst = 32'h10408000;
      20385: inst = 32'hc404fdc;
      20386: inst = 32'h8220000;
      20387: inst = 32'h10408000;
      20388: inst = 32'hc404fdd;
      20389: inst = 32'h8220000;
      20390: inst = 32'h10408000;
      20391: inst = 32'hc404fdf;
      20392: inst = 32'h8220000;
      20393: inst = 32'h10408000;
      20394: inst = 32'hc404fe0;
      20395: inst = 32'h8220000;
      20396: inst = 32'h10408000;
      20397: inst = 32'hc404fe1;
      20398: inst = 32'h8220000;
      20399: inst = 32'h10408000;
      20400: inst = 32'hc404fe2;
      20401: inst = 32'h8220000;
      20402: inst = 32'h10408000;
      20403: inst = 32'hc404fe9;
      20404: inst = 32'h8220000;
      20405: inst = 32'h10408000;
      20406: inst = 32'hc404fea;
      20407: inst = 32'h8220000;
      20408: inst = 32'h10408000;
      20409: inst = 32'hc404fec;
      20410: inst = 32'h8220000;
      20411: inst = 32'h10408000;
      20412: inst = 32'hc404fed;
      20413: inst = 32'h8220000;
      20414: inst = 32'h10408000;
      20415: inst = 32'hc404fee;
      20416: inst = 32'h8220000;
      20417: inst = 32'h10408000;
      20418: inst = 32'hc404fef;
      20419: inst = 32'h8220000;
      20420: inst = 32'h10408000;
      20421: inst = 32'hc404ff0;
      20422: inst = 32'h8220000;
      20423: inst = 32'h10408000;
      20424: inst = 32'hc40500b;
      20425: inst = 32'h8220000;
      20426: inst = 32'h10408000;
      20427: inst = 32'hc40500c;
      20428: inst = 32'h8220000;
      20429: inst = 32'h10408000;
      20430: inst = 32'hc40501d;
      20431: inst = 32'h8220000;
      20432: inst = 32'h10408000;
      20433: inst = 32'hc40501e;
      20434: inst = 32'h8220000;
      20435: inst = 32'h10408000;
      20436: inst = 32'hc40501f;
      20437: inst = 32'h8220000;
      20438: inst = 32'h10408000;
      20439: inst = 32'hc405024;
      20440: inst = 32'h8220000;
      20441: inst = 32'h10408000;
      20442: inst = 32'hc405025;
      20443: inst = 32'h8220000;
      20444: inst = 32'h10408000;
      20445: inst = 32'hc405030;
      20446: inst = 32'h8220000;
      20447: inst = 32'h10408000;
      20448: inst = 32'hc405031;
      20449: inst = 32'h8220000;
      20450: inst = 32'h10408000;
      20451: inst = 32'hc405032;
      20452: inst = 32'h8220000;
      20453: inst = 32'h10408000;
      20454: inst = 32'hc405033;
      20455: inst = 32'h8220000;
      20456: inst = 32'h10408000;
      20457: inst = 32'hc405034;
      20458: inst = 32'h8220000;
      20459: inst = 32'h10408000;
      20460: inst = 32'hc405035;
      20461: inst = 32'h8220000;
      20462: inst = 32'h10408000;
      20463: inst = 32'hc405036;
      20464: inst = 32'h8220000;
      20465: inst = 32'h10408000;
      20466: inst = 32'hc405037;
      20467: inst = 32'h8220000;
      20468: inst = 32'h10408000;
      20469: inst = 32'hc405038;
      20470: inst = 32'h8220000;
      20471: inst = 32'h10408000;
      20472: inst = 32'hc40503c;
      20473: inst = 32'h8220000;
      20474: inst = 32'h10408000;
      20475: inst = 32'hc40503d;
      20476: inst = 32'h8220000;
      20477: inst = 32'h10408000;
      20478: inst = 32'hc405049;
      20479: inst = 32'h8220000;
      20480: inst = 32'h10408000;
      20481: inst = 32'hc40504a;
      20482: inst = 32'h8220000;
      20483: inst = 32'h10408000;
      20484: inst = 32'hc40506b;
      20485: inst = 32'h8220000;
      20486: inst = 32'h10408000;
      20487: inst = 32'hc40506c;
      20488: inst = 32'h8220000;
      20489: inst = 32'h10408000;
      20490: inst = 32'hc40506d;
      20491: inst = 32'h8220000;
      20492: inst = 32'h10408000;
      20493: inst = 32'hc40506e;
      20494: inst = 32'h8220000;
      20495: inst = 32'h10408000;
      20496: inst = 32'hc40506f;
      20497: inst = 32'h8220000;
      20498: inst = 32'h10408000;
      20499: inst = 32'hc405070;
      20500: inst = 32'h8220000;
      20501: inst = 32'h10408000;
      20502: inst = 32'hc405071;
      20503: inst = 32'h8220000;
      20504: inst = 32'h10408000;
      20505: inst = 32'hc405072;
      20506: inst = 32'h8220000;
      20507: inst = 32'h10408000;
      20508: inst = 32'hc405073;
      20509: inst = 32'h8220000;
      20510: inst = 32'h10408000;
      20511: inst = 32'hc405074;
      20512: inst = 32'h8220000;
      20513: inst = 32'h10408000;
      20514: inst = 32'hc405075;
      20515: inst = 32'h8220000;
      20516: inst = 32'h10408000;
      20517: inst = 32'hc405077;
      20518: inst = 32'h8220000;
      20519: inst = 32'h10408000;
      20520: inst = 32'hc405078;
      20521: inst = 32'h8220000;
      20522: inst = 32'h10408000;
      20523: inst = 32'hc405079;
      20524: inst = 32'h8220000;
      20525: inst = 32'h10408000;
      20526: inst = 32'hc40507a;
      20527: inst = 32'h8220000;
      20528: inst = 32'h10408000;
      20529: inst = 32'hc40507b;
      20530: inst = 32'h8220000;
      20531: inst = 32'h10408000;
      20532: inst = 32'hc40507c;
      20533: inst = 32'h8220000;
      20534: inst = 32'h10408000;
      20535: inst = 32'hc40507d;
      20536: inst = 32'h8220000;
      20537: inst = 32'h10408000;
      20538: inst = 32'hc40507e;
      20539: inst = 32'h8220000;
      20540: inst = 32'h10408000;
      20541: inst = 32'hc40507f;
      20542: inst = 32'h8220000;
      20543: inst = 32'h10408000;
      20544: inst = 32'hc405080;
      20545: inst = 32'h8220000;
      20546: inst = 32'h10408000;
      20547: inst = 32'hc405084;
      20548: inst = 32'h8220000;
      20549: inst = 32'h10408000;
      20550: inst = 32'hc405085;
      20551: inst = 32'h8220000;
      20552: inst = 32'h10408000;
      20553: inst = 32'hc405086;
      20554: inst = 32'h8220000;
      20555: inst = 32'h10408000;
      20556: inst = 32'hc405087;
      20557: inst = 32'h8220000;
      20558: inst = 32'h10408000;
      20559: inst = 32'hc405088;
      20560: inst = 32'h8220000;
      20561: inst = 32'h10408000;
      20562: inst = 32'hc405089;
      20563: inst = 32'h8220000;
      20564: inst = 32'h10408000;
      20565: inst = 32'hc40508a;
      20566: inst = 32'h8220000;
      20567: inst = 32'h10408000;
      20568: inst = 32'hc40508b;
      20569: inst = 32'h8220000;
      20570: inst = 32'h10408000;
      20571: inst = 32'hc40508c;
      20572: inst = 32'h8220000;
      20573: inst = 32'h10408000;
      20574: inst = 32'hc40508d;
      20575: inst = 32'h8220000;
      20576: inst = 32'h10408000;
      20577: inst = 32'hc405090;
      20578: inst = 32'h8220000;
      20579: inst = 32'h10408000;
      20580: inst = 32'hc405091;
      20581: inst = 32'h8220000;
      20582: inst = 32'h10408000;
      20583: inst = 32'hc405096;
      20584: inst = 32'h8220000;
      20585: inst = 32'h10408000;
      20586: inst = 32'hc405097;
      20587: inst = 32'h8220000;
      20588: inst = 32'h10408000;
      20589: inst = 32'hc405098;
      20590: inst = 32'h8220000;
      20591: inst = 32'h10408000;
      20592: inst = 32'hc405099;
      20593: inst = 32'h8220000;
      20594: inst = 32'h10408000;
      20595: inst = 32'hc40509c;
      20596: inst = 32'h8220000;
      20597: inst = 32'h10408000;
      20598: inst = 32'hc40509d;
      20599: inst = 32'h8220000;
      20600: inst = 32'h10408000;
      20601: inst = 32'hc4050a9;
      20602: inst = 32'h8220000;
      20603: inst = 32'h10408000;
      20604: inst = 32'hc4050aa;
      20605: inst = 32'h8220000;
      20606: inst = 32'h10408000;
      20607: inst = 32'hc4050ab;
      20608: inst = 32'h8220000;
      20609: inst = 32'h10408000;
      20610: inst = 32'hc4050ac;
      20611: inst = 32'h8220000;
      20612: inst = 32'h10408000;
      20613: inst = 32'hc4050ad;
      20614: inst = 32'h8220000;
      20615: inst = 32'h10408000;
      20616: inst = 32'hc4050ae;
      20617: inst = 32'h8220000;
      20618: inst = 32'h10408000;
      20619: inst = 32'hc4050af;
      20620: inst = 32'h8220000;
      20621: inst = 32'h10408000;
      20622: inst = 32'hc4050b0;
      20623: inst = 32'h8220000;
      20624: inst = 32'h10408000;
      20625: inst = 32'hc4050b1;
      20626: inst = 32'h8220000;
      20627: inst = 32'h10408000;
      20628: inst = 32'hc4050b2;
      20629: inst = 32'h8220000;
      20630: inst = 32'h10408000;
      20631: inst = 32'hc4050b3;
      20632: inst = 32'h8220000;
      20633: inst = 32'h10408000;
      20634: inst = 32'hc4050cb;
      20635: inst = 32'h8220000;
      20636: inst = 32'h10408000;
      20637: inst = 32'hc4050cc;
      20638: inst = 32'h8220000;
      20639: inst = 32'h10408000;
      20640: inst = 32'hc4050cd;
      20641: inst = 32'h8220000;
      20642: inst = 32'h10408000;
      20643: inst = 32'hc4050ce;
      20644: inst = 32'h8220000;
      20645: inst = 32'h10408000;
      20646: inst = 32'hc4050cf;
      20647: inst = 32'h8220000;
      20648: inst = 32'h10408000;
      20649: inst = 32'hc4050d0;
      20650: inst = 32'h8220000;
      20651: inst = 32'h10408000;
      20652: inst = 32'hc4050d1;
      20653: inst = 32'h8220000;
      20654: inst = 32'h10408000;
      20655: inst = 32'hc4050d2;
      20656: inst = 32'h8220000;
      20657: inst = 32'h10408000;
      20658: inst = 32'hc4050d3;
      20659: inst = 32'h8220000;
      20660: inst = 32'h10408000;
      20661: inst = 32'hc4050d4;
      20662: inst = 32'h8220000;
      20663: inst = 32'h10408000;
      20664: inst = 32'hc4050d7;
      20665: inst = 32'h8220000;
      20666: inst = 32'h10408000;
      20667: inst = 32'hc4050d8;
      20668: inst = 32'h8220000;
      20669: inst = 32'h10408000;
      20670: inst = 32'hc4050d9;
      20671: inst = 32'h8220000;
      20672: inst = 32'h10408000;
      20673: inst = 32'hc4050da;
      20674: inst = 32'h8220000;
      20675: inst = 32'h10408000;
      20676: inst = 32'hc4050db;
      20677: inst = 32'h8220000;
      20678: inst = 32'h10408000;
      20679: inst = 32'hc4050dc;
      20680: inst = 32'h8220000;
      20681: inst = 32'h10408000;
      20682: inst = 32'hc4050dd;
      20683: inst = 32'h8220000;
      20684: inst = 32'h10408000;
      20685: inst = 32'hc4050de;
      20686: inst = 32'h8220000;
      20687: inst = 32'h10408000;
      20688: inst = 32'hc4050df;
      20689: inst = 32'h8220000;
      20690: inst = 32'h10408000;
      20691: inst = 32'hc4050e0;
      20692: inst = 32'h8220000;
      20693: inst = 32'h10408000;
      20694: inst = 32'hc4050e1;
      20695: inst = 32'h8220000;
      20696: inst = 32'h10408000;
      20697: inst = 32'hc4050e5;
      20698: inst = 32'h8220000;
      20699: inst = 32'h10408000;
      20700: inst = 32'hc4050e6;
      20701: inst = 32'h8220000;
      20702: inst = 32'h10408000;
      20703: inst = 32'hc4050e7;
      20704: inst = 32'h8220000;
      20705: inst = 32'h10408000;
      20706: inst = 32'hc4050e8;
      20707: inst = 32'h8220000;
      20708: inst = 32'h10408000;
      20709: inst = 32'hc4050e9;
      20710: inst = 32'h8220000;
      20711: inst = 32'h10408000;
      20712: inst = 32'hc4050ea;
      20713: inst = 32'h8220000;
      20714: inst = 32'h10408000;
      20715: inst = 32'hc4050eb;
      20716: inst = 32'h8220000;
      20717: inst = 32'h10408000;
      20718: inst = 32'hc4050ec;
      20719: inst = 32'h8220000;
      20720: inst = 32'h10408000;
      20721: inst = 32'hc4050ed;
      20722: inst = 32'h8220000;
      20723: inst = 32'h10408000;
      20724: inst = 32'hc4050f0;
      20725: inst = 32'h8220000;
      20726: inst = 32'h10408000;
      20727: inst = 32'hc4050f1;
      20728: inst = 32'h8220000;
      20729: inst = 32'h10408000;
      20730: inst = 32'hc4050f6;
      20731: inst = 32'h8220000;
      20732: inst = 32'h10408000;
      20733: inst = 32'hc4050f7;
      20734: inst = 32'h8220000;
      20735: inst = 32'h10408000;
      20736: inst = 32'hc4050f8;
      20737: inst = 32'h8220000;
      20738: inst = 32'h10408000;
      20739: inst = 32'hc4050f9;
      20740: inst = 32'h8220000;
      20741: inst = 32'h10408000;
      20742: inst = 32'hc4050fa;
      20743: inst = 32'h8220000;
      20744: inst = 32'h10408000;
      20745: inst = 32'hc4050fc;
      20746: inst = 32'h8220000;
      20747: inst = 32'h10408000;
      20748: inst = 32'hc4050fd;
      20749: inst = 32'h8220000;
      20750: inst = 32'h10408000;
      20751: inst = 32'hc405109;
      20752: inst = 32'h8220000;
      20753: inst = 32'h10408000;
      20754: inst = 32'hc40510a;
      20755: inst = 32'h8220000;
      20756: inst = 32'h10408000;
      20757: inst = 32'hc40510b;
      20758: inst = 32'h8220000;
      20759: inst = 32'h10408000;
      20760: inst = 32'hc40510c;
      20761: inst = 32'h8220000;
      20762: inst = 32'h10408000;
      20763: inst = 32'hc40510d;
      20764: inst = 32'h8220000;
      20765: inst = 32'h10408000;
      20766: inst = 32'hc40510e;
      20767: inst = 32'h8220000;
      20768: inst = 32'h10408000;
      20769: inst = 32'hc40510f;
      20770: inst = 32'h8220000;
      20771: inst = 32'h10408000;
      20772: inst = 32'hc405110;
      20773: inst = 32'h8220000;
      20774: inst = 32'h10408000;
      20775: inst = 32'hc405111;
      20776: inst = 32'h8220000;
      20777: inst = 32'h10408000;
      20778: inst = 32'hc405112;
      20779: inst = 32'h8220000;
      20780: inst = 32'h10408000;
      20781: inst = 32'hc405113;
      20782: inst = 32'h8220000;
      20783: inst = 32'h58000000;
      20784: inst = 32'h29c20000;
      20785: inst = 32'h29e30000;
      20786: inst = 32'h11600000;
      20787: inst = 32'hd600060;
      20788: inst = 32'h12208000;
      20789: inst = 32'he203fe0;
      20790: inst = 32'h13e00000;
      20791: inst = 32'hfe0514e;
      20792: inst = 32'h20200000;
      20793: inst = 32'h5be00000;
      20794: inst = 32'h13e00000;
      20795: inst = 32'hfe05d1d;
      20796: inst = 32'h20200001;
      20797: inst = 32'h5be00000;
      20798: inst = 32'h13e00000;
      20799: inst = 32'hfe05d1d;
      20800: inst = 32'h20200002;
      20801: inst = 32'h5be00000;
      20802: inst = 32'h13e00000;
      20803: inst = 32'hfe05943;
      20804: inst = 32'h20200003;
      20805: inst = 32'h5be00000;
      20806: inst = 32'h13e00000;
      20807: inst = 32'hfe05943;
      20808: inst = 32'h20200004;
      20809: inst = 32'h5be00000;
      20810: inst = 32'h13e00000;
      20811: inst = 32'hfe05553;
      20812: inst = 32'h20200005;
      20813: inst = 32'h5be00000;
      20814: inst = 32'hc6018c3;
      20815: inst = 32'h2a0e0000;
      20816: inst = 32'h294f0000;
      20817: inst = 32'h11200000;
      20818: inst = 32'hd205156;
      20819: inst = 32'h13e00000;
      20820: inst = 32'hfe0a9ea;
      20821: inst = 32'h5be00000;
      20822: inst = 32'h244c8000;
      20823: inst = 32'h24428800;
      20824: inst = 32'h8620000;
      20825: inst = 32'h2a0e0001;
      20826: inst = 32'h294f0000;
      20827: inst = 32'h11200000;
      20828: inst = 32'hd205160;
      20829: inst = 32'h13e00000;
      20830: inst = 32'hfe0a9ea;
      20831: inst = 32'h5be00000;
      20832: inst = 32'h244c8000;
      20833: inst = 32'h24428800;
      20834: inst = 32'h8620000;
      20835: inst = 32'h2a0e0002;
      20836: inst = 32'h294f0000;
      20837: inst = 32'h11200000;
      20838: inst = 32'hd20516a;
      20839: inst = 32'h13e00000;
      20840: inst = 32'hfe0a9ea;
      20841: inst = 32'h5be00000;
      20842: inst = 32'h244c8000;
      20843: inst = 32'h24428800;
      20844: inst = 32'h8620000;
      20845: inst = 32'h2a0e0003;
      20846: inst = 32'h294f0000;
      20847: inst = 32'h11200000;
      20848: inst = 32'hd205174;
      20849: inst = 32'h13e00000;
      20850: inst = 32'hfe0a9ea;
      20851: inst = 32'h5be00000;
      20852: inst = 32'h244c8000;
      20853: inst = 32'h24428800;
      20854: inst = 32'h8620000;
      20855: inst = 32'h2a0e0004;
      20856: inst = 32'h294f0000;
      20857: inst = 32'h11200000;
      20858: inst = 32'hd20517e;
      20859: inst = 32'h13e00000;
      20860: inst = 32'hfe0a9ea;
      20861: inst = 32'h5be00000;
      20862: inst = 32'h244c8000;
      20863: inst = 32'h24428800;
      20864: inst = 32'h8620000;
      20865: inst = 32'h2a0e0005;
      20866: inst = 32'h294f0000;
      20867: inst = 32'h11200000;
      20868: inst = 32'hd205188;
      20869: inst = 32'h13e00000;
      20870: inst = 32'hfe0a9ea;
      20871: inst = 32'h5be00000;
      20872: inst = 32'h244c8000;
      20873: inst = 32'h24428800;
      20874: inst = 32'h8620000;
      20875: inst = 32'h2a0e0006;
      20876: inst = 32'h294f0000;
      20877: inst = 32'h11200000;
      20878: inst = 32'hd205192;
      20879: inst = 32'h13e00000;
      20880: inst = 32'hfe0a9ea;
      20881: inst = 32'h5be00000;
      20882: inst = 32'h244c8000;
      20883: inst = 32'h24428800;
      20884: inst = 32'h8620000;
      20885: inst = 32'h2a0e0007;
      20886: inst = 32'h294f0000;
      20887: inst = 32'h11200000;
      20888: inst = 32'hd20519c;
      20889: inst = 32'h13e00000;
      20890: inst = 32'hfe0a9ea;
      20891: inst = 32'h5be00000;
      20892: inst = 32'h244c8000;
      20893: inst = 32'h24428800;
      20894: inst = 32'h8620000;
      20895: inst = 32'h2a0e0008;
      20896: inst = 32'h294f0000;
      20897: inst = 32'h11200000;
      20898: inst = 32'hd2051a6;
      20899: inst = 32'h13e00000;
      20900: inst = 32'hfe0a9ea;
      20901: inst = 32'h5be00000;
      20902: inst = 32'h244c8000;
      20903: inst = 32'h24428800;
      20904: inst = 32'h8620000;
      20905: inst = 32'h2a0e0009;
      20906: inst = 32'h294f0000;
      20907: inst = 32'h11200000;
      20908: inst = 32'hd2051b0;
      20909: inst = 32'h13e00000;
      20910: inst = 32'hfe0a9ea;
      20911: inst = 32'h5be00000;
      20912: inst = 32'h244c8000;
      20913: inst = 32'h24428800;
      20914: inst = 32'h8620000;
      20915: inst = 32'h2a0e0000;
      20916: inst = 32'h294f0001;
      20917: inst = 32'h11200000;
      20918: inst = 32'hd2051ba;
      20919: inst = 32'h13e00000;
      20920: inst = 32'hfe0a9ea;
      20921: inst = 32'h5be00000;
      20922: inst = 32'h244c8000;
      20923: inst = 32'h24428800;
      20924: inst = 32'h8620000;
      20925: inst = 32'h2a0e0001;
      20926: inst = 32'h294f0001;
      20927: inst = 32'h11200000;
      20928: inst = 32'hd2051c4;
      20929: inst = 32'h13e00000;
      20930: inst = 32'hfe0a9ea;
      20931: inst = 32'h5be00000;
      20932: inst = 32'h244c8000;
      20933: inst = 32'h24428800;
      20934: inst = 32'h8620000;
      20935: inst = 32'h2a0e0002;
      20936: inst = 32'h294f0001;
      20937: inst = 32'h11200000;
      20938: inst = 32'hd2051ce;
      20939: inst = 32'h13e00000;
      20940: inst = 32'hfe0a9ea;
      20941: inst = 32'h5be00000;
      20942: inst = 32'h244c8000;
      20943: inst = 32'h24428800;
      20944: inst = 32'h8620000;
      20945: inst = 32'h2a0e0003;
      20946: inst = 32'h294f0001;
      20947: inst = 32'h11200000;
      20948: inst = 32'hd2051d8;
      20949: inst = 32'h13e00000;
      20950: inst = 32'hfe0a9ea;
      20951: inst = 32'h5be00000;
      20952: inst = 32'h244c8000;
      20953: inst = 32'h24428800;
      20954: inst = 32'h8620000;
      20955: inst = 32'h2a0e0004;
      20956: inst = 32'h294f0001;
      20957: inst = 32'h11200000;
      20958: inst = 32'hd2051e2;
      20959: inst = 32'h13e00000;
      20960: inst = 32'hfe0a9ea;
      20961: inst = 32'h5be00000;
      20962: inst = 32'h244c8000;
      20963: inst = 32'h24428800;
      20964: inst = 32'h8620000;
      20965: inst = 32'h2a0e0005;
      20966: inst = 32'h294f0001;
      20967: inst = 32'h11200000;
      20968: inst = 32'hd2051ec;
      20969: inst = 32'h13e00000;
      20970: inst = 32'hfe0a9ea;
      20971: inst = 32'h5be00000;
      20972: inst = 32'h244c8000;
      20973: inst = 32'h24428800;
      20974: inst = 32'h8620000;
      20975: inst = 32'h2a0e0006;
      20976: inst = 32'h294f0001;
      20977: inst = 32'h11200000;
      20978: inst = 32'hd2051f6;
      20979: inst = 32'h13e00000;
      20980: inst = 32'hfe0a9ea;
      20981: inst = 32'h5be00000;
      20982: inst = 32'h244c8000;
      20983: inst = 32'h24428800;
      20984: inst = 32'h8620000;
      20985: inst = 32'h2a0e0007;
      20986: inst = 32'h294f0001;
      20987: inst = 32'h11200000;
      20988: inst = 32'hd205200;
      20989: inst = 32'h13e00000;
      20990: inst = 32'hfe0a9ea;
      20991: inst = 32'h5be00000;
      20992: inst = 32'h244c8000;
      20993: inst = 32'h24428800;
      20994: inst = 32'h8620000;
      20995: inst = 32'h2a0e0008;
      20996: inst = 32'h294f0001;
      20997: inst = 32'h11200000;
      20998: inst = 32'hd20520a;
      20999: inst = 32'h13e00000;
      21000: inst = 32'hfe0a9ea;
      21001: inst = 32'h5be00000;
      21002: inst = 32'h244c8000;
      21003: inst = 32'h24428800;
      21004: inst = 32'h8620000;
      21005: inst = 32'h2a0e0009;
      21006: inst = 32'h294f0001;
      21007: inst = 32'h11200000;
      21008: inst = 32'hd205214;
      21009: inst = 32'h13e00000;
      21010: inst = 32'hfe0a9ea;
      21011: inst = 32'h5be00000;
      21012: inst = 32'h244c8000;
      21013: inst = 32'h24428800;
      21014: inst = 32'h8620000;
      21015: inst = 32'h2a0e0000;
      21016: inst = 32'h294f0002;
      21017: inst = 32'h11200000;
      21018: inst = 32'hd20521e;
      21019: inst = 32'h13e00000;
      21020: inst = 32'hfe0a9ea;
      21021: inst = 32'h5be00000;
      21022: inst = 32'h244c8000;
      21023: inst = 32'h24428800;
      21024: inst = 32'h8620000;
      21025: inst = 32'h2a0e0009;
      21026: inst = 32'h294f0002;
      21027: inst = 32'h11200000;
      21028: inst = 32'hd205228;
      21029: inst = 32'h13e00000;
      21030: inst = 32'hfe0a9ea;
      21031: inst = 32'h5be00000;
      21032: inst = 32'h244c8000;
      21033: inst = 32'h24428800;
      21034: inst = 32'h8620000;
      21035: inst = 32'h2a0e0000;
      21036: inst = 32'h294f0003;
      21037: inst = 32'h11200000;
      21038: inst = 32'hd205232;
      21039: inst = 32'h13e00000;
      21040: inst = 32'hfe0a9ea;
      21041: inst = 32'h5be00000;
      21042: inst = 32'h244c8000;
      21043: inst = 32'h24428800;
      21044: inst = 32'h8620000;
      21045: inst = 32'h2a0e0002;
      21046: inst = 32'h294f0003;
      21047: inst = 32'h11200000;
      21048: inst = 32'hd20523c;
      21049: inst = 32'h13e00000;
      21050: inst = 32'hfe0a9ea;
      21051: inst = 32'h5be00000;
      21052: inst = 32'h244c8000;
      21053: inst = 32'h24428800;
      21054: inst = 32'h8620000;
      21055: inst = 32'h2a0e0007;
      21056: inst = 32'h294f0003;
      21057: inst = 32'h11200000;
      21058: inst = 32'hd205246;
      21059: inst = 32'h13e00000;
      21060: inst = 32'hfe0a9ea;
      21061: inst = 32'h5be00000;
      21062: inst = 32'h244c8000;
      21063: inst = 32'h24428800;
      21064: inst = 32'h8620000;
      21065: inst = 32'h2a0e0009;
      21066: inst = 32'h294f0003;
      21067: inst = 32'h11200000;
      21068: inst = 32'hd205250;
      21069: inst = 32'h13e00000;
      21070: inst = 32'hfe0a9ea;
      21071: inst = 32'h5be00000;
      21072: inst = 32'h244c8000;
      21073: inst = 32'h24428800;
      21074: inst = 32'h8620000;
      21075: inst = 32'h2a0e0000;
      21076: inst = 32'h294f0004;
      21077: inst = 32'h11200000;
      21078: inst = 32'hd20525a;
      21079: inst = 32'h13e00000;
      21080: inst = 32'hfe0a9ea;
      21081: inst = 32'h5be00000;
      21082: inst = 32'h244c8000;
      21083: inst = 32'h24428800;
      21084: inst = 32'h8620000;
      21085: inst = 32'h2a0e0002;
      21086: inst = 32'h294f0004;
      21087: inst = 32'h11200000;
      21088: inst = 32'hd205264;
      21089: inst = 32'h13e00000;
      21090: inst = 32'hfe0a9ea;
      21091: inst = 32'h5be00000;
      21092: inst = 32'h244c8000;
      21093: inst = 32'h24428800;
      21094: inst = 32'h8620000;
      21095: inst = 32'h2a0e0007;
      21096: inst = 32'h294f0004;
      21097: inst = 32'h11200000;
      21098: inst = 32'hd20526e;
      21099: inst = 32'h13e00000;
      21100: inst = 32'hfe0a9ea;
      21101: inst = 32'h5be00000;
      21102: inst = 32'h244c8000;
      21103: inst = 32'h24428800;
      21104: inst = 32'h8620000;
      21105: inst = 32'h2a0e0009;
      21106: inst = 32'h294f0004;
      21107: inst = 32'h11200000;
      21108: inst = 32'hd205278;
      21109: inst = 32'h13e00000;
      21110: inst = 32'hfe0a9ea;
      21111: inst = 32'h5be00000;
      21112: inst = 32'h244c8000;
      21113: inst = 32'h24428800;
      21114: inst = 32'h8620000;
      21115: inst = 32'h2a0e0000;
      21116: inst = 32'h294f0005;
      21117: inst = 32'h11200000;
      21118: inst = 32'hd205282;
      21119: inst = 32'h13e00000;
      21120: inst = 32'hfe0a9ea;
      21121: inst = 32'h5be00000;
      21122: inst = 32'h244c8000;
      21123: inst = 32'h24428800;
      21124: inst = 32'h8620000;
      21125: inst = 32'h2a0e0009;
      21126: inst = 32'h294f0005;
      21127: inst = 32'h11200000;
      21128: inst = 32'hd20528c;
      21129: inst = 32'h13e00000;
      21130: inst = 32'hfe0a9ea;
      21131: inst = 32'h5be00000;
      21132: inst = 32'h244c8000;
      21133: inst = 32'h24428800;
      21134: inst = 32'h8620000;
      21135: inst = 32'h2a0e0000;
      21136: inst = 32'h294f0006;
      21137: inst = 32'h11200000;
      21138: inst = 32'hd205296;
      21139: inst = 32'h13e00000;
      21140: inst = 32'hfe0a9ea;
      21141: inst = 32'h5be00000;
      21142: inst = 32'h244c8000;
      21143: inst = 32'h24428800;
      21144: inst = 32'h8620000;
      21145: inst = 32'h2a0e0009;
      21146: inst = 32'h294f0006;
      21147: inst = 32'h11200000;
      21148: inst = 32'hd2052a0;
      21149: inst = 32'h13e00000;
      21150: inst = 32'hfe0a9ea;
      21151: inst = 32'h5be00000;
      21152: inst = 32'h244c8000;
      21153: inst = 32'h24428800;
      21154: inst = 32'h8620000;
      21155: inst = 32'hc60f4ce;
      21156: inst = 32'h2a0e0001;
      21157: inst = 32'h294f0002;
      21158: inst = 32'h11200000;
      21159: inst = 32'hd2052ab;
      21160: inst = 32'h13e00000;
      21161: inst = 32'hfe0a9ea;
      21162: inst = 32'h5be00000;
      21163: inst = 32'h244c8000;
      21164: inst = 32'h24428800;
      21165: inst = 32'h8620000;
      21166: inst = 32'h2a0e0002;
      21167: inst = 32'h294f0002;
      21168: inst = 32'h11200000;
      21169: inst = 32'hd2052b5;
      21170: inst = 32'h13e00000;
      21171: inst = 32'hfe0a9ea;
      21172: inst = 32'h5be00000;
      21173: inst = 32'h244c8000;
      21174: inst = 32'h24428800;
      21175: inst = 32'h8620000;
      21176: inst = 32'h2a0e0003;
      21177: inst = 32'h294f0002;
      21178: inst = 32'h11200000;
      21179: inst = 32'hd2052bf;
      21180: inst = 32'h13e00000;
      21181: inst = 32'hfe0a9ea;
      21182: inst = 32'h5be00000;
      21183: inst = 32'h244c8000;
      21184: inst = 32'h24428800;
      21185: inst = 32'h8620000;
      21186: inst = 32'h2a0e0004;
      21187: inst = 32'h294f0002;
      21188: inst = 32'h11200000;
      21189: inst = 32'hd2052c9;
      21190: inst = 32'h13e00000;
      21191: inst = 32'hfe0a9ea;
      21192: inst = 32'h5be00000;
      21193: inst = 32'h244c8000;
      21194: inst = 32'h24428800;
      21195: inst = 32'h8620000;
      21196: inst = 32'h2a0e0005;
      21197: inst = 32'h294f0002;
      21198: inst = 32'h11200000;
      21199: inst = 32'hd2052d3;
      21200: inst = 32'h13e00000;
      21201: inst = 32'hfe0a9ea;
      21202: inst = 32'h5be00000;
      21203: inst = 32'h244c8000;
      21204: inst = 32'h24428800;
      21205: inst = 32'h8620000;
      21206: inst = 32'h2a0e0006;
      21207: inst = 32'h294f0002;
      21208: inst = 32'h11200000;
      21209: inst = 32'hd2052dd;
      21210: inst = 32'h13e00000;
      21211: inst = 32'hfe0a9ea;
      21212: inst = 32'h5be00000;
      21213: inst = 32'h244c8000;
      21214: inst = 32'h24428800;
      21215: inst = 32'h8620000;
      21216: inst = 32'h2a0e0007;
      21217: inst = 32'h294f0002;
      21218: inst = 32'h11200000;
      21219: inst = 32'hd2052e7;
      21220: inst = 32'h13e00000;
      21221: inst = 32'hfe0a9ea;
      21222: inst = 32'h5be00000;
      21223: inst = 32'h244c8000;
      21224: inst = 32'h24428800;
      21225: inst = 32'h8620000;
      21226: inst = 32'h2a0e0008;
      21227: inst = 32'h294f0002;
      21228: inst = 32'h11200000;
      21229: inst = 32'hd2052f1;
      21230: inst = 32'h13e00000;
      21231: inst = 32'hfe0a9ea;
      21232: inst = 32'h5be00000;
      21233: inst = 32'h244c8000;
      21234: inst = 32'h24428800;
      21235: inst = 32'h8620000;
      21236: inst = 32'h2a0e0001;
      21237: inst = 32'h294f0003;
      21238: inst = 32'h11200000;
      21239: inst = 32'hd2052fb;
      21240: inst = 32'h13e00000;
      21241: inst = 32'hfe0a9ea;
      21242: inst = 32'h5be00000;
      21243: inst = 32'h244c8000;
      21244: inst = 32'h24428800;
      21245: inst = 32'h8620000;
      21246: inst = 32'h2a0e0003;
      21247: inst = 32'h294f0003;
      21248: inst = 32'h11200000;
      21249: inst = 32'hd205305;
      21250: inst = 32'h13e00000;
      21251: inst = 32'hfe0a9ea;
      21252: inst = 32'h5be00000;
      21253: inst = 32'h244c8000;
      21254: inst = 32'h24428800;
      21255: inst = 32'h8620000;
      21256: inst = 32'h2a0e0004;
      21257: inst = 32'h294f0003;
      21258: inst = 32'h11200000;
      21259: inst = 32'hd20530f;
      21260: inst = 32'h13e00000;
      21261: inst = 32'hfe0a9ea;
      21262: inst = 32'h5be00000;
      21263: inst = 32'h244c8000;
      21264: inst = 32'h24428800;
      21265: inst = 32'h8620000;
      21266: inst = 32'h2a0e0005;
      21267: inst = 32'h294f0003;
      21268: inst = 32'h11200000;
      21269: inst = 32'hd205319;
      21270: inst = 32'h13e00000;
      21271: inst = 32'hfe0a9ea;
      21272: inst = 32'h5be00000;
      21273: inst = 32'h244c8000;
      21274: inst = 32'h24428800;
      21275: inst = 32'h8620000;
      21276: inst = 32'h2a0e0006;
      21277: inst = 32'h294f0003;
      21278: inst = 32'h11200000;
      21279: inst = 32'hd205323;
      21280: inst = 32'h13e00000;
      21281: inst = 32'hfe0a9ea;
      21282: inst = 32'h5be00000;
      21283: inst = 32'h244c8000;
      21284: inst = 32'h24428800;
      21285: inst = 32'h8620000;
      21286: inst = 32'h2a0e0008;
      21287: inst = 32'h294f0003;
      21288: inst = 32'h11200000;
      21289: inst = 32'hd20532d;
      21290: inst = 32'h13e00000;
      21291: inst = 32'hfe0a9ea;
      21292: inst = 32'h5be00000;
      21293: inst = 32'h244c8000;
      21294: inst = 32'h24428800;
      21295: inst = 32'h8620000;
      21296: inst = 32'h2a0e0001;
      21297: inst = 32'h294f0004;
      21298: inst = 32'h11200000;
      21299: inst = 32'hd205337;
      21300: inst = 32'h13e00000;
      21301: inst = 32'hfe0a9ea;
      21302: inst = 32'h5be00000;
      21303: inst = 32'h244c8000;
      21304: inst = 32'h24428800;
      21305: inst = 32'h8620000;
      21306: inst = 32'h2a0e0003;
      21307: inst = 32'h294f0004;
      21308: inst = 32'h11200000;
      21309: inst = 32'hd205341;
      21310: inst = 32'h13e00000;
      21311: inst = 32'hfe0a9ea;
      21312: inst = 32'h5be00000;
      21313: inst = 32'h244c8000;
      21314: inst = 32'h24428800;
      21315: inst = 32'h8620000;
      21316: inst = 32'h2a0e0004;
      21317: inst = 32'h294f0004;
      21318: inst = 32'h11200000;
      21319: inst = 32'hd20534b;
      21320: inst = 32'h13e00000;
      21321: inst = 32'hfe0a9ea;
      21322: inst = 32'h5be00000;
      21323: inst = 32'h244c8000;
      21324: inst = 32'h24428800;
      21325: inst = 32'h8620000;
      21326: inst = 32'h2a0e0005;
      21327: inst = 32'h294f0004;
      21328: inst = 32'h11200000;
      21329: inst = 32'hd205355;
      21330: inst = 32'h13e00000;
      21331: inst = 32'hfe0a9ea;
      21332: inst = 32'h5be00000;
      21333: inst = 32'h244c8000;
      21334: inst = 32'h24428800;
      21335: inst = 32'h8620000;
      21336: inst = 32'h2a0e0006;
      21337: inst = 32'h294f0004;
      21338: inst = 32'h11200000;
      21339: inst = 32'hd20535f;
      21340: inst = 32'h13e00000;
      21341: inst = 32'hfe0a9ea;
      21342: inst = 32'h5be00000;
      21343: inst = 32'h244c8000;
      21344: inst = 32'h24428800;
      21345: inst = 32'h8620000;
      21346: inst = 32'h2a0e0008;
      21347: inst = 32'h294f0004;
      21348: inst = 32'h11200000;
      21349: inst = 32'hd205369;
      21350: inst = 32'h13e00000;
      21351: inst = 32'hfe0a9ea;
      21352: inst = 32'h5be00000;
      21353: inst = 32'h244c8000;
      21354: inst = 32'h24428800;
      21355: inst = 32'h8620000;
      21356: inst = 32'h2a0e0001;
      21357: inst = 32'h294f0005;
      21358: inst = 32'h11200000;
      21359: inst = 32'hd205373;
      21360: inst = 32'h13e00000;
      21361: inst = 32'hfe0a9ea;
      21362: inst = 32'h5be00000;
      21363: inst = 32'h244c8000;
      21364: inst = 32'h24428800;
      21365: inst = 32'h8620000;
      21366: inst = 32'h2a0e0002;
      21367: inst = 32'h294f0005;
      21368: inst = 32'h11200000;
      21369: inst = 32'hd20537d;
      21370: inst = 32'h13e00000;
      21371: inst = 32'hfe0a9ea;
      21372: inst = 32'h5be00000;
      21373: inst = 32'h244c8000;
      21374: inst = 32'h24428800;
      21375: inst = 32'h8620000;
      21376: inst = 32'h2a0e0003;
      21377: inst = 32'h294f0005;
      21378: inst = 32'h11200000;
      21379: inst = 32'hd205387;
      21380: inst = 32'h13e00000;
      21381: inst = 32'hfe0a9ea;
      21382: inst = 32'h5be00000;
      21383: inst = 32'h244c8000;
      21384: inst = 32'h24428800;
      21385: inst = 32'h8620000;
      21386: inst = 32'h2a0e0004;
      21387: inst = 32'h294f0005;
      21388: inst = 32'h11200000;
      21389: inst = 32'hd205391;
      21390: inst = 32'h13e00000;
      21391: inst = 32'hfe0a9ea;
      21392: inst = 32'h5be00000;
      21393: inst = 32'h244c8000;
      21394: inst = 32'h24428800;
      21395: inst = 32'h8620000;
      21396: inst = 32'h2a0e0005;
      21397: inst = 32'h294f0005;
      21398: inst = 32'h11200000;
      21399: inst = 32'hd20539b;
      21400: inst = 32'h13e00000;
      21401: inst = 32'hfe0a9ea;
      21402: inst = 32'h5be00000;
      21403: inst = 32'h244c8000;
      21404: inst = 32'h24428800;
      21405: inst = 32'h8620000;
      21406: inst = 32'h2a0e0006;
      21407: inst = 32'h294f0005;
      21408: inst = 32'h11200000;
      21409: inst = 32'hd2053a5;
      21410: inst = 32'h13e00000;
      21411: inst = 32'hfe0a9ea;
      21412: inst = 32'h5be00000;
      21413: inst = 32'h244c8000;
      21414: inst = 32'h24428800;
      21415: inst = 32'h8620000;
      21416: inst = 32'h2a0e0007;
      21417: inst = 32'h294f0005;
      21418: inst = 32'h11200000;
      21419: inst = 32'hd2053af;
      21420: inst = 32'h13e00000;
      21421: inst = 32'hfe0a9ea;
      21422: inst = 32'h5be00000;
      21423: inst = 32'h244c8000;
      21424: inst = 32'h24428800;
      21425: inst = 32'h8620000;
      21426: inst = 32'h2a0e0008;
      21427: inst = 32'h294f0005;
      21428: inst = 32'h11200000;
      21429: inst = 32'hd2053b9;
      21430: inst = 32'h13e00000;
      21431: inst = 32'hfe0a9ea;
      21432: inst = 32'h5be00000;
      21433: inst = 32'h244c8000;
      21434: inst = 32'h24428800;
      21435: inst = 32'h8620000;
      21436: inst = 32'h2a0e0001;
      21437: inst = 32'h294f0006;
      21438: inst = 32'h11200000;
      21439: inst = 32'hd2053c3;
      21440: inst = 32'h13e00000;
      21441: inst = 32'hfe0a9ea;
      21442: inst = 32'h5be00000;
      21443: inst = 32'h244c8000;
      21444: inst = 32'h24428800;
      21445: inst = 32'h8620000;
      21446: inst = 32'h2a0e0002;
      21447: inst = 32'h294f0006;
      21448: inst = 32'h11200000;
      21449: inst = 32'hd2053cd;
      21450: inst = 32'h13e00000;
      21451: inst = 32'hfe0a9ea;
      21452: inst = 32'h5be00000;
      21453: inst = 32'h244c8000;
      21454: inst = 32'h24428800;
      21455: inst = 32'h8620000;
      21456: inst = 32'h2a0e0003;
      21457: inst = 32'h294f0006;
      21458: inst = 32'h11200000;
      21459: inst = 32'hd2053d7;
      21460: inst = 32'h13e00000;
      21461: inst = 32'hfe0a9ea;
      21462: inst = 32'h5be00000;
      21463: inst = 32'h244c8000;
      21464: inst = 32'h24428800;
      21465: inst = 32'h8620000;
      21466: inst = 32'h2a0e0004;
      21467: inst = 32'h294f0006;
      21468: inst = 32'h11200000;
      21469: inst = 32'hd2053e1;
      21470: inst = 32'h13e00000;
      21471: inst = 32'hfe0a9ea;
      21472: inst = 32'h5be00000;
      21473: inst = 32'h244c8000;
      21474: inst = 32'h24428800;
      21475: inst = 32'h8620000;
      21476: inst = 32'h2a0e0005;
      21477: inst = 32'h294f0006;
      21478: inst = 32'h11200000;
      21479: inst = 32'hd2053eb;
      21480: inst = 32'h13e00000;
      21481: inst = 32'hfe0a9ea;
      21482: inst = 32'h5be00000;
      21483: inst = 32'h244c8000;
      21484: inst = 32'h24428800;
      21485: inst = 32'h8620000;
      21486: inst = 32'h2a0e0006;
      21487: inst = 32'h294f0006;
      21488: inst = 32'h11200000;
      21489: inst = 32'hd2053f5;
      21490: inst = 32'h13e00000;
      21491: inst = 32'hfe0a9ea;
      21492: inst = 32'h5be00000;
      21493: inst = 32'h244c8000;
      21494: inst = 32'h24428800;
      21495: inst = 32'h8620000;
      21496: inst = 32'h2a0e0007;
      21497: inst = 32'h294f0006;
      21498: inst = 32'h11200000;
      21499: inst = 32'hd2053ff;
      21500: inst = 32'h13e00000;
      21501: inst = 32'hfe0a9ea;
      21502: inst = 32'h5be00000;
      21503: inst = 32'h244c8000;
      21504: inst = 32'h24428800;
      21505: inst = 32'h8620000;
      21506: inst = 32'h2a0e0008;
      21507: inst = 32'h294f0006;
      21508: inst = 32'h11200000;
      21509: inst = 32'hd205409;
      21510: inst = 32'h13e00000;
      21511: inst = 32'hfe0a9ea;
      21512: inst = 32'h5be00000;
      21513: inst = 32'h244c8000;
      21514: inst = 32'h24428800;
      21515: inst = 32'h8620000;
      21516: inst = 32'h2a0e0000;
      21517: inst = 32'h294f0008;
      21518: inst = 32'h11200000;
      21519: inst = 32'hd205413;
      21520: inst = 32'h13e00000;
      21521: inst = 32'hfe0a9ea;
      21522: inst = 32'h5be00000;
      21523: inst = 32'h244c8000;
      21524: inst = 32'h24428800;
      21525: inst = 32'h8620000;
      21526: inst = 32'h2a0e0001;
      21527: inst = 32'h294f0008;
      21528: inst = 32'h11200000;
      21529: inst = 32'hd20541d;
      21530: inst = 32'h13e00000;
      21531: inst = 32'hfe0a9ea;
      21532: inst = 32'h5be00000;
      21533: inst = 32'h244c8000;
      21534: inst = 32'h24428800;
      21535: inst = 32'h8620000;
      21536: inst = 32'h2a0e0008;
      21537: inst = 32'h294f0008;
      21538: inst = 32'h11200000;
      21539: inst = 32'hd205427;
      21540: inst = 32'h13e00000;
      21541: inst = 32'hfe0a9ea;
      21542: inst = 32'h5be00000;
      21543: inst = 32'h244c8000;
      21544: inst = 32'h24428800;
      21545: inst = 32'h8620000;
      21546: inst = 32'h2a0e0009;
      21547: inst = 32'h294f0008;
      21548: inst = 32'h11200000;
      21549: inst = 32'hd205431;
      21550: inst = 32'h13e00000;
      21551: inst = 32'hfe0a9ea;
      21552: inst = 32'h5be00000;
      21553: inst = 32'h244c8000;
      21554: inst = 32'h24428800;
      21555: inst = 32'h8620000;
      21556: inst = 32'h2a0e0003;
      21557: inst = 32'h294f000c;
      21558: inst = 32'h11200000;
      21559: inst = 32'hd20543b;
      21560: inst = 32'h13e00000;
      21561: inst = 32'hfe0a9ea;
      21562: inst = 32'h5be00000;
      21563: inst = 32'h244c8000;
      21564: inst = 32'h24428800;
      21565: inst = 32'h8620000;
      21566: inst = 32'h2a0e0006;
      21567: inst = 32'h294f000c;
      21568: inst = 32'h11200000;
      21569: inst = 32'hd205445;
      21570: inst = 32'h13e00000;
      21571: inst = 32'hfe0a9ea;
      21572: inst = 32'h5be00000;
      21573: inst = 32'h244c8000;
      21574: inst = 32'h24428800;
      21575: inst = 32'h8620000;
      21576: inst = 32'hc607800;
      21577: inst = 32'h2a0e0002;
      21578: inst = 32'h294f0007;
      21579: inst = 32'h11200000;
      21580: inst = 32'hd205450;
      21581: inst = 32'h13e00000;
      21582: inst = 32'hfe0a9ea;
      21583: inst = 32'h5be00000;
      21584: inst = 32'h244c8000;
      21585: inst = 32'h24428800;
      21586: inst = 32'h8620000;
      21587: inst = 32'h2a0e0003;
      21588: inst = 32'h294f0007;
      21589: inst = 32'h11200000;
      21590: inst = 32'hd20545a;
      21591: inst = 32'h13e00000;
      21592: inst = 32'hfe0a9ea;
      21593: inst = 32'h5be00000;
      21594: inst = 32'h244c8000;
      21595: inst = 32'h24428800;
      21596: inst = 32'h8620000;
      21597: inst = 32'h2a0e0006;
      21598: inst = 32'h294f0007;
      21599: inst = 32'h11200000;
      21600: inst = 32'hd205464;
      21601: inst = 32'h13e00000;
      21602: inst = 32'hfe0a9ea;
      21603: inst = 32'h5be00000;
      21604: inst = 32'h244c8000;
      21605: inst = 32'h24428800;
      21606: inst = 32'h8620000;
      21607: inst = 32'h2a0e0007;
      21608: inst = 32'h294f0007;
      21609: inst = 32'h11200000;
      21610: inst = 32'hd20546e;
      21611: inst = 32'h13e00000;
      21612: inst = 32'hfe0a9ea;
      21613: inst = 32'h5be00000;
      21614: inst = 32'h244c8000;
      21615: inst = 32'h24428800;
      21616: inst = 32'h8620000;
      21617: inst = 32'hc60a000;
      21618: inst = 32'h2a0e0004;
      21619: inst = 32'h294f0007;
      21620: inst = 32'h11200000;
      21621: inst = 32'hd205479;
      21622: inst = 32'h13e00000;
      21623: inst = 32'hfe0a9ea;
      21624: inst = 32'h5be00000;
      21625: inst = 32'h244c8000;
      21626: inst = 32'h24428800;
      21627: inst = 32'h8620000;
      21628: inst = 32'h2a0e0005;
      21629: inst = 32'h294f0007;
      21630: inst = 32'h11200000;
      21631: inst = 32'hd205483;
      21632: inst = 32'h13e00000;
      21633: inst = 32'hfe0a9ea;
      21634: inst = 32'h5be00000;
      21635: inst = 32'h244c8000;
      21636: inst = 32'h24428800;
      21637: inst = 32'h8620000;
      21638: inst = 32'h2a0e0002;
      21639: inst = 32'h294f0008;
      21640: inst = 32'h11200000;
      21641: inst = 32'hd20548d;
      21642: inst = 32'h13e00000;
      21643: inst = 32'hfe0a9ea;
      21644: inst = 32'h5be00000;
      21645: inst = 32'h244c8000;
      21646: inst = 32'h24428800;
      21647: inst = 32'h8620000;
      21648: inst = 32'h2a0e0003;
      21649: inst = 32'h294f0008;
      21650: inst = 32'h11200000;
      21651: inst = 32'hd205497;
      21652: inst = 32'h13e00000;
      21653: inst = 32'hfe0a9ea;
      21654: inst = 32'h5be00000;
      21655: inst = 32'h244c8000;
      21656: inst = 32'h24428800;
      21657: inst = 32'h8620000;
      21658: inst = 32'h2a0e0004;
      21659: inst = 32'h294f0008;
      21660: inst = 32'h11200000;
      21661: inst = 32'hd2054a1;
      21662: inst = 32'h13e00000;
      21663: inst = 32'hfe0a9ea;
      21664: inst = 32'h5be00000;
      21665: inst = 32'h244c8000;
      21666: inst = 32'h24428800;
      21667: inst = 32'h8620000;
      21668: inst = 32'h2a0e0005;
      21669: inst = 32'h294f0008;
      21670: inst = 32'h11200000;
      21671: inst = 32'hd2054ab;
      21672: inst = 32'h13e00000;
      21673: inst = 32'hfe0a9ea;
      21674: inst = 32'h5be00000;
      21675: inst = 32'h244c8000;
      21676: inst = 32'h24428800;
      21677: inst = 32'h8620000;
      21678: inst = 32'h2a0e0006;
      21679: inst = 32'h294f0008;
      21680: inst = 32'h11200000;
      21681: inst = 32'hd2054b5;
      21682: inst = 32'h13e00000;
      21683: inst = 32'hfe0a9ea;
      21684: inst = 32'h5be00000;
      21685: inst = 32'h244c8000;
      21686: inst = 32'h24428800;
      21687: inst = 32'h8620000;
      21688: inst = 32'h2a0e0007;
      21689: inst = 32'h294f0008;
      21690: inst = 32'h11200000;
      21691: inst = 32'hd2054bf;
      21692: inst = 32'h13e00000;
      21693: inst = 32'hfe0a9ea;
      21694: inst = 32'h5be00000;
      21695: inst = 32'h244c8000;
      21696: inst = 32'h24428800;
      21697: inst = 32'h8620000;
      21698: inst = 32'h2a0e0002;
      21699: inst = 32'h294f0009;
      21700: inst = 32'h11200000;
      21701: inst = 32'hd2054c9;
      21702: inst = 32'h13e00000;
      21703: inst = 32'hfe0a9ea;
      21704: inst = 32'h5be00000;
      21705: inst = 32'h244c8000;
      21706: inst = 32'h24428800;
      21707: inst = 32'h8620000;
      21708: inst = 32'h2a0e0003;
      21709: inst = 32'h294f0009;
      21710: inst = 32'h11200000;
      21711: inst = 32'hd2054d3;
      21712: inst = 32'h13e00000;
      21713: inst = 32'hfe0a9ea;
      21714: inst = 32'h5be00000;
      21715: inst = 32'h244c8000;
      21716: inst = 32'h24428800;
      21717: inst = 32'h8620000;
      21718: inst = 32'h2a0e0004;
      21719: inst = 32'h294f0009;
      21720: inst = 32'h11200000;
      21721: inst = 32'hd2054dd;
      21722: inst = 32'h13e00000;
      21723: inst = 32'hfe0a9ea;
      21724: inst = 32'h5be00000;
      21725: inst = 32'h244c8000;
      21726: inst = 32'h24428800;
      21727: inst = 32'h8620000;
      21728: inst = 32'h2a0e0005;
      21729: inst = 32'h294f0009;
      21730: inst = 32'h11200000;
      21731: inst = 32'hd2054e7;
      21732: inst = 32'h13e00000;
      21733: inst = 32'hfe0a9ea;
      21734: inst = 32'h5be00000;
      21735: inst = 32'h244c8000;
      21736: inst = 32'h24428800;
      21737: inst = 32'h8620000;
      21738: inst = 32'h2a0e0006;
      21739: inst = 32'h294f0009;
      21740: inst = 32'h11200000;
      21741: inst = 32'hd2054f1;
      21742: inst = 32'h13e00000;
      21743: inst = 32'hfe0a9ea;
      21744: inst = 32'h5be00000;
      21745: inst = 32'h244c8000;
      21746: inst = 32'h24428800;
      21747: inst = 32'h8620000;
      21748: inst = 32'h2a0e0007;
      21749: inst = 32'h294f0009;
      21750: inst = 32'h11200000;
      21751: inst = 32'hd2054fb;
      21752: inst = 32'h13e00000;
      21753: inst = 32'hfe0a9ea;
      21754: inst = 32'h5be00000;
      21755: inst = 32'h244c8000;
      21756: inst = 32'h24428800;
      21757: inst = 32'h8620000;
      21758: inst = 32'hc6010ac;
      21759: inst = 32'h2a0e0002;
      21760: inst = 32'h294f000a;
      21761: inst = 32'h11200000;
      21762: inst = 32'hd205506;
      21763: inst = 32'h13e00000;
      21764: inst = 32'hfe0a9ea;
      21765: inst = 32'h5be00000;
      21766: inst = 32'h244c8000;
      21767: inst = 32'h24428800;
      21768: inst = 32'h8620000;
      21769: inst = 32'h2a0e0003;
      21770: inst = 32'h294f000a;
      21771: inst = 32'h11200000;
      21772: inst = 32'hd205510;
      21773: inst = 32'h13e00000;
      21774: inst = 32'hfe0a9ea;
      21775: inst = 32'h5be00000;
      21776: inst = 32'h244c8000;
      21777: inst = 32'h24428800;
      21778: inst = 32'h8620000;
      21779: inst = 32'h2a0e0004;
      21780: inst = 32'h294f000a;
      21781: inst = 32'h11200000;
      21782: inst = 32'hd20551a;
      21783: inst = 32'h13e00000;
      21784: inst = 32'hfe0a9ea;
      21785: inst = 32'h5be00000;
      21786: inst = 32'h244c8000;
      21787: inst = 32'h24428800;
      21788: inst = 32'h8620000;
      21789: inst = 32'h2a0e0005;
      21790: inst = 32'h294f000a;
      21791: inst = 32'h11200000;
      21792: inst = 32'hd205524;
      21793: inst = 32'h13e00000;
      21794: inst = 32'hfe0a9ea;
      21795: inst = 32'h5be00000;
      21796: inst = 32'h244c8000;
      21797: inst = 32'h24428800;
      21798: inst = 32'h8620000;
      21799: inst = 32'h2a0e0006;
      21800: inst = 32'h294f000a;
      21801: inst = 32'h11200000;
      21802: inst = 32'hd20552e;
      21803: inst = 32'h13e00000;
      21804: inst = 32'hfe0a9ea;
      21805: inst = 32'h5be00000;
      21806: inst = 32'h244c8000;
      21807: inst = 32'h24428800;
      21808: inst = 32'h8620000;
      21809: inst = 32'h2a0e0007;
      21810: inst = 32'h294f000a;
      21811: inst = 32'h11200000;
      21812: inst = 32'hd205538;
      21813: inst = 32'h13e00000;
      21814: inst = 32'hfe0a9ea;
      21815: inst = 32'h5be00000;
      21816: inst = 32'h244c8000;
      21817: inst = 32'h24428800;
      21818: inst = 32'h8620000;
      21819: inst = 32'hc60d42c;
      21820: inst = 32'h2a0e0003;
      21821: inst = 32'h294f000b;
      21822: inst = 32'h11200000;
      21823: inst = 32'hd205543;
      21824: inst = 32'h13e00000;
      21825: inst = 32'hfe0a9ea;
      21826: inst = 32'h5be00000;
      21827: inst = 32'h244c8000;
      21828: inst = 32'h24428800;
      21829: inst = 32'h8620000;
      21830: inst = 32'h2a0e0006;
      21831: inst = 32'h294f000b;
      21832: inst = 32'h11200000;
      21833: inst = 32'hd20554d;
      21834: inst = 32'h13e00000;
      21835: inst = 32'hfe0a9ea;
      21836: inst = 32'h5be00000;
      21837: inst = 32'h244c8000;
      21838: inst = 32'h24428800;
      21839: inst = 32'h8620000;
      21840: inst = 32'h13e00000;
      21841: inst = 32'hfe060f7;
      21842: inst = 32'h5be00000;
      21843: inst = 32'hc6018c3;
      21844: inst = 32'h2a0e0000;
      21845: inst = 32'h294f0000;
      21846: inst = 32'h11200000;
      21847: inst = 32'hd20555b;
      21848: inst = 32'h13e00000;
      21849: inst = 32'hfe0a9ea;
      21850: inst = 32'h5be00000;
      21851: inst = 32'h244c8000;
      21852: inst = 32'h24428800;
      21853: inst = 32'h8620000;
      21854: inst = 32'h2a0e0001;
      21855: inst = 32'h294f0000;
      21856: inst = 32'h11200000;
      21857: inst = 32'hd205565;
      21858: inst = 32'h13e00000;
      21859: inst = 32'hfe0a9ea;
      21860: inst = 32'h5be00000;
      21861: inst = 32'h244c8000;
      21862: inst = 32'h24428800;
      21863: inst = 32'h8620000;
      21864: inst = 32'h2a0e0002;
      21865: inst = 32'h294f0000;
      21866: inst = 32'h11200000;
      21867: inst = 32'hd20556f;
      21868: inst = 32'h13e00000;
      21869: inst = 32'hfe0a9ea;
      21870: inst = 32'h5be00000;
      21871: inst = 32'h244c8000;
      21872: inst = 32'h24428800;
      21873: inst = 32'h8620000;
      21874: inst = 32'h2a0e0003;
      21875: inst = 32'h294f0000;
      21876: inst = 32'h11200000;
      21877: inst = 32'hd205579;
      21878: inst = 32'h13e00000;
      21879: inst = 32'hfe0a9ea;
      21880: inst = 32'h5be00000;
      21881: inst = 32'h244c8000;
      21882: inst = 32'h24428800;
      21883: inst = 32'h8620000;
      21884: inst = 32'h2a0e0004;
      21885: inst = 32'h294f0000;
      21886: inst = 32'h11200000;
      21887: inst = 32'hd205583;
      21888: inst = 32'h13e00000;
      21889: inst = 32'hfe0a9ea;
      21890: inst = 32'h5be00000;
      21891: inst = 32'h244c8000;
      21892: inst = 32'h24428800;
      21893: inst = 32'h8620000;
      21894: inst = 32'h2a0e0005;
      21895: inst = 32'h294f0000;
      21896: inst = 32'h11200000;
      21897: inst = 32'hd20558d;
      21898: inst = 32'h13e00000;
      21899: inst = 32'hfe0a9ea;
      21900: inst = 32'h5be00000;
      21901: inst = 32'h244c8000;
      21902: inst = 32'h24428800;
      21903: inst = 32'h8620000;
      21904: inst = 32'h2a0e0006;
      21905: inst = 32'h294f0000;
      21906: inst = 32'h11200000;
      21907: inst = 32'hd205597;
      21908: inst = 32'h13e00000;
      21909: inst = 32'hfe0a9ea;
      21910: inst = 32'h5be00000;
      21911: inst = 32'h244c8000;
      21912: inst = 32'h24428800;
      21913: inst = 32'h8620000;
      21914: inst = 32'h2a0e0007;
      21915: inst = 32'h294f0000;
      21916: inst = 32'h11200000;
      21917: inst = 32'hd2055a1;
      21918: inst = 32'h13e00000;
      21919: inst = 32'hfe0a9ea;
      21920: inst = 32'h5be00000;
      21921: inst = 32'h244c8000;
      21922: inst = 32'h24428800;
      21923: inst = 32'h8620000;
      21924: inst = 32'h2a0e0008;
      21925: inst = 32'h294f0000;
      21926: inst = 32'h11200000;
      21927: inst = 32'hd2055ab;
      21928: inst = 32'h13e00000;
      21929: inst = 32'hfe0a9ea;
      21930: inst = 32'h5be00000;
      21931: inst = 32'h244c8000;
      21932: inst = 32'h24428800;
      21933: inst = 32'h8620000;
      21934: inst = 32'h2a0e0009;
      21935: inst = 32'h294f0000;
      21936: inst = 32'h11200000;
      21937: inst = 32'hd2055b5;
      21938: inst = 32'h13e00000;
      21939: inst = 32'hfe0a9ea;
      21940: inst = 32'h5be00000;
      21941: inst = 32'h244c8000;
      21942: inst = 32'h24428800;
      21943: inst = 32'h8620000;
      21944: inst = 32'h2a0e0000;
      21945: inst = 32'h294f0001;
      21946: inst = 32'h11200000;
      21947: inst = 32'hd2055bf;
      21948: inst = 32'h13e00000;
      21949: inst = 32'hfe0a9ea;
      21950: inst = 32'h5be00000;
      21951: inst = 32'h244c8000;
      21952: inst = 32'h24428800;
      21953: inst = 32'h8620000;
      21954: inst = 32'h2a0e0001;
      21955: inst = 32'h294f0001;
      21956: inst = 32'h11200000;
      21957: inst = 32'hd2055c9;
      21958: inst = 32'h13e00000;
      21959: inst = 32'hfe0a9ea;
      21960: inst = 32'h5be00000;
      21961: inst = 32'h244c8000;
      21962: inst = 32'h24428800;
      21963: inst = 32'h8620000;
      21964: inst = 32'h2a0e0002;
      21965: inst = 32'h294f0001;
      21966: inst = 32'h11200000;
      21967: inst = 32'hd2055d3;
      21968: inst = 32'h13e00000;
      21969: inst = 32'hfe0a9ea;
      21970: inst = 32'h5be00000;
      21971: inst = 32'h244c8000;
      21972: inst = 32'h24428800;
      21973: inst = 32'h8620000;
      21974: inst = 32'h2a0e0003;
      21975: inst = 32'h294f0001;
      21976: inst = 32'h11200000;
      21977: inst = 32'hd2055dd;
      21978: inst = 32'h13e00000;
      21979: inst = 32'hfe0a9ea;
      21980: inst = 32'h5be00000;
      21981: inst = 32'h244c8000;
      21982: inst = 32'h24428800;
      21983: inst = 32'h8620000;
      21984: inst = 32'h2a0e0004;
      21985: inst = 32'h294f0001;
      21986: inst = 32'h11200000;
      21987: inst = 32'hd2055e7;
      21988: inst = 32'h13e00000;
      21989: inst = 32'hfe0a9ea;
      21990: inst = 32'h5be00000;
      21991: inst = 32'h244c8000;
      21992: inst = 32'h24428800;
      21993: inst = 32'h8620000;
      21994: inst = 32'h2a0e0005;
      21995: inst = 32'h294f0001;
      21996: inst = 32'h11200000;
      21997: inst = 32'hd2055f1;
      21998: inst = 32'h13e00000;
      21999: inst = 32'hfe0a9ea;
      22000: inst = 32'h5be00000;
      22001: inst = 32'h244c8000;
      22002: inst = 32'h24428800;
      22003: inst = 32'h8620000;
      22004: inst = 32'h2a0e0006;
      22005: inst = 32'h294f0001;
      22006: inst = 32'h11200000;
      22007: inst = 32'hd2055fb;
      22008: inst = 32'h13e00000;
      22009: inst = 32'hfe0a9ea;
      22010: inst = 32'h5be00000;
      22011: inst = 32'h244c8000;
      22012: inst = 32'h24428800;
      22013: inst = 32'h8620000;
      22014: inst = 32'h2a0e0007;
      22015: inst = 32'h294f0001;
      22016: inst = 32'h11200000;
      22017: inst = 32'hd205605;
      22018: inst = 32'h13e00000;
      22019: inst = 32'hfe0a9ea;
      22020: inst = 32'h5be00000;
      22021: inst = 32'h244c8000;
      22022: inst = 32'h24428800;
      22023: inst = 32'h8620000;
      22024: inst = 32'h2a0e0008;
      22025: inst = 32'h294f0001;
      22026: inst = 32'h11200000;
      22027: inst = 32'hd20560f;
      22028: inst = 32'h13e00000;
      22029: inst = 32'hfe0a9ea;
      22030: inst = 32'h5be00000;
      22031: inst = 32'h244c8000;
      22032: inst = 32'h24428800;
      22033: inst = 32'h8620000;
      22034: inst = 32'h2a0e0009;
      22035: inst = 32'h294f0001;
      22036: inst = 32'h11200000;
      22037: inst = 32'hd205619;
      22038: inst = 32'h13e00000;
      22039: inst = 32'hfe0a9ea;
      22040: inst = 32'h5be00000;
      22041: inst = 32'h244c8000;
      22042: inst = 32'h24428800;
      22043: inst = 32'h8620000;
      22044: inst = 32'h2a0e0000;
      22045: inst = 32'h294f0002;
      22046: inst = 32'h11200000;
      22047: inst = 32'hd205623;
      22048: inst = 32'h13e00000;
      22049: inst = 32'hfe0a9ea;
      22050: inst = 32'h5be00000;
      22051: inst = 32'h244c8000;
      22052: inst = 32'h24428800;
      22053: inst = 32'h8620000;
      22054: inst = 32'h2a0e0001;
      22055: inst = 32'h294f0002;
      22056: inst = 32'h11200000;
      22057: inst = 32'hd20562d;
      22058: inst = 32'h13e00000;
      22059: inst = 32'hfe0a9ea;
      22060: inst = 32'h5be00000;
      22061: inst = 32'h244c8000;
      22062: inst = 32'h24428800;
      22063: inst = 32'h8620000;
      22064: inst = 32'h2a0e0002;
      22065: inst = 32'h294f0002;
      22066: inst = 32'h11200000;
      22067: inst = 32'hd205637;
      22068: inst = 32'h13e00000;
      22069: inst = 32'hfe0a9ea;
      22070: inst = 32'h5be00000;
      22071: inst = 32'h244c8000;
      22072: inst = 32'h24428800;
      22073: inst = 32'h8620000;
      22074: inst = 32'h2a0e0003;
      22075: inst = 32'h294f0002;
      22076: inst = 32'h11200000;
      22077: inst = 32'hd205641;
      22078: inst = 32'h13e00000;
      22079: inst = 32'hfe0a9ea;
      22080: inst = 32'h5be00000;
      22081: inst = 32'h244c8000;
      22082: inst = 32'h24428800;
      22083: inst = 32'h8620000;
      22084: inst = 32'h2a0e0004;
      22085: inst = 32'h294f0002;
      22086: inst = 32'h11200000;
      22087: inst = 32'hd20564b;
      22088: inst = 32'h13e00000;
      22089: inst = 32'hfe0a9ea;
      22090: inst = 32'h5be00000;
      22091: inst = 32'h244c8000;
      22092: inst = 32'h24428800;
      22093: inst = 32'h8620000;
      22094: inst = 32'h2a0e0005;
      22095: inst = 32'h294f0002;
      22096: inst = 32'h11200000;
      22097: inst = 32'hd205655;
      22098: inst = 32'h13e00000;
      22099: inst = 32'hfe0a9ea;
      22100: inst = 32'h5be00000;
      22101: inst = 32'h244c8000;
      22102: inst = 32'h24428800;
      22103: inst = 32'h8620000;
      22104: inst = 32'h2a0e0006;
      22105: inst = 32'h294f0002;
      22106: inst = 32'h11200000;
      22107: inst = 32'hd20565f;
      22108: inst = 32'h13e00000;
      22109: inst = 32'hfe0a9ea;
      22110: inst = 32'h5be00000;
      22111: inst = 32'h244c8000;
      22112: inst = 32'h24428800;
      22113: inst = 32'h8620000;
      22114: inst = 32'h2a0e0007;
      22115: inst = 32'h294f0002;
      22116: inst = 32'h11200000;
      22117: inst = 32'hd205669;
      22118: inst = 32'h13e00000;
      22119: inst = 32'hfe0a9ea;
      22120: inst = 32'h5be00000;
      22121: inst = 32'h244c8000;
      22122: inst = 32'h24428800;
      22123: inst = 32'h8620000;
      22124: inst = 32'h2a0e0008;
      22125: inst = 32'h294f0002;
      22126: inst = 32'h11200000;
      22127: inst = 32'hd205673;
      22128: inst = 32'h13e00000;
      22129: inst = 32'hfe0a9ea;
      22130: inst = 32'h5be00000;
      22131: inst = 32'h244c8000;
      22132: inst = 32'h24428800;
      22133: inst = 32'h8620000;
      22134: inst = 32'h2a0e0009;
      22135: inst = 32'h294f0002;
      22136: inst = 32'h11200000;
      22137: inst = 32'hd20567d;
      22138: inst = 32'h13e00000;
      22139: inst = 32'hfe0a9ea;
      22140: inst = 32'h5be00000;
      22141: inst = 32'h244c8000;
      22142: inst = 32'h24428800;
      22143: inst = 32'h8620000;
      22144: inst = 32'h2a0e0000;
      22145: inst = 32'h294f0003;
      22146: inst = 32'h11200000;
      22147: inst = 32'hd205687;
      22148: inst = 32'h13e00000;
      22149: inst = 32'hfe0a9ea;
      22150: inst = 32'h5be00000;
      22151: inst = 32'h244c8000;
      22152: inst = 32'h24428800;
      22153: inst = 32'h8620000;
      22154: inst = 32'h2a0e0001;
      22155: inst = 32'h294f0003;
      22156: inst = 32'h11200000;
      22157: inst = 32'hd205691;
      22158: inst = 32'h13e00000;
      22159: inst = 32'hfe0a9ea;
      22160: inst = 32'h5be00000;
      22161: inst = 32'h244c8000;
      22162: inst = 32'h24428800;
      22163: inst = 32'h8620000;
      22164: inst = 32'h2a0e0002;
      22165: inst = 32'h294f0003;
      22166: inst = 32'h11200000;
      22167: inst = 32'hd20569b;
      22168: inst = 32'h13e00000;
      22169: inst = 32'hfe0a9ea;
      22170: inst = 32'h5be00000;
      22171: inst = 32'h244c8000;
      22172: inst = 32'h24428800;
      22173: inst = 32'h8620000;
      22174: inst = 32'h2a0e0003;
      22175: inst = 32'h294f0003;
      22176: inst = 32'h11200000;
      22177: inst = 32'hd2056a5;
      22178: inst = 32'h13e00000;
      22179: inst = 32'hfe0a9ea;
      22180: inst = 32'h5be00000;
      22181: inst = 32'h244c8000;
      22182: inst = 32'h24428800;
      22183: inst = 32'h8620000;
      22184: inst = 32'h2a0e0004;
      22185: inst = 32'h294f0003;
      22186: inst = 32'h11200000;
      22187: inst = 32'hd2056af;
      22188: inst = 32'h13e00000;
      22189: inst = 32'hfe0a9ea;
      22190: inst = 32'h5be00000;
      22191: inst = 32'h244c8000;
      22192: inst = 32'h24428800;
      22193: inst = 32'h8620000;
      22194: inst = 32'h2a0e0005;
      22195: inst = 32'h294f0003;
      22196: inst = 32'h11200000;
      22197: inst = 32'hd2056b9;
      22198: inst = 32'h13e00000;
      22199: inst = 32'hfe0a9ea;
      22200: inst = 32'h5be00000;
      22201: inst = 32'h244c8000;
      22202: inst = 32'h24428800;
      22203: inst = 32'h8620000;
      22204: inst = 32'h2a0e0006;
      22205: inst = 32'h294f0003;
      22206: inst = 32'h11200000;
      22207: inst = 32'hd2056c3;
      22208: inst = 32'h13e00000;
      22209: inst = 32'hfe0a9ea;
      22210: inst = 32'h5be00000;
      22211: inst = 32'h244c8000;
      22212: inst = 32'h24428800;
      22213: inst = 32'h8620000;
      22214: inst = 32'h2a0e0007;
      22215: inst = 32'h294f0003;
      22216: inst = 32'h11200000;
      22217: inst = 32'hd2056cd;
      22218: inst = 32'h13e00000;
      22219: inst = 32'hfe0a9ea;
      22220: inst = 32'h5be00000;
      22221: inst = 32'h244c8000;
      22222: inst = 32'h24428800;
      22223: inst = 32'h8620000;
      22224: inst = 32'h2a0e0008;
      22225: inst = 32'h294f0003;
      22226: inst = 32'h11200000;
      22227: inst = 32'hd2056d7;
      22228: inst = 32'h13e00000;
      22229: inst = 32'hfe0a9ea;
      22230: inst = 32'h5be00000;
      22231: inst = 32'h244c8000;
      22232: inst = 32'h24428800;
      22233: inst = 32'h8620000;
      22234: inst = 32'h2a0e0009;
      22235: inst = 32'h294f0003;
      22236: inst = 32'h11200000;
      22237: inst = 32'hd2056e1;
      22238: inst = 32'h13e00000;
      22239: inst = 32'hfe0a9ea;
      22240: inst = 32'h5be00000;
      22241: inst = 32'h244c8000;
      22242: inst = 32'h24428800;
      22243: inst = 32'h8620000;
      22244: inst = 32'h2a0e0000;
      22245: inst = 32'h294f0004;
      22246: inst = 32'h11200000;
      22247: inst = 32'hd2056eb;
      22248: inst = 32'h13e00000;
      22249: inst = 32'hfe0a9ea;
      22250: inst = 32'h5be00000;
      22251: inst = 32'h244c8000;
      22252: inst = 32'h24428800;
      22253: inst = 32'h8620000;
      22254: inst = 32'h2a0e0001;
      22255: inst = 32'h294f0004;
      22256: inst = 32'h11200000;
      22257: inst = 32'hd2056f5;
      22258: inst = 32'h13e00000;
      22259: inst = 32'hfe0a9ea;
      22260: inst = 32'h5be00000;
      22261: inst = 32'h244c8000;
      22262: inst = 32'h24428800;
      22263: inst = 32'h8620000;
      22264: inst = 32'h2a0e0002;
      22265: inst = 32'h294f0004;
      22266: inst = 32'h11200000;
      22267: inst = 32'hd2056ff;
      22268: inst = 32'h13e00000;
      22269: inst = 32'hfe0a9ea;
      22270: inst = 32'h5be00000;
      22271: inst = 32'h244c8000;
      22272: inst = 32'h24428800;
      22273: inst = 32'h8620000;
      22274: inst = 32'h2a0e0003;
      22275: inst = 32'h294f0004;
      22276: inst = 32'h11200000;
      22277: inst = 32'hd205709;
      22278: inst = 32'h13e00000;
      22279: inst = 32'hfe0a9ea;
      22280: inst = 32'h5be00000;
      22281: inst = 32'h244c8000;
      22282: inst = 32'h24428800;
      22283: inst = 32'h8620000;
      22284: inst = 32'h2a0e0004;
      22285: inst = 32'h294f0004;
      22286: inst = 32'h11200000;
      22287: inst = 32'hd205713;
      22288: inst = 32'h13e00000;
      22289: inst = 32'hfe0a9ea;
      22290: inst = 32'h5be00000;
      22291: inst = 32'h244c8000;
      22292: inst = 32'h24428800;
      22293: inst = 32'h8620000;
      22294: inst = 32'h2a0e0005;
      22295: inst = 32'h294f0004;
      22296: inst = 32'h11200000;
      22297: inst = 32'hd20571d;
      22298: inst = 32'h13e00000;
      22299: inst = 32'hfe0a9ea;
      22300: inst = 32'h5be00000;
      22301: inst = 32'h244c8000;
      22302: inst = 32'h24428800;
      22303: inst = 32'h8620000;
      22304: inst = 32'h2a0e0006;
      22305: inst = 32'h294f0004;
      22306: inst = 32'h11200000;
      22307: inst = 32'hd205727;
      22308: inst = 32'h13e00000;
      22309: inst = 32'hfe0a9ea;
      22310: inst = 32'h5be00000;
      22311: inst = 32'h244c8000;
      22312: inst = 32'h24428800;
      22313: inst = 32'h8620000;
      22314: inst = 32'h2a0e0007;
      22315: inst = 32'h294f0004;
      22316: inst = 32'h11200000;
      22317: inst = 32'hd205731;
      22318: inst = 32'h13e00000;
      22319: inst = 32'hfe0a9ea;
      22320: inst = 32'h5be00000;
      22321: inst = 32'h244c8000;
      22322: inst = 32'h24428800;
      22323: inst = 32'h8620000;
      22324: inst = 32'h2a0e0008;
      22325: inst = 32'h294f0004;
      22326: inst = 32'h11200000;
      22327: inst = 32'hd20573b;
      22328: inst = 32'h13e00000;
      22329: inst = 32'hfe0a9ea;
      22330: inst = 32'h5be00000;
      22331: inst = 32'h244c8000;
      22332: inst = 32'h24428800;
      22333: inst = 32'h8620000;
      22334: inst = 32'h2a0e0009;
      22335: inst = 32'h294f0004;
      22336: inst = 32'h11200000;
      22337: inst = 32'hd205745;
      22338: inst = 32'h13e00000;
      22339: inst = 32'hfe0a9ea;
      22340: inst = 32'h5be00000;
      22341: inst = 32'h244c8000;
      22342: inst = 32'h24428800;
      22343: inst = 32'h8620000;
      22344: inst = 32'h2a0e0000;
      22345: inst = 32'h294f0005;
      22346: inst = 32'h11200000;
      22347: inst = 32'hd20574f;
      22348: inst = 32'h13e00000;
      22349: inst = 32'hfe0a9ea;
      22350: inst = 32'h5be00000;
      22351: inst = 32'h244c8000;
      22352: inst = 32'h24428800;
      22353: inst = 32'h8620000;
      22354: inst = 32'h2a0e0001;
      22355: inst = 32'h294f0005;
      22356: inst = 32'h11200000;
      22357: inst = 32'hd205759;
      22358: inst = 32'h13e00000;
      22359: inst = 32'hfe0a9ea;
      22360: inst = 32'h5be00000;
      22361: inst = 32'h244c8000;
      22362: inst = 32'h24428800;
      22363: inst = 32'h8620000;
      22364: inst = 32'h2a0e0002;
      22365: inst = 32'h294f0005;
      22366: inst = 32'h11200000;
      22367: inst = 32'hd205763;
      22368: inst = 32'h13e00000;
      22369: inst = 32'hfe0a9ea;
      22370: inst = 32'h5be00000;
      22371: inst = 32'h244c8000;
      22372: inst = 32'h24428800;
      22373: inst = 32'h8620000;
      22374: inst = 32'h2a0e0003;
      22375: inst = 32'h294f0005;
      22376: inst = 32'h11200000;
      22377: inst = 32'hd20576d;
      22378: inst = 32'h13e00000;
      22379: inst = 32'hfe0a9ea;
      22380: inst = 32'h5be00000;
      22381: inst = 32'h244c8000;
      22382: inst = 32'h24428800;
      22383: inst = 32'h8620000;
      22384: inst = 32'h2a0e0004;
      22385: inst = 32'h294f0005;
      22386: inst = 32'h11200000;
      22387: inst = 32'hd205777;
      22388: inst = 32'h13e00000;
      22389: inst = 32'hfe0a9ea;
      22390: inst = 32'h5be00000;
      22391: inst = 32'h244c8000;
      22392: inst = 32'h24428800;
      22393: inst = 32'h8620000;
      22394: inst = 32'h2a0e0005;
      22395: inst = 32'h294f0005;
      22396: inst = 32'h11200000;
      22397: inst = 32'hd205781;
      22398: inst = 32'h13e00000;
      22399: inst = 32'hfe0a9ea;
      22400: inst = 32'h5be00000;
      22401: inst = 32'h244c8000;
      22402: inst = 32'h24428800;
      22403: inst = 32'h8620000;
      22404: inst = 32'h2a0e0006;
      22405: inst = 32'h294f0005;
      22406: inst = 32'h11200000;
      22407: inst = 32'hd20578b;
      22408: inst = 32'h13e00000;
      22409: inst = 32'hfe0a9ea;
      22410: inst = 32'h5be00000;
      22411: inst = 32'h244c8000;
      22412: inst = 32'h24428800;
      22413: inst = 32'h8620000;
      22414: inst = 32'h2a0e0007;
      22415: inst = 32'h294f0005;
      22416: inst = 32'h11200000;
      22417: inst = 32'hd205795;
      22418: inst = 32'h13e00000;
      22419: inst = 32'hfe0a9ea;
      22420: inst = 32'h5be00000;
      22421: inst = 32'h244c8000;
      22422: inst = 32'h24428800;
      22423: inst = 32'h8620000;
      22424: inst = 32'h2a0e0008;
      22425: inst = 32'h294f0005;
      22426: inst = 32'h11200000;
      22427: inst = 32'hd20579f;
      22428: inst = 32'h13e00000;
      22429: inst = 32'hfe0a9ea;
      22430: inst = 32'h5be00000;
      22431: inst = 32'h244c8000;
      22432: inst = 32'h24428800;
      22433: inst = 32'h8620000;
      22434: inst = 32'h2a0e0009;
      22435: inst = 32'h294f0005;
      22436: inst = 32'h11200000;
      22437: inst = 32'hd2057a9;
      22438: inst = 32'h13e00000;
      22439: inst = 32'hfe0a9ea;
      22440: inst = 32'h5be00000;
      22441: inst = 32'h244c8000;
      22442: inst = 32'h24428800;
      22443: inst = 32'h8620000;
      22444: inst = 32'h2a0e0000;
      22445: inst = 32'h294f0006;
      22446: inst = 32'h11200000;
      22447: inst = 32'hd2057b3;
      22448: inst = 32'h13e00000;
      22449: inst = 32'hfe0a9ea;
      22450: inst = 32'h5be00000;
      22451: inst = 32'h244c8000;
      22452: inst = 32'h24428800;
      22453: inst = 32'h8620000;
      22454: inst = 32'h2a0e0001;
      22455: inst = 32'h294f0006;
      22456: inst = 32'h11200000;
      22457: inst = 32'hd2057bd;
      22458: inst = 32'h13e00000;
      22459: inst = 32'hfe0a9ea;
      22460: inst = 32'h5be00000;
      22461: inst = 32'h244c8000;
      22462: inst = 32'h24428800;
      22463: inst = 32'h8620000;
      22464: inst = 32'h2a0e0002;
      22465: inst = 32'h294f0006;
      22466: inst = 32'h11200000;
      22467: inst = 32'hd2057c7;
      22468: inst = 32'h13e00000;
      22469: inst = 32'hfe0a9ea;
      22470: inst = 32'h5be00000;
      22471: inst = 32'h244c8000;
      22472: inst = 32'h24428800;
      22473: inst = 32'h8620000;
      22474: inst = 32'h2a0e0003;
      22475: inst = 32'h294f0006;
      22476: inst = 32'h11200000;
      22477: inst = 32'hd2057d1;
      22478: inst = 32'h13e00000;
      22479: inst = 32'hfe0a9ea;
      22480: inst = 32'h5be00000;
      22481: inst = 32'h244c8000;
      22482: inst = 32'h24428800;
      22483: inst = 32'h8620000;
      22484: inst = 32'h2a0e0004;
      22485: inst = 32'h294f0006;
      22486: inst = 32'h11200000;
      22487: inst = 32'hd2057db;
      22488: inst = 32'h13e00000;
      22489: inst = 32'hfe0a9ea;
      22490: inst = 32'h5be00000;
      22491: inst = 32'h244c8000;
      22492: inst = 32'h24428800;
      22493: inst = 32'h8620000;
      22494: inst = 32'h2a0e0005;
      22495: inst = 32'h294f0006;
      22496: inst = 32'h11200000;
      22497: inst = 32'hd2057e5;
      22498: inst = 32'h13e00000;
      22499: inst = 32'hfe0a9ea;
      22500: inst = 32'h5be00000;
      22501: inst = 32'h244c8000;
      22502: inst = 32'h24428800;
      22503: inst = 32'h8620000;
      22504: inst = 32'h2a0e0006;
      22505: inst = 32'h294f0006;
      22506: inst = 32'h11200000;
      22507: inst = 32'hd2057ef;
      22508: inst = 32'h13e00000;
      22509: inst = 32'hfe0a9ea;
      22510: inst = 32'h5be00000;
      22511: inst = 32'h244c8000;
      22512: inst = 32'h24428800;
      22513: inst = 32'h8620000;
      22514: inst = 32'h2a0e0007;
      22515: inst = 32'h294f0006;
      22516: inst = 32'h11200000;
      22517: inst = 32'hd2057f9;
      22518: inst = 32'h13e00000;
      22519: inst = 32'hfe0a9ea;
      22520: inst = 32'h5be00000;
      22521: inst = 32'h244c8000;
      22522: inst = 32'h24428800;
      22523: inst = 32'h8620000;
      22524: inst = 32'h2a0e0008;
      22525: inst = 32'h294f0006;
      22526: inst = 32'h11200000;
      22527: inst = 32'hd205803;
      22528: inst = 32'h13e00000;
      22529: inst = 32'hfe0a9ea;
      22530: inst = 32'h5be00000;
      22531: inst = 32'h244c8000;
      22532: inst = 32'h24428800;
      22533: inst = 32'h8620000;
      22534: inst = 32'h2a0e0009;
      22535: inst = 32'h294f0006;
      22536: inst = 32'h11200000;
      22537: inst = 32'hd20580d;
      22538: inst = 32'h13e00000;
      22539: inst = 32'hfe0a9ea;
      22540: inst = 32'h5be00000;
      22541: inst = 32'h244c8000;
      22542: inst = 32'h24428800;
      22543: inst = 32'h8620000;
      22544: inst = 32'hc60f4ce;
      22545: inst = 32'h2a0e0001;
      22546: inst = 32'h294f0007;
      22547: inst = 32'h11200000;
      22548: inst = 32'hd205818;
      22549: inst = 32'h13e00000;
      22550: inst = 32'hfe0a9ea;
      22551: inst = 32'h5be00000;
      22552: inst = 32'h244c8000;
      22553: inst = 32'h24428800;
      22554: inst = 32'h8620000;
      22555: inst = 32'h2a0e0008;
      22556: inst = 32'h294f0007;
      22557: inst = 32'h11200000;
      22558: inst = 32'hd205822;
      22559: inst = 32'h13e00000;
      22560: inst = 32'hfe0a9ea;
      22561: inst = 32'h5be00000;
      22562: inst = 32'h244c8000;
      22563: inst = 32'h24428800;
      22564: inst = 32'h8620000;
      22565: inst = 32'h2a0e0001;
      22566: inst = 32'h294f0008;
      22567: inst = 32'h11200000;
      22568: inst = 32'hd20582c;
      22569: inst = 32'h13e00000;
      22570: inst = 32'hfe0a9ea;
      22571: inst = 32'h5be00000;
      22572: inst = 32'h244c8000;
      22573: inst = 32'h24428800;
      22574: inst = 32'h8620000;
      22575: inst = 32'h2a0e0008;
      22576: inst = 32'h294f0008;
      22577: inst = 32'h11200000;
      22578: inst = 32'hd205836;
      22579: inst = 32'h13e00000;
      22580: inst = 32'hfe0a9ea;
      22581: inst = 32'h5be00000;
      22582: inst = 32'h244c8000;
      22583: inst = 32'h24428800;
      22584: inst = 32'h8620000;
      22585: inst = 32'hc607841;
      22586: inst = 32'h2a0e0002;
      22587: inst = 32'h294f0007;
      22588: inst = 32'h11200000;
      22589: inst = 32'hd205841;
      22590: inst = 32'h13e00000;
      22591: inst = 32'hfe0a9ea;
      22592: inst = 32'h5be00000;
      22593: inst = 32'h244c8000;
      22594: inst = 32'h24428800;
      22595: inst = 32'h8620000;
      22596: inst = 32'h2a0e0003;
      22597: inst = 32'h294f0007;
      22598: inst = 32'h11200000;
      22599: inst = 32'hd20584b;
      22600: inst = 32'h13e00000;
      22601: inst = 32'hfe0a9ea;
      22602: inst = 32'h5be00000;
      22603: inst = 32'h244c8000;
      22604: inst = 32'h24428800;
      22605: inst = 32'h8620000;
      22606: inst = 32'h2a0e0004;
      22607: inst = 32'h294f0007;
      22608: inst = 32'h11200000;
      22609: inst = 32'hd205855;
      22610: inst = 32'h13e00000;
      22611: inst = 32'hfe0a9ea;
      22612: inst = 32'h5be00000;
      22613: inst = 32'h244c8000;
      22614: inst = 32'h24428800;
      22615: inst = 32'h8620000;
      22616: inst = 32'h2a0e0005;
      22617: inst = 32'h294f0007;
      22618: inst = 32'h11200000;
      22619: inst = 32'hd20585f;
      22620: inst = 32'h13e00000;
      22621: inst = 32'hfe0a9ea;
      22622: inst = 32'h5be00000;
      22623: inst = 32'h244c8000;
      22624: inst = 32'h24428800;
      22625: inst = 32'h8620000;
      22626: inst = 32'h2a0e0006;
      22627: inst = 32'h294f0007;
      22628: inst = 32'h11200000;
      22629: inst = 32'hd205869;
      22630: inst = 32'h13e00000;
      22631: inst = 32'hfe0a9ea;
      22632: inst = 32'h5be00000;
      22633: inst = 32'h244c8000;
      22634: inst = 32'h24428800;
      22635: inst = 32'h8620000;
      22636: inst = 32'h2a0e0007;
      22637: inst = 32'h294f0007;
      22638: inst = 32'h11200000;
      22639: inst = 32'hd205873;
      22640: inst = 32'h13e00000;
      22641: inst = 32'hfe0a9ea;
      22642: inst = 32'h5be00000;
      22643: inst = 32'h244c8000;
      22644: inst = 32'h24428800;
      22645: inst = 32'h8620000;
      22646: inst = 32'h2a0e0002;
      22647: inst = 32'h294f0008;
      22648: inst = 32'h11200000;
      22649: inst = 32'hd20587d;
      22650: inst = 32'h13e00000;
      22651: inst = 32'hfe0a9ea;
      22652: inst = 32'h5be00000;
      22653: inst = 32'h244c8000;
      22654: inst = 32'h24428800;
      22655: inst = 32'h8620000;
      22656: inst = 32'h2a0e0003;
      22657: inst = 32'h294f0008;
      22658: inst = 32'h11200000;
      22659: inst = 32'hd205887;
      22660: inst = 32'h13e00000;
      22661: inst = 32'hfe0a9ea;
      22662: inst = 32'h5be00000;
      22663: inst = 32'h244c8000;
      22664: inst = 32'h24428800;
      22665: inst = 32'h8620000;
      22666: inst = 32'h2a0e0004;
      22667: inst = 32'h294f0008;
      22668: inst = 32'h11200000;
      22669: inst = 32'hd205891;
      22670: inst = 32'h13e00000;
      22671: inst = 32'hfe0a9ea;
      22672: inst = 32'h5be00000;
      22673: inst = 32'h244c8000;
      22674: inst = 32'h24428800;
      22675: inst = 32'h8620000;
      22676: inst = 32'h2a0e0005;
      22677: inst = 32'h294f0008;
      22678: inst = 32'h11200000;
      22679: inst = 32'hd20589b;
      22680: inst = 32'h13e00000;
      22681: inst = 32'hfe0a9ea;
      22682: inst = 32'h5be00000;
      22683: inst = 32'h244c8000;
      22684: inst = 32'h24428800;
      22685: inst = 32'h8620000;
      22686: inst = 32'h2a0e0006;
      22687: inst = 32'h294f0008;
      22688: inst = 32'h11200000;
      22689: inst = 32'hd2058a5;
      22690: inst = 32'h13e00000;
      22691: inst = 32'hfe0a9ea;
      22692: inst = 32'h5be00000;
      22693: inst = 32'h244c8000;
      22694: inst = 32'h24428800;
      22695: inst = 32'h8620000;
      22696: inst = 32'h2a0e0007;
      22697: inst = 32'h294f0008;
      22698: inst = 32'h11200000;
      22699: inst = 32'hd2058af;
      22700: inst = 32'h13e00000;
      22701: inst = 32'hfe0a9ea;
      22702: inst = 32'h5be00000;
      22703: inst = 32'h244c8000;
      22704: inst = 32'h24428800;
      22705: inst = 32'h8620000;
      22706: inst = 32'h2a0e0002;
      22707: inst = 32'h294f0009;
      22708: inst = 32'h11200000;
      22709: inst = 32'hd2058b9;
      22710: inst = 32'h13e00000;
      22711: inst = 32'hfe0a9ea;
      22712: inst = 32'h5be00000;
      22713: inst = 32'h244c8000;
      22714: inst = 32'h24428800;
      22715: inst = 32'h8620000;
      22716: inst = 32'h2a0e0003;
      22717: inst = 32'h294f0009;
      22718: inst = 32'h11200000;
      22719: inst = 32'hd2058c3;
      22720: inst = 32'h13e00000;
      22721: inst = 32'hfe0a9ea;
      22722: inst = 32'h5be00000;
      22723: inst = 32'h244c8000;
      22724: inst = 32'h24428800;
      22725: inst = 32'h8620000;
      22726: inst = 32'h2a0e0004;
      22727: inst = 32'h294f0009;
      22728: inst = 32'h11200000;
      22729: inst = 32'hd2058cd;
      22730: inst = 32'h13e00000;
      22731: inst = 32'hfe0a9ea;
      22732: inst = 32'h5be00000;
      22733: inst = 32'h244c8000;
      22734: inst = 32'h24428800;
      22735: inst = 32'h8620000;
      22736: inst = 32'h2a0e0005;
      22737: inst = 32'h294f0009;
      22738: inst = 32'h11200000;
      22739: inst = 32'hd2058d7;
      22740: inst = 32'h13e00000;
      22741: inst = 32'hfe0a9ea;
      22742: inst = 32'h5be00000;
      22743: inst = 32'h244c8000;
      22744: inst = 32'h24428800;
      22745: inst = 32'h8620000;
      22746: inst = 32'h2a0e0006;
      22747: inst = 32'h294f0009;
      22748: inst = 32'h11200000;
      22749: inst = 32'hd2058e1;
      22750: inst = 32'h13e00000;
      22751: inst = 32'hfe0a9ea;
      22752: inst = 32'h5be00000;
      22753: inst = 32'h244c8000;
      22754: inst = 32'h24428800;
      22755: inst = 32'h8620000;
      22756: inst = 32'h2a0e0007;
      22757: inst = 32'h294f0009;
      22758: inst = 32'h11200000;
      22759: inst = 32'hd2058eb;
      22760: inst = 32'h13e00000;
      22761: inst = 32'hfe0a9ea;
      22762: inst = 32'h5be00000;
      22763: inst = 32'h244c8000;
      22764: inst = 32'h24428800;
      22765: inst = 32'h8620000;
      22766: inst = 32'hc6010ac;
      22767: inst = 32'h2a0e0002;
      22768: inst = 32'h294f000a;
      22769: inst = 32'h11200000;
      22770: inst = 32'hd2058f6;
      22771: inst = 32'h13e00000;
      22772: inst = 32'hfe0a9ea;
      22773: inst = 32'h5be00000;
      22774: inst = 32'h244c8000;
      22775: inst = 32'h24428800;
      22776: inst = 32'h8620000;
      22777: inst = 32'h2a0e0003;
      22778: inst = 32'h294f000a;
      22779: inst = 32'h11200000;
      22780: inst = 32'hd205900;
      22781: inst = 32'h13e00000;
      22782: inst = 32'hfe0a9ea;
      22783: inst = 32'h5be00000;
      22784: inst = 32'h244c8000;
      22785: inst = 32'h24428800;
      22786: inst = 32'h8620000;
      22787: inst = 32'h2a0e0004;
      22788: inst = 32'h294f000a;
      22789: inst = 32'h11200000;
      22790: inst = 32'hd20590a;
      22791: inst = 32'h13e00000;
      22792: inst = 32'hfe0a9ea;
      22793: inst = 32'h5be00000;
      22794: inst = 32'h244c8000;
      22795: inst = 32'h24428800;
      22796: inst = 32'h8620000;
      22797: inst = 32'h2a0e0005;
      22798: inst = 32'h294f000a;
      22799: inst = 32'h11200000;
      22800: inst = 32'hd205914;
      22801: inst = 32'h13e00000;
      22802: inst = 32'hfe0a9ea;
      22803: inst = 32'h5be00000;
      22804: inst = 32'h244c8000;
      22805: inst = 32'h24428800;
      22806: inst = 32'h8620000;
      22807: inst = 32'h2a0e0006;
      22808: inst = 32'h294f000a;
      22809: inst = 32'h11200000;
      22810: inst = 32'hd20591e;
      22811: inst = 32'h13e00000;
      22812: inst = 32'hfe0a9ea;
      22813: inst = 32'h5be00000;
      22814: inst = 32'h244c8000;
      22815: inst = 32'h24428800;
      22816: inst = 32'h8620000;
      22817: inst = 32'h2a0e0007;
      22818: inst = 32'h294f000a;
      22819: inst = 32'h11200000;
      22820: inst = 32'hd205928;
      22821: inst = 32'h13e00000;
      22822: inst = 32'hfe0a9ea;
      22823: inst = 32'h5be00000;
      22824: inst = 32'h244c8000;
      22825: inst = 32'h24428800;
      22826: inst = 32'h8620000;
      22827: inst = 32'hc60d42c;
      22828: inst = 32'h2a0e0003;
      22829: inst = 32'h294f000b;
      22830: inst = 32'h11200000;
      22831: inst = 32'hd205933;
      22832: inst = 32'h13e00000;
      22833: inst = 32'hfe0a9ea;
      22834: inst = 32'h5be00000;
      22835: inst = 32'h244c8000;
      22836: inst = 32'h24428800;
      22837: inst = 32'h8620000;
      22838: inst = 32'h2a0e0006;
      22839: inst = 32'h294f000b;
      22840: inst = 32'h11200000;
      22841: inst = 32'hd20593d;
      22842: inst = 32'h13e00000;
      22843: inst = 32'hfe0a9ea;
      22844: inst = 32'h5be00000;
      22845: inst = 32'h244c8000;
      22846: inst = 32'h24428800;
      22847: inst = 32'h8620000;
      22848: inst = 32'h13e00000;
      22849: inst = 32'hfe060f7;
      22850: inst = 32'h5be00000;
      22851: inst = 32'hc6018c3;
      22852: inst = 32'h2a0e0000;
      22853: inst = 32'h294f0000;
      22854: inst = 32'h11200000;
      22855: inst = 32'hd20594b;
      22856: inst = 32'h13e00000;
      22857: inst = 32'hfe0a9ea;
      22858: inst = 32'h5be00000;
      22859: inst = 32'h244c8000;
      22860: inst = 32'h24428800;
      22861: inst = 32'h8620000;
      22862: inst = 32'h2a0e0001;
      22863: inst = 32'h294f0000;
      22864: inst = 32'h11200000;
      22865: inst = 32'hd205955;
      22866: inst = 32'h13e00000;
      22867: inst = 32'hfe0a9ea;
      22868: inst = 32'h5be00000;
      22869: inst = 32'h244c8000;
      22870: inst = 32'h24428800;
      22871: inst = 32'h8620000;
      22872: inst = 32'h2a0e0002;
      22873: inst = 32'h294f0000;
      22874: inst = 32'h11200000;
      22875: inst = 32'hd20595f;
      22876: inst = 32'h13e00000;
      22877: inst = 32'hfe0a9ea;
      22878: inst = 32'h5be00000;
      22879: inst = 32'h244c8000;
      22880: inst = 32'h24428800;
      22881: inst = 32'h8620000;
      22882: inst = 32'h2a0e0003;
      22883: inst = 32'h294f0000;
      22884: inst = 32'h11200000;
      22885: inst = 32'hd205969;
      22886: inst = 32'h13e00000;
      22887: inst = 32'hfe0a9ea;
      22888: inst = 32'h5be00000;
      22889: inst = 32'h244c8000;
      22890: inst = 32'h24428800;
      22891: inst = 32'h8620000;
      22892: inst = 32'h2a0e0004;
      22893: inst = 32'h294f0000;
      22894: inst = 32'h11200000;
      22895: inst = 32'hd205973;
      22896: inst = 32'h13e00000;
      22897: inst = 32'hfe0a9ea;
      22898: inst = 32'h5be00000;
      22899: inst = 32'h244c8000;
      22900: inst = 32'h24428800;
      22901: inst = 32'h8620000;
      22902: inst = 32'h2a0e0005;
      22903: inst = 32'h294f0000;
      22904: inst = 32'h11200000;
      22905: inst = 32'hd20597d;
      22906: inst = 32'h13e00000;
      22907: inst = 32'hfe0a9ea;
      22908: inst = 32'h5be00000;
      22909: inst = 32'h244c8000;
      22910: inst = 32'h24428800;
      22911: inst = 32'h8620000;
      22912: inst = 32'h2a0e0006;
      22913: inst = 32'h294f0000;
      22914: inst = 32'h11200000;
      22915: inst = 32'hd205987;
      22916: inst = 32'h13e00000;
      22917: inst = 32'hfe0a9ea;
      22918: inst = 32'h5be00000;
      22919: inst = 32'h244c8000;
      22920: inst = 32'h24428800;
      22921: inst = 32'h8620000;
      22922: inst = 32'h2a0e0007;
      22923: inst = 32'h294f0000;
      22924: inst = 32'h11200000;
      22925: inst = 32'hd205991;
      22926: inst = 32'h13e00000;
      22927: inst = 32'hfe0a9ea;
      22928: inst = 32'h5be00000;
      22929: inst = 32'h244c8000;
      22930: inst = 32'h24428800;
      22931: inst = 32'h8620000;
      22932: inst = 32'h2a0e0008;
      22933: inst = 32'h294f0000;
      22934: inst = 32'h11200000;
      22935: inst = 32'hd20599b;
      22936: inst = 32'h13e00000;
      22937: inst = 32'hfe0a9ea;
      22938: inst = 32'h5be00000;
      22939: inst = 32'h244c8000;
      22940: inst = 32'h24428800;
      22941: inst = 32'h8620000;
      22942: inst = 32'h2a0e0009;
      22943: inst = 32'h294f0000;
      22944: inst = 32'h11200000;
      22945: inst = 32'hd2059a5;
      22946: inst = 32'h13e00000;
      22947: inst = 32'hfe0a9ea;
      22948: inst = 32'h5be00000;
      22949: inst = 32'h244c8000;
      22950: inst = 32'h24428800;
      22951: inst = 32'h8620000;
      22952: inst = 32'h2a0e0000;
      22953: inst = 32'h294f0001;
      22954: inst = 32'h11200000;
      22955: inst = 32'hd2059af;
      22956: inst = 32'h13e00000;
      22957: inst = 32'hfe0a9ea;
      22958: inst = 32'h5be00000;
      22959: inst = 32'h244c8000;
      22960: inst = 32'h24428800;
      22961: inst = 32'h8620000;
      22962: inst = 32'h2a0e0001;
      22963: inst = 32'h294f0001;
      22964: inst = 32'h11200000;
      22965: inst = 32'hd2059b9;
      22966: inst = 32'h13e00000;
      22967: inst = 32'hfe0a9ea;
      22968: inst = 32'h5be00000;
      22969: inst = 32'h244c8000;
      22970: inst = 32'h24428800;
      22971: inst = 32'h8620000;
      22972: inst = 32'h2a0e0002;
      22973: inst = 32'h294f0001;
      22974: inst = 32'h11200000;
      22975: inst = 32'hd2059c3;
      22976: inst = 32'h13e00000;
      22977: inst = 32'hfe0a9ea;
      22978: inst = 32'h5be00000;
      22979: inst = 32'h244c8000;
      22980: inst = 32'h24428800;
      22981: inst = 32'h8620000;
      22982: inst = 32'h2a0e0003;
      22983: inst = 32'h294f0001;
      22984: inst = 32'h11200000;
      22985: inst = 32'hd2059cd;
      22986: inst = 32'h13e00000;
      22987: inst = 32'hfe0a9ea;
      22988: inst = 32'h5be00000;
      22989: inst = 32'h244c8000;
      22990: inst = 32'h24428800;
      22991: inst = 32'h8620000;
      22992: inst = 32'h2a0e0004;
      22993: inst = 32'h294f0001;
      22994: inst = 32'h11200000;
      22995: inst = 32'hd2059d7;
      22996: inst = 32'h13e00000;
      22997: inst = 32'hfe0a9ea;
      22998: inst = 32'h5be00000;
      22999: inst = 32'h244c8000;
      23000: inst = 32'h24428800;
      23001: inst = 32'h8620000;
      23002: inst = 32'h2a0e0005;
      23003: inst = 32'h294f0001;
      23004: inst = 32'h11200000;
      23005: inst = 32'hd2059e1;
      23006: inst = 32'h13e00000;
      23007: inst = 32'hfe0a9ea;
      23008: inst = 32'h5be00000;
      23009: inst = 32'h244c8000;
      23010: inst = 32'h24428800;
      23011: inst = 32'h8620000;
      23012: inst = 32'h2a0e0006;
      23013: inst = 32'h294f0001;
      23014: inst = 32'h11200000;
      23015: inst = 32'hd2059eb;
      23016: inst = 32'h13e00000;
      23017: inst = 32'hfe0a9ea;
      23018: inst = 32'h5be00000;
      23019: inst = 32'h244c8000;
      23020: inst = 32'h24428800;
      23021: inst = 32'h8620000;
      23022: inst = 32'h2a0e0007;
      23023: inst = 32'h294f0001;
      23024: inst = 32'h11200000;
      23025: inst = 32'hd2059f5;
      23026: inst = 32'h13e00000;
      23027: inst = 32'hfe0a9ea;
      23028: inst = 32'h5be00000;
      23029: inst = 32'h244c8000;
      23030: inst = 32'h24428800;
      23031: inst = 32'h8620000;
      23032: inst = 32'h2a0e0008;
      23033: inst = 32'h294f0001;
      23034: inst = 32'h11200000;
      23035: inst = 32'hd2059ff;
      23036: inst = 32'h13e00000;
      23037: inst = 32'hfe0a9ea;
      23038: inst = 32'h5be00000;
      23039: inst = 32'h244c8000;
      23040: inst = 32'h24428800;
      23041: inst = 32'h8620000;
      23042: inst = 32'h2a0e0009;
      23043: inst = 32'h294f0001;
      23044: inst = 32'h11200000;
      23045: inst = 32'hd205a09;
      23046: inst = 32'h13e00000;
      23047: inst = 32'hfe0a9ea;
      23048: inst = 32'h5be00000;
      23049: inst = 32'h244c8000;
      23050: inst = 32'h24428800;
      23051: inst = 32'h8620000;
      23052: inst = 32'h2a0e0000;
      23053: inst = 32'h294f0002;
      23054: inst = 32'h11200000;
      23055: inst = 32'hd205a13;
      23056: inst = 32'h13e00000;
      23057: inst = 32'hfe0a9ea;
      23058: inst = 32'h5be00000;
      23059: inst = 32'h244c8000;
      23060: inst = 32'h24428800;
      23061: inst = 32'h8620000;
      23062: inst = 32'h2a0e0001;
      23063: inst = 32'h294f0002;
      23064: inst = 32'h11200000;
      23065: inst = 32'hd205a1d;
      23066: inst = 32'h13e00000;
      23067: inst = 32'hfe0a9ea;
      23068: inst = 32'h5be00000;
      23069: inst = 32'h244c8000;
      23070: inst = 32'h24428800;
      23071: inst = 32'h8620000;
      23072: inst = 32'h2a0e0000;
      23073: inst = 32'h294f0003;
      23074: inst = 32'h11200000;
      23075: inst = 32'hd205a27;
      23076: inst = 32'h13e00000;
      23077: inst = 32'hfe0a9ea;
      23078: inst = 32'h5be00000;
      23079: inst = 32'h244c8000;
      23080: inst = 32'h24428800;
      23081: inst = 32'h8620000;
      23082: inst = 32'h2a0e0008;
      23083: inst = 32'h294f0003;
      23084: inst = 32'h11200000;
      23085: inst = 32'hd205a31;
      23086: inst = 32'h13e00000;
      23087: inst = 32'hfe0a9ea;
      23088: inst = 32'h5be00000;
      23089: inst = 32'h244c8000;
      23090: inst = 32'h24428800;
      23091: inst = 32'h8620000;
      23092: inst = 32'h2a0e0000;
      23093: inst = 32'h294f0004;
      23094: inst = 32'h11200000;
      23095: inst = 32'hd205a3b;
      23096: inst = 32'h13e00000;
      23097: inst = 32'hfe0a9ea;
      23098: inst = 32'h5be00000;
      23099: inst = 32'h244c8000;
      23100: inst = 32'h24428800;
      23101: inst = 32'h8620000;
      23102: inst = 32'h2a0e0008;
      23103: inst = 32'h294f0004;
      23104: inst = 32'h11200000;
      23105: inst = 32'hd205a45;
      23106: inst = 32'h13e00000;
      23107: inst = 32'hfe0a9ea;
      23108: inst = 32'h5be00000;
      23109: inst = 32'h244c8000;
      23110: inst = 32'h24428800;
      23111: inst = 32'h8620000;
      23112: inst = 32'h2a0e0000;
      23113: inst = 32'h294f0005;
      23114: inst = 32'h11200000;
      23115: inst = 32'hd205a4f;
      23116: inst = 32'h13e00000;
      23117: inst = 32'hfe0a9ea;
      23118: inst = 32'h5be00000;
      23119: inst = 32'h244c8000;
      23120: inst = 32'h24428800;
      23121: inst = 32'h8620000;
      23122: inst = 32'h2a0e0001;
      23123: inst = 32'h294f0005;
      23124: inst = 32'h11200000;
      23125: inst = 32'hd205a59;
      23126: inst = 32'h13e00000;
      23127: inst = 32'hfe0a9ea;
      23128: inst = 32'h5be00000;
      23129: inst = 32'h244c8000;
      23130: inst = 32'h24428800;
      23131: inst = 32'h8620000;
      23132: inst = 32'h2a0e0000;
      23133: inst = 32'h294f0006;
      23134: inst = 32'h11200000;
      23135: inst = 32'hd205a63;
      23136: inst = 32'h13e00000;
      23137: inst = 32'hfe0a9ea;
      23138: inst = 32'h5be00000;
      23139: inst = 32'h244c8000;
      23140: inst = 32'h24428800;
      23141: inst = 32'h8620000;
      23142: inst = 32'h2a0e0001;
      23143: inst = 32'h294f0006;
      23144: inst = 32'h11200000;
      23145: inst = 32'hd205a6d;
      23146: inst = 32'h13e00000;
      23147: inst = 32'hfe0a9ea;
      23148: inst = 32'h5be00000;
      23149: inst = 32'h244c8000;
      23150: inst = 32'h24428800;
      23151: inst = 32'h8620000;
      23152: inst = 32'hc60d42c;
      23153: inst = 32'h2a0e0002;
      23154: inst = 32'h294f0002;
      23155: inst = 32'h11200000;
      23156: inst = 32'hd205a78;
      23157: inst = 32'h13e00000;
      23158: inst = 32'hfe0a9ea;
      23159: inst = 32'h5be00000;
      23160: inst = 32'h244c8000;
      23161: inst = 32'h24428800;
      23162: inst = 32'h8620000;
      23163: inst = 32'h2a0e0003;
      23164: inst = 32'h294f0002;
      23165: inst = 32'h11200000;
      23166: inst = 32'hd205a82;
      23167: inst = 32'h13e00000;
      23168: inst = 32'hfe0a9ea;
      23169: inst = 32'h5be00000;
      23170: inst = 32'h244c8000;
      23171: inst = 32'h24428800;
      23172: inst = 32'h8620000;
      23173: inst = 32'h2a0e0004;
      23174: inst = 32'h294f0002;
      23175: inst = 32'h11200000;
      23176: inst = 32'hd205a8c;
      23177: inst = 32'h13e00000;
      23178: inst = 32'hfe0a9ea;
      23179: inst = 32'h5be00000;
      23180: inst = 32'h244c8000;
      23181: inst = 32'h24428800;
      23182: inst = 32'h8620000;
      23183: inst = 32'h2a0e0005;
      23184: inst = 32'h294f0002;
      23185: inst = 32'h11200000;
      23186: inst = 32'hd205a96;
      23187: inst = 32'h13e00000;
      23188: inst = 32'hfe0a9ea;
      23189: inst = 32'h5be00000;
      23190: inst = 32'h244c8000;
      23191: inst = 32'h24428800;
      23192: inst = 32'h8620000;
      23193: inst = 32'h2a0e0006;
      23194: inst = 32'h294f0002;
      23195: inst = 32'h11200000;
      23196: inst = 32'hd205aa0;
      23197: inst = 32'h13e00000;
      23198: inst = 32'hfe0a9ea;
      23199: inst = 32'h5be00000;
      23200: inst = 32'h244c8000;
      23201: inst = 32'h24428800;
      23202: inst = 32'h8620000;
      23203: inst = 32'h2a0e0007;
      23204: inst = 32'h294f0002;
      23205: inst = 32'h11200000;
      23206: inst = 32'hd205aaa;
      23207: inst = 32'h13e00000;
      23208: inst = 32'hfe0a9ea;
      23209: inst = 32'h5be00000;
      23210: inst = 32'h244c8000;
      23211: inst = 32'h24428800;
      23212: inst = 32'h8620000;
      23213: inst = 32'h2a0e0008;
      23214: inst = 32'h294f0002;
      23215: inst = 32'h11200000;
      23216: inst = 32'hd205ab4;
      23217: inst = 32'h13e00000;
      23218: inst = 32'hfe0a9ea;
      23219: inst = 32'h5be00000;
      23220: inst = 32'h244c8000;
      23221: inst = 32'h24428800;
      23222: inst = 32'h8620000;
      23223: inst = 32'h2a0e0009;
      23224: inst = 32'h294f0002;
      23225: inst = 32'h11200000;
      23226: inst = 32'hd205abe;
      23227: inst = 32'h13e00000;
      23228: inst = 32'hfe0a9ea;
      23229: inst = 32'h5be00000;
      23230: inst = 32'h244c8000;
      23231: inst = 32'h24428800;
      23232: inst = 32'h8620000;
      23233: inst = 32'h2a0e0002;
      23234: inst = 32'h294f0005;
      23235: inst = 32'h11200000;
      23236: inst = 32'hd205ac8;
      23237: inst = 32'h13e00000;
      23238: inst = 32'hfe0a9ea;
      23239: inst = 32'h5be00000;
      23240: inst = 32'h244c8000;
      23241: inst = 32'h24428800;
      23242: inst = 32'h8620000;
      23243: inst = 32'h2a0e0002;
      23244: inst = 32'h294f0006;
      23245: inst = 32'h11200000;
      23246: inst = 32'hd205ad2;
      23247: inst = 32'h13e00000;
      23248: inst = 32'hfe0a9ea;
      23249: inst = 32'h5be00000;
      23250: inst = 32'h244c8000;
      23251: inst = 32'h24428800;
      23252: inst = 32'h8620000;
      23253: inst = 32'h2a0e0003;
      23254: inst = 32'h294f000b;
      23255: inst = 32'h11200000;
      23256: inst = 32'hd205adc;
      23257: inst = 32'h13e00000;
      23258: inst = 32'hfe0a9ea;
      23259: inst = 32'h5be00000;
      23260: inst = 32'h244c8000;
      23261: inst = 32'h24428800;
      23262: inst = 32'h8620000;
      23263: inst = 32'h2a0e0006;
      23264: inst = 32'h294f000b;
      23265: inst = 32'h11200000;
      23266: inst = 32'hd205ae6;
      23267: inst = 32'h13e00000;
      23268: inst = 32'hfe0a9ea;
      23269: inst = 32'h5be00000;
      23270: inst = 32'h244c8000;
      23271: inst = 32'h24428800;
      23272: inst = 32'h8620000;
      23273: inst = 32'hc60f4ce;
      23274: inst = 32'h2a0e0001;
      23275: inst = 32'h294f0003;
      23276: inst = 32'h11200000;
      23277: inst = 32'hd205af1;
      23278: inst = 32'h13e00000;
      23279: inst = 32'hfe0a9ea;
      23280: inst = 32'h5be00000;
      23281: inst = 32'h244c8000;
      23282: inst = 32'h24428800;
      23283: inst = 32'h8620000;
      23284: inst = 32'h2a0e0002;
      23285: inst = 32'h294f0003;
      23286: inst = 32'h11200000;
      23287: inst = 32'hd205afb;
      23288: inst = 32'h13e00000;
      23289: inst = 32'hfe0a9ea;
      23290: inst = 32'h5be00000;
      23291: inst = 32'h244c8000;
      23292: inst = 32'h24428800;
      23293: inst = 32'h8620000;
      23294: inst = 32'h2a0e0003;
      23295: inst = 32'h294f0003;
      23296: inst = 32'h11200000;
      23297: inst = 32'hd205b05;
      23298: inst = 32'h13e00000;
      23299: inst = 32'hfe0a9ea;
      23300: inst = 32'h5be00000;
      23301: inst = 32'h244c8000;
      23302: inst = 32'h24428800;
      23303: inst = 32'h8620000;
      23304: inst = 32'h2a0e0004;
      23305: inst = 32'h294f0003;
      23306: inst = 32'h11200000;
      23307: inst = 32'hd205b0f;
      23308: inst = 32'h13e00000;
      23309: inst = 32'hfe0a9ea;
      23310: inst = 32'h5be00000;
      23311: inst = 32'h244c8000;
      23312: inst = 32'h24428800;
      23313: inst = 32'h8620000;
      23314: inst = 32'h2a0e0005;
      23315: inst = 32'h294f0003;
      23316: inst = 32'h11200000;
      23317: inst = 32'hd205b19;
      23318: inst = 32'h13e00000;
      23319: inst = 32'hfe0a9ea;
      23320: inst = 32'h5be00000;
      23321: inst = 32'h244c8000;
      23322: inst = 32'h24428800;
      23323: inst = 32'h8620000;
      23324: inst = 32'h2a0e0006;
      23325: inst = 32'h294f0003;
      23326: inst = 32'h11200000;
      23327: inst = 32'hd205b23;
      23328: inst = 32'h13e00000;
      23329: inst = 32'hfe0a9ea;
      23330: inst = 32'h5be00000;
      23331: inst = 32'h244c8000;
      23332: inst = 32'h24428800;
      23333: inst = 32'h8620000;
      23334: inst = 32'h2a0e0007;
      23335: inst = 32'h294f0003;
      23336: inst = 32'h11200000;
      23337: inst = 32'hd205b2d;
      23338: inst = 32'h13e00000;
      23339: inst = 32'hfe0a9ea;
      23340: inst = 32'h5be00000;
      23341: inst = 32'h244c8000;
      23342: inst = 32'h24428800;
      23343: inst = 32'h8620000;
      23344: inst = 32'h2a0e0009;
      23345: inst = 32'h294f0003;
      23346: inst = 32'h11200000;
      23347: inst = 32'hd205b37;
      23348: inst = 32'h13e00000;
      23349: inst = 32'hfe0a9ea;
      23350: inst = 32'h5be00000;
      23351: inst = 32'h244c8000;
      23352: inst = 32'h24428800;
      23353: inst = 32'h8620000;
      23354: inst = 32'h2a0e0001;
      23355: inst = 32'h294f0004;
      23356: inst = 32'h11200000;
      23357: inst = 32'hd205b41;
      23358: inst = 32'h13e00000;
      23359: inst = 32'hfe0a9ea;
      23360: inst = 32'h5be00000;
      23361: inst = 32'h244c8000;
      23362: inst = 32'h24428800;
      23363: inst = 32'h8620000;
      23364: inst = 32'h2a0e0002;
      23365: inst = 32'h294f0004;
      23366: inst = 32'h11200000;
      23367: inst = 32'hd205b4b;
      23368: inst = 32'h13e00000;
      23369: inst = 32'hfe0a9ea;
      23370: inst = 32'h5be00000;
      23371: inst = 32'h244c8000;
      23372: inst = 32'h24428800;
      23373: inst = 32'h8620000;
      23374: inst = 32'h2a0e0003;
      23375: inst = 32'h294f0004;
      23376: inst = 32'h11200000;
      23377: inst = 32'hd205b55;
      23378: inst = 32'h13e00000;
      23379: inst = 32'hfe0a9ea;
      23380: inst = 32'h5be00000;
      23381: inst = 32'h244c8000;
      23382: inst = 32'h24428800;
      23383: inst = 32'h8620000;
      23384: inst = 32'h2a0e0004;
      23385: inst = 32'h294f0004;
      23386: inst = 32'h11200000;
      23387: inst = 32'hd205b5f;
      23388: inst = 32'h13e00000;
      23389: inst = 32'hfe0a9ea;
      23390: inst = 32'h5be00000;
      23391: inst = 32'h244c8000;
      23392: inst = 32'h24428800;
      23393: inst = 32'h8620000;
      23394: inst = 32'h2a0e0005;
      23395: inst = 32'h294f0004;
      23396: inst = 32'h11200000;
      23397: inst = 32'hd205b69;
      23398: inst = 32'h13e00000;
      23399: inst = 32'hfe0a9ea;
      23400: inst = 32'h5be00000;
      23401: inst = 32'h244c8000;
      23402: inst = 32'h24428800;
      23403: inst = 32'h8620000;
      23404: inst = 32'h2a0e0006;
      23405: inst = 32'h294f0004;
      23406: inst = 32'h11200000;
      23407: inst = 32'hd205b73;
      23408: inst = 32'h13e00000;
      23409: inst = 32'hfe0a9ea;
      23410: inst = 32'h5be00000;
      23411: inst = 32'h244c8000;
      23412: inst = 32'h24428800;
      23413: inst = 32'h8620000;
      23414: inst = 32'h2a0e0007;
      23415: inst = 32'h294f0004;
      23416: inst = 32'h11200000;
      23417: inst = 32'hd205b7d;
      23418: inst = 32'h13e00000;
      23419: inst = 32'hfe0a9ea;
      23420: inst = 32'h5be00000;
      23421: inst = 32'h244c8000;
      23422: inst = 32'h24428800;
      23423: inst = 32'h8620000;
      23424: inst = 32'h2a0e0009;
      23425: inst = 32'h294f0004;
      23426: inst = 32'h11200000;
      23427: inst = 32'hd205b87;
      23428: inst = 32'h13e00000;
      23429: inst = 32'hfe0a9ea;
      23430: inst = 32'h5be00000;
      23431: inst = 32'h244c8000;
      23432: inst = 32'h24428800;
      23433: inst = 32'h8620000;
      23434: inst = 32'h2a0e0003;
      23435: inst = 32'h294f0005;
      23436: inst = 32'h11200000;
      23437: inst = 32'hd205b91;
      23438: inst = 32'h13e00000;
      23439: inst = 32'hfe0a9ea;
      23440: inst = 32'h5be00000;
      23441: inst = 32'h244c8000;
      23442: inst = 32'h24428800;
      23443: inst = 32'h8620000;
      23444: inst = 32'h2a0e0004;
      23445: inst = 32'h294f0005;
      23446: inst = 32'h11200000;
      23447: inst = 32'hd205b9b;
      23448: inst = 32'h13e00000;
      23449: inst = 32'hfe0a9ea;
      23450: inst = 32'h5be00000;
      23451: inst = 32'h244c8000;
      23452: inst = 32'h24428800;
      23453: inst = 32'h8620000;
      23454: inst = 32'h2a0e0005;
      23455: inst = 32'h294f0005;
      23456: inst = 32'h11200000;
      23457: inst = 32'hd205ba5;
      23458: inst = 32'h13e00000;
      23459: inst = 32'hfe0a9ea;
      23460: inst = 32'h5be00000;
      23461: inst = 32'h244c8000;
      23462: inst = 32'h24428800;
      23463: inst = 32'h8620000;
      23464: inst = 32'h2a0e0006;
      23465: inst = 32'h294f0005;
      23466: inst = 32'h11200000;
      23467: inst = 32'hd205baf;
      23468: inst = 32'h13e00000;
      23469: inst = 32'hfe0a9ea;
      23470: inst = 32'h5be00000;
      23471: inst = 32'h244c8000;
      23472: inst = 32'h24428800;
      23473: inst = 32'h8620000;
      23474: inst = 32'h2a0e0007;
      23475: inst = 32'h294f0005;
      23476: inst = 32'h11200000;
      23477: inst = 32'hd205bb9;
      23478: inst = 32'h13e00000;
      23479: inst = 32'hfe0a9ea;
      23480: inst = 32'h5be00000;
      23481: inst = 32'h244c8000;
      23482: inst = 32'h24428800;
      23483: inst = 32'h8620000;
      23484: inst = 32'h2a0e0008;
      23485: inst = 32'h294f0005;
      23486: inst = 32'h11200000;
      23487: inst = 32'hd205bc3;
      23488: inst = 32'h13e00000;
      23489: inst = 32'hfe0a9ea;
      23490: inst = 32'h5be00000;
      23491: inst = 32'h244c8000;
      23492: inst = 32'h24428800;
      23493: inst = 32'h8620000;
      23494: inst = 32'h2a0e0009;
      23495: inst = 32'h294f0005;
      23496: inst = 32'h11200000;
      23497: inst = 32'hd205bcd;
      23498: inst = 32'h13e00000;
      23499: inst = 32'hfe0a9ea;
      23500: inst = 32'h5be00000;
      23501: inst = 32'h244c8000;
      23502: inst = 32'h24428800;
      23503: inst = 32'h8620000;
      23504: inst = 32'h2a0e0003;
      23505: inst = 32'h294f0006;
      23506: inst = 32'h11200000;
      23507: inst = 32'hd205bd7;
      23508: inst = 32'h13e00000;
      23509: inst = 32'hfe0a9ea;
      23510: inst = 32'h5be00000;
      23511: inst = 32'h244c8000;
      23512: inst = 32'h24428800;
      23513: inst = 32'h8620000;
      23514: inst = 32'h2a0e0004;
      23515: inst = 32'h294f0006;
      23516: inst = 32'h11200000;
      23517: inst = 32'hd205be1;
      23518: inst = 32'h13e00000;
      23519: inst = 32'hfe0a9ea;
      23520: inst = 32'h5be00000;
      23521: inst = 32'h244c8000;
      23522: inst = 32'h24428800;
      23523: inst = 32'h8620000;
      23524: inst = 32'h2a0e0005;
      23525: inst = 32'h294f0006;
      23526: inst = 32'h11200000;
      23527: inst = 32'hd205beb;
      23528: inst = 32'h13e00000;
      23529: inst = 32'hfe0a9ea;
      23530: inst = 32'h5be00000;
      23531: inst = 32'h244c8000;
      23532: inst = 32'h24428800;
      23533: inst = 32'h8620000;
      23534: inst = 32'h2a0e0006;
      23535: inst = 32'h294f0006;
      23536: inst = 32'h11200000;
      23537: inst = 32'hd205bf5;
      23538: inst = 32'h13e00000;
      23539: inst = 32'hfe0a9ea;
      23540: inst = 32'h5be00000;
      23541: inst = 32'h244c8000;
      23542: inst = 32'h24428800;
      23543: inst = 32'h8620000;
      23544: inst = 32'h2a0e0007;
      23545: inst = 32'h294f0006;
      23546: inst = 32'h11200000;
      23547: inst = 32'hd205bff;
      23548: inst = 32'h13e00000;
      23549: inst = 32'hfe0a9ea;
      23550: inst = 32'h5be00000;
      23551: inst = 32'h244c8000;
      23552: inst = 32'h24428800;
      23553: inst = 32'h8620000;
      23554: inst = 32'h2a0e0008;
      23555: inst = 32'h294f0006;
      23556: inst = 32'h11200000;
      23557: inst = 32'hd205c09;
      23558: inst = 32'h13e00000;
      23559: inst = 32'hfe0a9ea;
      23560: inst = 32'h5be00000;
      23561: inst = 32'h244c8000;
      23562: inst = 32'h24428800;
      23563: inst = 32'h8620000;
      23564: inst = 32'h2a0e0009;
      23565: inst = 32'h294f0006;
      23566: inst = 32'h11200000;
      23567: inst = 32'hd205c13;
      23568: inst = 32'h13e00000;
      23569: inst = 32'hfe0a9ea;
      23570: inst = 32'h5be00000;
      23571: inst = 32'h244c8000;
      23572: inst = 32'h24428800;
      23573: inst = 32'h8620000;
      23574: inst = 32'h2a0e0004;
      23575: inst = 32'h294f0008;
      23576: inst = 32'h11200000;
      23577: inst = 32'hd205c1d;
      23578: inst = 32'h13e00000;
      23579: inst = 32'hfe0a9ea;
      23580: inst = 32'h5be00000;
      23581: inst = 32'h244c8000;
      23582: inst = 32'h24428800;
      23583: inst = 32'h8620000;
      23584: inst = 32'h2a0e0008;
      23585: inst = 32'h294f0008;
      23586: inst = 32'h11200000;
      23587: inst = 32'hd205c27;
      23588: inst = 32'h13e00000;
      23589: inst = 32'hfe0a9ea;
      23590: inst = 32'h5be00000;
      23591: inst = 32'h244c8000;
      23592: inst = 32'h24428800;
      23593: inst = 32'h8620000;
      23594: inst = 32'h2a0e0004;
      23595: inst = 32'h294f0009;
      23596: inst = 32'h11200000;
      23597: inst = 32'hd205c31;
      23598: inst = 32'h13e00000;
      23599: inst = 32'hfe0a9ea;
      23600: inst = 32'h5be00000;
      23601: inst = 32'h244c8000;
      23602: inst = 32'h24428800;
      23603: inst = 32'h8620000;
      23604: inst = 32'hc607841;
      23605: inst = 32'h2a0e0002;
      23606: inst = 32'h294f0007;
      23607: inst = 32'h11200000;
      23608: inst = 32'hd205c3c;
      23609: inst = 32'h13e00000;
      23610: inst = 32'hfe0a9ea;
      23611: inst = 32'h5be00000;
      23612: inst = 32'h244c8000;
      23613: inst = 32'h24428800;
      23614: inst = 32'h8620000;
      23615: inst = 32'h2a0e0002;
      23616: inst = 32'h294f0008;
      23617: inst = 32'h11200000;
      23618: inst = 32'hd205c46;
      23619: inst = 32'h13e00000;
      23620: inst = 32'hfe0a9ea;
      23621: inst = 32'h5be00000;
      23622: inst = 32'h244c8000;
      23623: inst = 32'h24428800;
      23624: inst = 32'h8620000;
      23625: inst = 32'hc60a000;
      23626: inst = 32'h2a0e0003;
      23627: inst = 32'h294f0007;
      23628: inst = 32'h11200000;
      23629: inst = 32'hd205c51;
      23630: inst = 32'h13e00000;
      23631: inst = 32'hfe0a9ea;
      23632: inst = 32'h5be00000;
      23633: inst = 32'h244c8000;
      23634: inst = 32'h24428800;
      23635: inst = 32'h8620000;
      23636: inst = 32'h2a0e0004;
      23637: inst = 32'h294f0007;
      23638: inst = 32'h11200000;
      23639: inst = 32'hd205c5b;
      23640: inst = 32'h13e00000;
      23641: inst = 32'hfe0a9ea;
      23642: inst = 32'h5be00000;
      23643: inst = 32'h244c8000;
      23644: inst = 32'h24428800;
      23645: inst = 32'h8620000;
      23646: inst = 32'h2a0e0005;
      23647: inst = 32'h294f0007;
      23648: inst = 32'h11200000;
      23649: inst = 32'hd205c65;
      23650: inst = 32'h13e00000;
      23651: inst = 32'hfe0a9ea;
      23652: inst = 32'h5be00000;
      23653: inst = 32'h244c8000;
      23654: inst = 32'h24428800;
      23655: inst = 32'h8620000;
      23656: inst = 32'h2a0e0006;
      23657: inst = 32'h294f0007;
      23658: inst = 32'h11200000;
      23659: inst = 32'hd205c6f;
      23660: inst = 32'h13e00000;
      23661: inst = 32'hfe0a9ea;
      23662: inst = 32'h5be00000;
      23663: inst = 32'h244c8000;
      23664: inst = 32'h24428800;
      23665: inst = 32'h8620000;
      23666: inst = 32'h2a0e0007;
      23667: inst = 32'h294f0007;
      23668: inst = 32'h11200000;
      23669: inst = 32'hd205c79;
      23670: inst = 32'h13e00000;
      23671: inst = 32'hfe0a9ea;
      23672: inst = 32'h5be00000;
      23673: inst = 32'h244c8000;
      23674: inst = 32'h24428800;
      23675: inst = 32'h8620000;
      23676: inst = 32'h2a0e0003;
      23677: inst = 32'h294f0008;
      23678: inst = 32'h11200000;
      23679: inst = 32'hd205c83;
      23680: inst = 32'h13e00000;
      23681: inst = 32'hfe0a9ea;
      23682: inst = 32'h5be00000;
      23683: inst = 32'h244c8000;
      23684: inst = 32'h24428800;
      23685: inst = 32'h8620000;
      23686: inst = 32'h2a0e0005;
      23687: inst = 32'h294f0008;
      23688: inst = 32'h11200000;
      23689: inst = 32'hd205c8d;
      23690: inst = 32'h13e00000;
      23691: inst = 32'hfe0a9ea;
      23692: inst = 32'h5be00000;
      23693: inst = 32'h244c8000;
      23694: inst = 32'h24428800;
      23695: inst = 32'h8620000;
      23696: inst = 32'h2a0e0006;
      23697: inst = 32'h294f0008;
      23698: inst = 32'h11200000;
      23699: inst = 32'hd205c97;
      23700: inst = 32'h13e00000;
      23701: inst = 32'hfe0a9ea;
      23702: inst = 32'h5be00000;
      23703: inst = 32'h244c8000;
      23704: inst = 32'h24428800;
      23705: inst = 32'h8620000;
      23706: inst = 32'h2a0e0007;
      23707: inst = 32'h294f0008;
      23708: inst = 32'h11200000;
      23709: inst = 32'hd205ca1;
      23710: inst = 32'h13e00000;
      23711: inst = 32'hfe0a9ea;
      23712: inst = 32'h5be00000;
      23713: inst = 32'h244c8000;
      23714: inst = 32'h24428800;
      23715: inst = 32'h8620000;
      23716: inst = 32'h2a0e0002;
      23717: inst = 32'h294f0009;
      23718: inst = 32'h11200000;
      23719: inst = 32'hd205cab;
      23720: inst = 32'h13e00000;
      23721: inst = 32'hfe0a9ea;
      23722: inst = 32'h5be00000;
      23723: inst = 32'h244c8000;
      23724: inst = 32'h24428800;
      23725: inst = 32'h8620000;
      23726: inst = 32'h2a0e0003;
      23727: inst = 32'h294f0009;
      23728: inst = 32'h11200000;
      23729: inst = 32'hd205cb5;
      23730: inst = 32'h13e00000;
      23731: inst = 32'hfe0a9ea;
      23732: inst = 32'h5be00000;
      23733: inst = 32'h244c8000;
      23734: inst = 32'h24428800;
      23735: inst = 32'h8620000;
      23736: inst = 32'h2a0e0005;
      23737: inst = 32'h294f0009;
      23738: inst = 32'h11200000;
      23739: inst = 32'hd205cbf;
      23740: inst = 32'h13e00000;
      23741: inst = 32'hfe0a9ea;
      23742: inst = 32'h5be00000;
      23743: inst = 32'h244c8000;
      23744: inst = 32'h24428800;
      23745: inst = 32'h8620000;
      23746: inst = 32'h2a0e0006;
      23747: inst = 32'h294f0009;
      23748: inst = 32'h11200000;
      23749: inst = 32'hd205cc9;
      23750: inst = 32'h13e00000;
      23751: inst = 32'hfe0a9ea;
      23752: inst = 32'h5be00000;
      23753: inst = 32'h244c8000;
      23754: inst = 32'h24428800;
      23755: inst = 32'h8620000;
      23756: inst = 32'h2a0e0007;
      23757: inst = 32'h294f0009;
      23758: inst = 32'h11200000;
      23759: inst = 32'hd205cd3;
      23760: inst = 32'h13e00000;
      23761: inst = 32'hfe0a9ea;
      23762: inst = 32'h5be00000;
      23763: inst = 32'h244c8000;
      23764: inst = 32'h24428800;
      23765: inst = 32'h8620000;
      23766: inst = 32'hc6010ac;
      23767: inst = 32'h2a0e0002;
      23768: inst = 32'h294f000a;
      23769: inst = 32'h11200000;
      23770: inst = 32'hd205cde;
      23771: inst = 32'h13e00000;
      23772: inst = 32'hfe0a9ea;
      23773: inst = 32'h5be00000;
      23774: inst = 32'h244c8000;
      23775: inst = 32'h24428800;
      23776: inst = 32'h8620000;
      23777: inst = 32'h2a0e0003;
      23778: inst = 32'h294f000a;
      23779: inst = 32'h11200000;
      23780: inst = 32'hd205ce8;
      23781: inst = 32'h13e00000;
      23782: inst = 32'hfe0a9ea;
      23783: inst = 32'h5be00000;
      23784: inst = 32'h244c8000;
      23785: inst = 32'h24428800;
      23786: inst = 32'h8620000;
      23787: inst = 32'h2a0e0004;
      23788: inst = 32'h294f000a;
      23789: inst = 32'h11200000;
      23790: inst = 32'hd205cf2;
      23791: inst = 32'h13e00000;
      23792: inst = 32'hfe0a9ea;
      23793: inst = 32'h5be00000;
      23794: inst = 32'h244c8000;
      23795: inst = 32'h24428800;
      23796: inst = 32'h8620000;
      23797: inst = 32'h2a0e0005;
      23798: inst = 32'h294f000a;
      23799: inst = 32'h11200000;
      23800: inst = 32'hd205cfc;
      23801: inst = 32'h13e00000;
      23802: inst = 32'hfe0a9ea;
      23803: inst = 32'h5be00000;
      23804: inst = 32'h244c8000;
      23805: inst = 32'h24428800;
      23806: inst = 32'h8620000;
      23807: inst = 32'h2a0e0006;
      23808: inst = 32'h294f000a;
      23809: inst = 32'h11200000;
      23810: inst = 32'hd205d06;
      23811: inst = 32'h13e00000;
      23812: inst = 32'hfe0a9ea;
      23813: inst = 32'h5be00000;
      23814: inst = 32'h244c8000;
      23815: inst = 32'h24428800;
      23816: inst = 32'h8620000;
      23817: inst = 32'h2a0e0007;
      23818: inst = 32'h294f000a;
      23819: inst = 32'h11200000;
      23820: inst = 32'hd205d10;
      23821: inst = 32'h13e00000;
      23822: inst = 32'hfe0a9ea;
      23823: inst = 32'h5be00000;
      23824: inst = 32'h244c8000;
      23825: inst = 32'h24428800;
      23826: inst = 32'h8620000;
      23827: inst = 32'h13e00000;
      23828: inst = 32'hfe05d1a;
      23829: inst = 32'h20200003;
      23830: inst = 32'h5be00000;
      23831: inst = 32'h13e00000;
      23832: inst = 32'hfe060f7;
      23833: inst = 32'h5be00000;
      23834: inst = 32'h13e00000;
      23835: inst = 32'hfe060f7;
      23836: inst = 32'h5be00000;
      23837: inst = 32'hc6018c3;
      23838: inst = 32'h2a0e000a;
      23839: inst = 32'h294f0000;
      23840: inst = 32'h11200000;
      23841: inst = 32'hd205d25;
      23842: inst = 32'h13e00000;
      23843: inst = 32'hfe0a9ea;
      23844: inst = 32'h5be00000;
      23845: inst = 32'h244c8000;
      23846: inst = 32'h24428800;
      23847: inst = 32'h8620000;
      23848: inst = 32'h2a0e0009;
      23849: inst = 32'h294f0000;
      23850: inst = 32'h11200000;
      23851: inst = 32'hd205d2f;
      23852: inst = 32'h13e00000;
      23853: inst = 32'hfe0a9ea;
      23854: inst = 32'h5be00000;
      23855: inst = 32'h244c8000;
      23856: inst = 32'h24428800;
      23857: inst = 32'h8620000;
      23858: inst = 32'h2a0e0008;
      23859: inst = 32'h294f0000;
      23860: inst = 32'h11200000;
      23861: inst = 32'hd205d39;
      23862: inst = 32'h13e00000;
      23863: inst = 32'hfe0a9ea;
      23864: inst = 32'h5be00000;
      23865: inst = 32'h244c8000;
      23866: inst = 32'h24428800;
      23867: inst = 32'h8620000;
      23868: inst = 32'h2a0e0007;
      23869: inst = 32'h294f0000;
      23870: inst = 32'h11200000;
      23871: inst = 32'hd205d43;
      23872: inst = 32'h13e00000;
      23873: inst = 32'hfe0a9ea;
      23874: inst = 32'h5be00000;
      23875: inst = 32'h244c8000;
      23876: inst = 32'h24428800;
      23877: inst = 32'h8620000;
      23878: inst = 32'h2a0e0006;
      23879: inst = 32'h294f0000;
      23880: inst = 32'h11200000;
      23881: inst = 32'hd205d4d;
      23882: inst = 32'h13e00000;
      23883: inst = 32'hfe0a9ea;
      23884: inst = 32'h5be00000;
      23885: inst = 32'h244c8000;
      23886: inst = 32'h24428800;
      23887: inst = 32'h8620000;
      23888: inst = 32'h2a0e0005;
      23889: inst = 32'h294f0000;
      23890: inst = 32'h11200000;
      23891: inst = 32'hd205d57;
      23892: inst = 32'h13e00000;
      23893: inst = 32'hfe0a9ea;
      23894: inst = 32'h5be00000;
      23895: inst = 32'h244c8000;
      23896: inst = 32'h24428800;
      23897: inst = 32'h8620000;
      23898: inst = 32'h2a0e0004;
      23899: inst = 32'h294f0000;
      23900: inst = 32'h11200000;
      23901: inst = 32'hd205d61;
      23902: inst = 32'h13e00000;
      23903: inst = 32'hfe0a9ea;
      23904: inst = 32'h5be00000;
      23905: inst = 32'h244c8000;
      23906: inst = 32'h24428800;
      23907: inst = 32'h8620000;
      23908: inst = 32'h2a0e0003;
      23909: inst = 32'h294f0000;
      23910: inst = 32'h11200000;
      23911: inst = 32'hd205d6b;
      23912: inst = 32'h13e00000;
      23913: inst = 32'hfe0a9ea;
      23914: inst = 32'h5be00000;
      23915: inst = 32'h244c8000;
      23916: inst = 32'h24428800;
      23917: inst = 32'h8620000;
      23918: inst = 32'h2a0e0002;
      23919: inst = 32'h294f0000;
      23920: inst = 32'h11200000;
      23921: inst = 32'hd205d75;
      23922: inst = 32'h13e00000;
      23923: inst = 32'hfe0a9ea;
      23924: inst = 32'h5be00000;
      23925: inst = 32'h244c8000;
      23926: inst = 32'h24428800;
      23927: inst = 32'h8620000;
      23928: inst = 32'h2a0e0001;
      23929: inst = 32'h294f0000;
      23930: inst = 32'h11200000;
      23931: inst = 32'hd205d7f;
      23932: inst = 32'h13e00000;
      23933: inst = 32'hfe0a9ea;
      23934: inst = 32'h5be00000;
      23935: inst = 32'h244c8000;
      23936: inst = 32'h24428800;
      23937: inst = 32'h8620000;
      23938: inst = 32'h2a0e000a;
      23939: inst = 32'h294f0001;
      23940: inst = 32'h11200000;
      23941: inst = 32'hd205d89;
      23942: inst = 32'h13e00000;
      23943: inst = 32'hfe0a9ea;
      23944: inst = 32'h5be00000;
      23945: inst = 32'h244c8000;
      23946: inst = 32'h24428800;
      23947: inst = 32'h8620000;
      23948: inst = 32'h2a0e0009;
      23949: inst = 32'h294f0001;
      23950: inst = 32'h11200000;
      23951: inst = 32'hd205d93;
      23952: inst = 32'h13e00000;
      23953: inst = 32'hfe0a9ea;
      23954: inst = 32'h5be00000;
      23955: inst = 32'h244c8000;
      23956: inst = 32'h24428800;
      23957: inst = 32'h8620000;
      23958: inst = 32'h2a0e0008;
      23959: inst = 32'h294f0001;
      23960: inst = 32'h11200000;
      23961: inst = 32'hd205d9d;
      23962: inst = 32'h13e00000;
      23963: inst = 32'hfe0a9ea;
      23964: inst = 32'h5be00000;
      23965: inst = 32'h244c8000;
      23966: inst = 32'h24428800;
      23967: inst = 32'h8620000;
      23968: inst = 32'h2a0e0007;
      23969: inst = 32'h294f0001;
      23970: inst = 32'h11200000;
      23971: inst = 32'hd205da7;
      23972: inst = 32'h13e00000;
      23973: inst = 32'hfe0a9ea;
      23974: inst = 32'h5be00000;
      23975: inst = 32'h244c8000;
      23976: inst = 32'h24428800;
      23977: inst = 32'h8620000;
      23978: inst = 32'h2a0e0006;
      23979: inst = 32'h294f0001;
      23980: inst = 32'h11200000;
      23981: inst = 32'hd205db1;
      23982: inst = 32'h13e00000;
      23983: inst = 32'hfe0a9ea;
      23984: inst = 32'h5be00000;
      23985: inst = 32'h244c8000;
      23986: inst = 32'h24428800;
      23987: inst = 32'h8620000;
      23988: inst = 32'h2a0e0005;
      23989: inst = 32'h294f0001;
      23990: inst = 32'h11200000;
      23991: inst = 32'hd205dbb;
      23992: inst = 32'h13e00000;
      23993: inst = 32'hfe0a9ea;
      23994: inst = 32'h5be00000;
      23995: inst = 32'h244c8000;
      23996: inst = 32'h24428800;
      23997: inst = 32'h8620000;
      23998: inst = 32'h2a0e0004;
      23999: inst = 32'h294f0001;
      24000: inst = 32'h11200000;
      24001: inst = 32'hd205dc5;
      24002: inst = 32'h13e00000;
      24003: inst = 32'hfe0a9ea;
      24004: inst = 32'h5be00000;
      24005: inst = 32'h244c8000;
      24006: inst = 32'h24428800;
      24007: inst = 32'h8620000;
      24008: inst = 32'h2a0e0003;
      24009: inst = 32'h294f0001;
      24010: inst = 32'h11200000;
      24011: inst = 32'hd205dcf;
      24012: inst = 32'h13e00000;
      24013: inst = 32'hfe0a9ea;
      24014: inst = 32'h5be00000;
      24015: inst = 32'h244c8000;
      24016: inst = 32'h24428800;
      24017: inst = 32'h8620000;
      24018: inst = 32'h2a0e0002;
      24019: inst = 32'h294f0001;
      24020: inst = 32'h11200000;
      24021: inst = 32'hd205dd9;
      24022: inst = 32'h13e00000;
      24023: inst = 32'hfe0a9ea;
      24024: inst = 32'h5be00000;
      24025: inst = 32'h244c8000;
      24026: inst = 32'h24428800;
      24027: inst = 32'h8620000;
      24028: inst = 32'h2a0e0001;
      24029: inst = 32'h294f0001;
      24030: inst = 32'h11200000;
      24031: inst = 32'hd205de3;
      24032: inst = 32'h13e00000;
      24033: inst = 32'hfe0a9ea;
      24034: inst = 32'h5be00000;
      24035: inst = 32'h244c8000;
      24036: inst = 32'h24428800;
      24037: inst = 32'h8620000;
      24038: inst = 32'h2a0e000a;
      24039: inst = 32'h294f0002;
      24040: inst = 32'h11200000;
      24041: inst = 32'hd205ded;
      24042: inst = 32'h13e00000;
      24043: inst = 32'hfe0a9ea;
      24044: inst = 32'h5be00000;
      24045: inst = 32'h244c8000;
      24046: inst = 32'h24428800;
      24047: inst = 32'h8620000;
      24048: inst = 32'h2a0e0009;
      24049: inst = 32'h294f0002;
      24050: inst = 32'h11200000;
      24051: inst = 32'hd205df7;
      24052: inst = 32'h13e00000;
      24053: inst = 32'hfe0a9ea;
      24054: inst = 32'h5be00000;
      24055: inst = 32'h244c8000;
      24056: inst = 32'h24428800;
      24057: inst = 32'h8620000;
      24058: inst = 32'h2a0e000a;
      24059: inst = 32'h294f0003;
      24060: inst = 32'h11200000;
      24061: inst = 32'hd205e01;
      24062: inst = 32'h13e00000;
      24063: inst = 32'hfe0a9ea;
      24064: inst = 32'h5be00000;
      24065: inst = 32'h244c8000;
      24066: inst = 32'h24428800;
      24067: inst = 32'h8620000;
      24068: inst = 32'h2a0e0002;
      24069: inst = 32'h294f0003;
      24070: inst = 32'h11200000;
      24071: inst = 32'hd205e0b;
      24072: inst = 32'h13e00000;
      24073: inst = 32'hfe0a9ea;
      24074: inst = 32'h5be00000;
      24075: inst = 32'h244c8000;
      24076: inst = 32'h24428800;
      24077: inst = 32'h8620000;
      24078: inst = 32'h2a0e000a;
      24079: inst = 32'h294f0004;
      24080: inst = 32'h11200000;
      24081: inst = 32'hd205e15;
      24082: inst = 32'h13e00000;
      24083: inst = 32'hfe0a9ea;
      24084: inst = 32'h5be00000;
      24085: inst = 32'h244c8000;
      24086: inst = 32'h24428800;
      24087: inst = 32'h8620000;
      24088: inst = 32'h2a0e0002;
      24089: inst = 32'h294f0004;
      24090: inst = 32'h11200000;
      24091: inst = 32'hd205e1f;
      24092: inst = 32'h13e00000;
      24093: inst = 32'hfe0a9ea;
      24094: inst = 32'h5be00000;
      24095: inst = 32'h244c8000;
      24096: inst = 32'h24428800;
      24097: inst = 32'h8620000;
      24098: inst = 32'h2a0e000a;
      24099: inst = 32'h294f0005;
      24100: inst = 32'h11200000;
      24101: inst = 32'hd205e29;
      24102: inst = 32'h13e00000;
      24103: inst = 32'hfe0a9ea;
      24104: inst = 32'h5be00000;
      24105: inst = 32'h244c8000;
      24106: inst = 32'h24428800;
      24107: inst = 32'h8620000;
      24108: inst = 32'h2a0e0009;
      24109: inst = 32'h294f0005;
      24110: inst = 32'h11200000;
      24111: inst = 32'hd205e33;
      24112: inst = 32'h13e00000;
      24113: inst = 32'hfe0a9ea;
      24114: inst = 32'h5be00000;
      24115: inst = 32'h244c8000;
      24116: inst = 32'h24428800;
      24117: inst = 32'h8620000;
      24118: inst = 32'h2a0e000a;
      24119: inst = 32'h294f0006;
      24120: inst = 32'h11200000;
      24121: inst = 32'hd205e3d;
      24122: inst = 32'h13e00000;
      24123: inst = 32'hfe0a9ea;
      24124: inst = 32'h5be00000;
      24125: inst = 32'h244c8000;
      24126: inst = 32'h24428800;
      24127: inst = 32'h8620000;
      24128: inst = 32'h2a0e0009;
      24129: inst = 32'h294f0006;
      24130: inst = 32'h11200000;
      24131: inst = 32'hd205e47;
      24132: inst = 32'h13e00000;
      24133: inst = 32'hfe0a9ea;
      24134: inst = 32'h5be00000;
      24135: inst = 32'h244c8000;
      24136: inst = 32'h24428800;
      24137: inst = 32'h8620000;
      24138: inst = 32'hc60d42c;
      24139: inst = 32'h2a0e0008;
      24140: inst = 32'h294f0002;
      24141: inst = 32'h11200000;
      24142: inst = 32'hd205e52;
      24143: inst = 32'h13e00000;
      24144: inst = 32'hfe0a9ea;
      24145: inst = 32'h5be00000;
      24146: inst = 32'h244c8000;
      24147: inst = 32'h24428800;
      24148: inst = 32'h8620000;
      24149: inst = 32'h2a0e0007;
      24150: inst = 32'h294f0002;
      24151: inst = 32'h11200000;
      24152: inst = 32'hd205e5c;
      24153: inst = 32'h13e00000;
      24154: inst = 32'hfe0a9ea;
      24155: inst = 32'h5be00000;
      24156: inst = 32'h244c8000;
      24157: inst = 32'h24428800;
      24158: inst = 32'h8620000;
      24159: inst = 32'h2a0e0006;
      24160: inst = 32'h294f0002;
      24161: inst = 32'h11200000;
      24162: inst = 32'hd205e66;
      24163: inst = 32'h13e00000;
      24164: inst = 32'hfe0a9ea;
      24165: inst = 32'h5be00000;
      24166: inst = 32'h244c8000;
      24167: inst = 32'h24428800;
      24168: inst = 32'h8620000;
      24169: inst = 32'h2a0e0005;
      24170: inst = 32'h294f0002;
      24171: inst = 32'h11200000;
      24172: inst = 32'hd205e70;
      24173: inst = 32'h13e00000;
      24174: inst = 32'hfe0a9ea;
      24175: inst = 32'h5be00000;
      24176: inst = 32'h244c8000;
      24177: inst = 32'h24428800;
      24178: inst = 32'h8620000;
      24179: inst = 32'h2a0e0004;
      24180: inst = 32'h294f0002;
      24181: inst = 32'h11200000;
      24182: inst = 32'hd205e7a;
      24183: inst = 32'h13e00000;
      24184: inst = 32'hfe0a9ea;
      24185: inst = 32'h5be00000;
      24186: inst = 32'h244c8000;
      24187: inst = 32'h24428800;
      24188: inst = 32'h8620000;
      24189: inst = 32'h2a0e0003;
      24190: inst = 32'h294f0002;
      24191: inst = 32'h11200000;
      24192: inst = 32'hd205e84;
      24193: inst = 32'h13e00000;
      24194: inst = 32'hfe0a9ea;
      24195: inst = 32'h5be00000;
      24196: inst = 32'h244c8000;
      24197: inst = 32'h24428800;
      24198: inst = 32'h8620000;
      24199: inst = 32'h2a0e0002;
      24200: inst = 32'h294f0002;
      24201: inst = 32'h11200000;
      24202: inst = 32'hd205e8e;
      24203: inst = 32'h13e00000;
      24204: inst = 32'hfe0a9ea;
      24205: inst = 32'h5be00000;
      24206: inst = 32'h244c8000;
      24207: inst = 32'h24428800;
      24208: inst = 32'h8620000;
      24209: inst = 32'h2a0e0001;
      24210: inst = 32'h294f0002;
      24211: inst = 32'h11200000;
      24212: inst = 32'hd205e98;
      24213: inst = 32'h13e00000;
      24214: inst = 32'hfe0a9ea;
      24215: inst = 32'h5be00000;
      24216: inst = 32'h244c8000;
      24217: inst = 32'h24428800;
      24218: inst = 32'h8620000;
      24219: inst = 32'h2a0e0008;
      24220: inst = 32'h294f0005;
      24221: inst = 32'h11200000;
      24222: inst = 32'hd205ea2;
      24223: inst = 32'h13e00000;
      24224: inst = 32'hfe0a9ea;
      24225: inst = 32'h5be00000;
      24226: inst = 32'h244c8000;
      24227: inst = 32'h24428800;
      24228: inst = 32'h8620000;
      24229: inst = 32'h2a0e0008;
      24230: inst = 32'h294f0006;
      24231: inst = 32'h11200000;
      24232: inst = 32'hd205eac;
      24233: inst = 32'h13e00000;
      24234: inst = 32'hfe0a9ea;
      24235: inst = 32'h5be00000;
      24236: inst = 32'h244c8000;
      24237: inst = 32'h24428800;
      24238: inst = 32'h8620000;
      24239: inst = 32'h2a0e0007;
      24240: inst = 32'h294f000b;
      24241: inst = 32'h11200000;
      24242: inst = 32'hd205eb6;
      24243: inst = 32'h13e00000;
      24244: inst = 32'hfe0a9ea;
      24245: inst = 32'h5be00000;
      24246: inst = 32'h244c8000;
      24247: inst = 32'h24428800;
      24248: inst = 32'h8620000;
      24249: inst = 32'h2a0e0004;
      24250: inst = 32'h294f000b;
      24251: inst = 32'h11200000;
      24252: inst = 32'hd205ec0;
      24253: inst = 32'h13e00000;
      24254: inst = 32'hfe0a9ea;
      24255: inst = 32'h5be00000;
      24256: inst = 32'h244c8000;
      24257: inst = 32'h24428800;
      24258: inst = 32'h8620000;
      24259: inst = 32'hc60f4ce;
      24260: inst = 32'h2a0e0009;
      24261: inst = 32'h294f0003;
      24262: inst = 32'h11200000;
      24263: inst = 32'hd205ecb;
      24264: inst = 32'h13e00000;
      24265: inst = 32'hfe0a9ea;
      24266: inst = 32'h5be00000;
      24267: inst = 32'h244c8000;
      24268: inst = 32'h24428800;
      24269: inst = 32'h8620000;
      24270: inst = 32'h2a0e0008;
      24271: inst = 32'h294f0003;
      24272: inst = 32'h11200000;
      24273: inst = 32'hd205ed5;
      24274: inst = 32'h13e00000;
      24275: inst = 32'hfe0a9ea;
      24276: inst = 32'h5be00000;
      24277: inst = 32'h244c8000;
      24278: inst = 32'h24428800;
      24279: inst = 32'h8620000;
      24280: inst = 32'h2a0e0007;
      24281: inst = 32'h294f0003;
      24282: inst = 32'h11200000;
      24283: inst = 32'hd205edf;
      24284: inst = 32'h13e00000;
      24285: inst = 32'hfe0a9ea;
      24286: inst = 32'h5be00000;
      24287: inst = 32'h244c8000;
      24288: inst = 32'h24428800;
      24289: inst = 32'h8620000;
      24290: inst = 32'h2a0e0006;
      24291: inst = 32'h294f0003;
      24292: inst = 32'h11200000;
      24293: inst = 32'hd205ee9;
      24294: inst = 32'h13e00000;
      24295: inst = 32'hfe0a9ea;
      24296: inst = 32'h5be00000;
      24297: inst = 32'h244c8000;
      24298: inst = 32'h24428800;
      24299: inst = 32'h8620000;
      24300: inst = 32'h2a0e0005;
      24301: inst = 32'h294f0003;
      24302: inst = 32'h11200000;
      24303: inst = 32'hd205ef3;
      24304: inst = 32'h13e00000;
      24305: inst = 32'hfe0a9ea;
      24306: inst = 32'h5be00000;
      24307: inst = 32'h244c8000;
      24308: inst = 32'h24428800;
      24309: inst = 32'h8620000;
      24310: inst = 32'h2a0e0004;
      24311: inst = 32'h294f0003;
      24312: inst = 32'h11200000;
      24313: inst = 32'hd205efd;
      24314: inst = 32'h13e00000;
      24315: inst = 32'hfe0a9ea;
      24316: inst = 32'h5be00000;
      24317: inst = 32'h244c8000;
      24318: inst = 32'h24428800;
      24319: inst = 32'h8620000;
      24320: inst = 32'h2a0e0003;
      24321: inst = 32'h294f0003;
      24322: inst = 32'h11200000;
      24323: inst = 32'hd205f07;
      24324: inst = 32'h13e00000;
      24325: inst = 32'hfe0a9ea;
      24326: inst = 32'h5be00000;
      24327: inst = 32'h244c8000;
      24328: inst = 32'h24428800;
      24329: inst = 32'h8620000;
      24330: inst = 32'h2a0e0001;
      24331: inst = 32'h294f0003;
      24332: inst = 32'h11200000;
      24333: inst = 32'hd205f11;
      24334: inst = 32'h13e00000;
      24335: inst = 32'hfe0a9ea;
      24336: inst = 32'h5be00000;
      24337: inst = 32'h244c8000;
      24338: inst = 32'h24428800;
      24339: inst = 32'h8620000;
      24340: inst = 32'h2a0e0009;
      24341: inst = 32'h294f0004;
      24342: inst = 32'h11200000;
      24343: inst = 32'hd205f1b;
      24344: inst = 32'h13e00000;
      24345: inst = 32'hfe0a9ea;
      24346: inst = 32'h5be00000;
      24347: inst = 32'h244c8000;
      24348: inst = 32'h24428800;
      24349: inst = 32'h8620000;
      24350: inst = 32'h2a0e0008;
      24351: inst = 32'h294f0004;
      24352: inst = 32'h11200000;
      24353: inst = 32'hd205f25;
      24354: inst = 32'h13e00000;
      24355: inst = 32'hfe0a9ea;
      24356: inst = 32'h5be00000;
      24357: inst = 32'h244c8000;
      24358: inst = 32'h24428800;
      24359: inst = 32'h8620000;
      24360: inst = 32'h2a0e0007;
      24361: inst = 32'h294f0004;
      24362: inst = 32'h11200000;
      24363: inst = 32'hd205f2f;
      24364: inst = 32'h13e00000;
      24365: inst = 32'hfe0a9ea;
      24366: inst = 32'h5be00000;
      24367: inst = 32'h244c8000;
      24368: inst = 32'h24428800;
      24369: inst = 32'h8620000;
      24370: inst = 32'h2a0e0006;
      24371: inst = 32'h294f0004;
      24372: inst = 32'h11200000;
      24373: inst = 32'hd205f39;
      24374: inst = 32'h13e00000;
      24375: inst = 32'hfe0a9ea;
      24376: inst = 32'h5be00000;
      24377: inst = 32'h244c8000;
      24378: inst = 32'h24428800;
      24379: inst = 32'h8620000;
      24380: inst = 32'h2a0e0005;
      24381: inst = 32'h294f0004;
      24382: inst = 32'h11200000;
      24383: inst = 32'hd205f43;
      24384: inst = 32'h13e00000;
      24385: inst = 32'hfe0a9ea;
      24386: inst = 32'h5be00000;
      24387: inst = 32'h244c8000;
      24388: inst = 32'h24428800;
      24389: inst = 32'h8620000;
      24390: inst = 32'h2a0e0004;
      24391: inst = 32'h294f0004;
      24392: inst = 32'h11200000;
      24393: inst = 32'hd205f4d;
      24394: inst = 32'h13e00000;
      24395: inst = 32'hfe0a9ea;
      24396: inst = 32'h5be00000;
      24397: inst = 32'h244c8000;
      24398: inst = 32'h24428800;
      24399: inst = 32'h8620000;
      24400: inst = 32'h2a0e0003;
      24401: inst = 32'h294f0004;
      24402: inst = 32'h11200000;
      24403: inst = 32'hd205f57;
      24404: inst = 32'h13e00000;
      24405: inst = 32'hfe0a9ea;
      24406: inst = 32'h5be00000;
      24407: inst = 32'h244c8000;
      24408: inst = 32'h24428800;
      24409: inst = 32'h8620000;
      24410: inst = 32'h2a0e0001;
      24411: inst = 32'h294f0004;
      24412: inst = 32'h11200000;
      24413: inst = 32'hd205f61;
      24414: inst = 32'h13e00000;
      24415: inst = 32'hfe0a9ea;
      24416: inst = 32'h5be00000;
      24417: inst = 32'h244c8000;
      24418: inst = 32'h24428800;
      24419: inst = 32'h8620000;
      24420: inst = 32'h2a0e0007;
      24421: inst = 32'h294f0005;
      24422: inst = 32'h11200000;
      24423: inst = 32'hd205f6b;
      24424: inst = 32'h13e00000;
      24425: inst = 32'hfe0a9ea;
      24426: inst = 32'h5be00000;
      24427: inst = 32'h244c8000;
      24428: inst = 32'h24428800;
      24429: inst = 32'h8620000;
      24430: inst = 32'h2a0e0006;
      24431: inst = 32'h294f0005;
      24432: inst = 32'h11200000;
      24433: inst = 32'hd205f75;
      24434: inst = 32'h13e00000;
      24435: inst = 32'hfe0a9ea;
      24436: inst = 32'h5be00000;
      24437: inst = 32'h244c8000;
      24438: inst = 32'h24428800;
      24439: inst = 32'h8620000;
      24440: inst = 32'h2a0e0005;
      24441: inst = 32'h294f0005;
      24442: inst = 32'h11200000;
      24443: inst = 32'hd205f7f;
      24444: inst = 32'h13e00000;
      24445: inst = 32'hfe0a9ea;
      24446: inst = 32'h5be00000;
      24447: inst = 32'h244c8000;
      24448: inst = 32'h24428800;
      24449: inst = 32'h8620000;
      24450: inst = 32'h2a0e0004;
      24451: inst = 32'h294f0005;
      24452: inst = 32'h11200000;
      24453: inst = 32'hd205f89;
      24454: inst = 32'h13e00000;
      24455: inst = 32'hfe0a9ea;
      24456: inst = 32'h5be00000;
      24457: inst = 32'h244c8000;
      24458: inst = 32'h24428800;
      24459: inst = 32'h8620000;
      24460: inst = 32'h2a0e0003;
      24461: inst = 32'h294f0005;
      24462: inst = 32'h11200000;
      24463: inst = 32'hd205f93;
      24464: inst = 32'h13e00000;
      24465: inst = 32'hfe0a9ea;
      24466: inst = 32'h5be00000;
      24467: inst = 32'h244c8000;
      24468: inst = 32'h24428800;
      24469: inst = 32'h8620000;
      24470: inst = 32'h2a0e0002;
      24471: inst = 32'h294f0005;
      24472: inst = 32'h11200000;
      24473: inst = 32'hd205f9d;
      24474: inst = 32'h13e00000;
      24475: inst = 32'hfe0a9ea;
      24476: inst = 32'h5be00000;
      24477: inst = 32'h244c8000;
      24478: inst = 32'h24428800;
      24479: inst = 32'h8620000;
      24480: inst = 32'h2a0e0001;
      24481: inst = 32'h294f0005;
      24482: inst = 32'h11200000;
      24483: inst = 32'hd205fa7;
      24484: inst = 32'h13e00000;
      24485: inst = 32'hfe0a9ea;
      24486: inst = 32'h5be00000;
      24487: inst = 32'h244c8000;
      24488: inst = 32'h24428800;
      24489: inst = 32'h8620000;
      24490: inst = 32'h2a0e0007;
      24491: inst = 32'h294f0006;
      24492: inst = 32'h11200000;
      24493: inst = 32'hd205fb1;
      24494: inst = 32'h13e00000;
      24495: inst = 32'hfe0a9ea;
      24496: inst = 32'h5be00000;
      24497: inst = 32'h244c8000;
      24498: inst = 32'h24428800;
      24499: inst = 32'h8620000;
      24500: inst = 32'h2a0e0006;
      24501: inst = 32'h294f0006;
      24502: inst = 32'h11200000;
      24503: inst = 32'hd205fbb;
      24504: inst = 32'h13e00000;
      24505: inst = 32'hfe0a9ea;
      24506: inst = 32'h5be00000;
      24507: inst = 32'h244c8000;
      24508: inst = 32'h24428800;
      24509: inst = 32'h8620000;
      24510: inst = 32'h2a0e0005;
      24511: inst = 32'h294f0006;
      24512: inst = 32'h11200000;
      24513: inst = 32'hd205fc5;
      24514: inst = 32'h13e00000;
      24515: inst = 32'hfe0a9ea;
      24516: inst = 32'h5be00000;
      24517: inst = 32'h244c8000;
      24518: inst = 32'h24428800;
      24519: inst = 32'h8620000;
      24520: inst = 32'h2a0e0004;
      24521: inst = 32'h294f0006;
      24522: inst = 32'h11200000;
      24523: inst = 32'hd205fcf;
      24524: inst = 32'h13e00000;
      24525: inst = 32'hfe0a9ea;
      24526: inst = 32'h5be00000;
      24527: inst = 32'h244c8000;
      24528: inst = 32'h24428800;
      24529: inst = 32'h8620000;
      24530: inst = 32'h2a0e0003;
      24531: inst = 32'h294f0006;
      24532: inst = 32'h11200000;
      24533: inst = 32'hd205fd9;
      24534: inst = 32'h13e00000;
      24535: inst = 32'hfe0a9ea;
      24536: inst = 32'h5be00000;
      24537: inst = 32'h244c8000;
      24538: inst = 32'h24428800;
      24539: inst = 32'h8620000;
      24540: inst = 32'h2a0e0002;
      24541: inst = 32'h294f0006;
      24542: inst = 32'h11200000;
      24543: inst = 32'hd205fe3;
      24544: inst = 32'h13e00000;
      24545: inst = 32'hfe0a9ea;
      24546: inst = 32'h5be00000;
      24547: inst = 32'h244c8000;
      24548: inst = 32'h24428800;
      24549: inst = 32'h8620000;
      24550: inst = 32'h2a0e0001;
      24551: inst = 32'h294f0006;
      24552: inst = 32'h11200000;
      24553: inst = 32'hd205fed;
      24554: inst = 32'h13e00000;
      24555: inst = 32'hfe0a9ea;
      24556: inst = 32'h5be00000;
      24557: inst = 32'h244c8000;
      24558: inst = 32'h24428800;
      24559: inst = 32'h8620000;
      24560: inst = 32'h2a0e0006;
      24561: inst = 32'h294f0008;
      24562: inst = 32'h11200000;
      24563: inst = 32'hd205ff7;
      24564: inst = 32'h13e00000;
      24565: inst = 32'hfe0a9ea;
      24566: inst = 32'h5be00000;
      24567: inst = 32'h244c8000;
      24568: inst = 32'h24428800;
      24569: inst = 32'h8620000;
      24570: inst = 32'h2a0e0002;
      24571: inst = 32'h294f0008;
      24572: inst = 32'h11200000;
      24573: inst = 32'hd206001;
      24574: inst = 32'h13e00000;
      24575: inst = 32'hfe0a9ea;
      24576: inst = 32'h5be00000;
      24577: inst = 32'h244c8000;
      24578: inst = 32'h24428800;
      24579: inst = 32'h8620000;
      24580: inst = 32'h2a0e0006;
      24581: inst = 32'h294f0009;
      24582: inst = 32'h11200000;
      24583: inst = 32'hd20600b;
      24584: inst = 32'h13e00000;
      24585: inst = 32'hfe0a9ea;
      24586: inst = 32'h5be00000;
      24587: inst = 32'h244c8000;
      24588: inst = 32'h24428800;
      24589: inst = 32'h8620000;
      24590: inst = 32'hc607841;
      24591: inst = 32'h2a0e0008;
      24592: inst = 32'h294f0007;
      24593: inst = 32'h11200000;
      24594: inst = 32'hd206016;
      24595: inst = 32'h13e00000;
      24596: inst = 32'hfe0a9ea;
      24597: inst = 32'h5be00000;
      24598: inst = 32'h244c8000;
      24599: inst = 32'h24428800;
      24600: inst = 32'h8620000;
      24601: inst = 32'h2a0e0008;
      24602: inst = 32'h294f0008;
      24603: inst = 32'h11200000;
      24604: inst = 32'hd206020;
      24605: inst = 32'h13e00000;
      24606: inst = 32'hfe0a9ea;
      24607: inst = 32'h5be00000;
      24608: inst = 32'h244c8000;
      24609: inst = 32'h24428800;
      24610: inst = 32'h8620000;
      24611: inst = 32'hc60a000;
      24612: inst = 32'h2a0e0007;
      24613: inst = 32'h294f0007;
      24614: inst = 32'h11200000;
      24615: inst = 32'hd20602b;
      24616: inst = 32'h13e00000;
      24617: inst = 32'hfe0a9ea;
      24618: inst = 32'h5be00000;
      24619: inst = 32'h244c8000;
      24620: inst = 32'h24428800;
      24621: inst = 32'h8620000;
      24622: inst = 32'h2a0e0006;
      24623: inst = 32'h294f0007;
      24624: inst = 32'h11200000;
      24625: inst = 32'hd206035;
      24626: inst = 32'h13e00000;
      24627: inst = 32'hfe0a9ea;
      24628: inst = 32'h5be00000;
      24629: inst = 32'h244c8000;
      24630: inst = 32'h24428800;
      24631: inst = 32'h8620000;
      24632: inst = 32'h2a0e0005;
      24633: inst = 32'h294f0007;
      24634: inst = 32'h11200000;
      24635: inst = 32'hd20603f;
      24636: inst = 32'h13e00000;
      24637: inst = 32'hfe0a9ea;
      24638: inst = 32'h5be00000;
      24639: inst = 32'h244c8000;
      24640: inst = 32'h24428800;
      24641: inst = 32'h8620000;
      24642: inst = 32'h2a0e0004;
      24643: inst = 32'h294f0007;
      24644: inst = 32'h11200000;
      24645: inst = 32'hd206049;
      24646: inst = 32'h13e00000;
      24647: inst = 32'hfe0a9ea;
      24648: inst = 32'h5be00000;
      24649: inst = 32'h244c8000;
      24650: inst = 32'h24428800;
      24651: inst = 32'h8620000;
      24652: inst = 32'h2a0e0003;
      24653: inst = 32'h294f0007;
      24654: inst = 32'h11200000;
      24655: inst = 32'hd206053;
      24656: inst = 32'h13e00000;
      24657: inst = 32'hfe0a9ea;
      24658: inst = 32'h5be00000;
      24659: inst = 32'h244c8000;
      24660: inst = 32'h24428800;
      24661: inst = 32'h8620000;
      24662: inst = 32'h2a0e0007;
      24663: inst = 32'h294f0008;
      24664: inst = 32'h11200000;
      24665: inst = 32'hd20605d;
      24666: inst = 32'h13e00000;
      24667: inst = 32'hfe0a9ea;
      24668: inst = 32'h5be00000;
      24669: inst = 32'h244c8000;
      24670: inst = 32'h24428800;
      24671: inst = 32'h8620000;
      24672: inst = 32'h2a0e0005;
      24673: inst = 32'h294f0008;
      24674: inst = 32'h11200000;
      24675: inst = 32'hd206067;
      24676: inst = 32'h13e00000;
      24677: inst = 32'hfe0a9ea;
      24678: inst = 32'h5be00000;
      24679: inst = 32'h244c8000;
      24680: inst = 32'h24428800;
      24681: inst = 32'h8620000;
      24682: inst = 32'h2a0e0004;
      24683: inst = 32'h294f0008;
      24684: inst = 32'h11200000;
      24685: inst = 32'hd206071;
      24686: inst = 32'h13e00000;
      24687: inst = 32'hfe0a9ea;
      24688: inst = 32'h5be00000;
      24689: inst = 32'h244c8000;
      24690: inst = 32'h24428800;
      24691: inst = 32'h8620000;
      24692: inst = 32'h2a0e0003;
      24693: inst = 32'h294f0008;
      24694: inst = 32'h11200000;
      24695: inst = 32'hd20607b;
      24696: inst = 32'h13e00000;
      24697: inst = 32'hfe0a9ea;
      24698: inst = 32'h5be00000;
      24699: inst = 32'h244c8000;
      24700: inst = 32'h24428800;
      24701: inst = 32'h8620000;
      24702: inst = 32'h2a0e0008;
      24703: inst = 32'h294f0009;
      24704: inst = 32'h11200000;
      24705: inst = 32'hd206085;
      24706: inst = 32'h13e00000;
      24707: inst = 32'hfe0a9ea;
      24708: inst = 32'h5be00000;
      24709: inst = 32'h244c8000;
      24710: inst = 32'h24428800;
      24711: inst = 32'h8620000;
      24712: inst = 32'h2a0e0007;
      24713: inst = 32'h294f0009;
      24714: inst = 32'h11200000;
      24715: inst = 32'hd20608f;
      24716: inst = 32'h13e00000;
      24717: inst = 32'hfe0a9ea;
      24718: inst = 32'h5be00000;
      24719: inst = 32'h244c8000;
      24720: inst = 32'h24428800;
      24721: inst = 32'h8620000;
      24722: inst = 32'h2a0e0005;
      24723: inst = 32'h294f0009;
      24724: inst = 32'h11200000;
      24725: inst = 32'hd206099;
      24726: inst = 32'h13e00000;
      24727: inst = 32'hfe0a9ea;
      24728: inst = 32'h5be00000;
      24729: inst = 32'h244c8000;
      24730: inst = 32'h24428800;
      24731: inst = 32'h8620000;
      24732: inst = 32'h2a0e0004;
      24733: inst = 32'h294f0009;
      24734: inst = 32'h11200000;
      24735: inst = 32'hd2060a3;
      24736: inst = 32'h13e00000;
      24737: inst = 32'hfe0a9ea;
      24738: inst = 32'h5be00000;
      24739: inst = 32'h244c8000;
      24740: inst = 32'h24428800;
      24741: inst = 32'h8620000;
      24742: inst = 32'h2a0e0003;
      24743: inst = 32'h294f0009;
      24744: inst = 32'h11200000;
      24745: inst = 32'hd2060ad;
      24746: inst = 32'h13e00000;
      24747: inst = 32'hfe0a9ea;
      24748: inst = 32'h5be00000;
      24749: inst = 32'h244c8000;
      24750: inst = 32'h24428800;
      24751: inst = 32'h8620000;
      24752: inst = 32'hc6010ac;
      24753: inst = 32'h2a0e0008;
      24754: inst = 32'h294f000a;
      24755: inst = 32'h11200000;
      24756: inst = 32'hd2060b8;
      24757: inst = 32'h13e00000;
      24758: inst = 32'hfe0a9ea;
      24759: inst = 32'h5be00000;
      24760: inst = 32'h244c8000;
      24761: inst = 32'h24428800;
      24762: inst = 32'h8620000;
      24763: inst = 32'h2a0e0007;
      24764: inst = 32'h294f000a;
      24765: inst = 32'h11200000;
      24766: inst = 32'hd2060c2;
      24767: inst = 32'h13e00000;
      24768: inst = 32'hfe0a9ea;
      24769: inst = 32'h5be00000;
      24770: inst = 32'h244c8000;
      24771: inst = 32'h24428800;
      24772: inst = 32'h8620000;
      24773: inst = 32'h2a0e0006;
      24774: inst = 32'h294f000a;
      24775: inst = 32'h11200000;
      24776: inst = 32'hd2060cc;
      24777: inst = 32'h13e00000;
      24778: inst = 32'hfe0a9ea;
      24779: inst = 32'h5be00000;
      24780: inst = 32'h244c8000;
      24781: inst = 32'h24428800;
      24782: inst = 32'h8620000;
      24783: inst = 32'h2a0e0005;
      24784: inst = 32'h294f000a;
      24785: inst = 32'h11200000;
      24786: inst = 32'hd2060d6;
      24787: inst = 32'h13e00000;
      24788: inst = 32'hfe0a9ea;
      24789: inst = 32'h5be00000;
      24790: inst = 32'h244c8000;
      24791: inst = 32'h24428800;
      24792: inst = 32'h8620000;
      24793: inst = 32'h2a0e0004;
      24794: inst = 32'h294f000a;
      24795: inst = 32'h11200000;
      24796: inst = 32'hd2060e0;
      24797: inst = 32'h13e00000;
      24798: inst = 32'hfe0a9ea;
      24799: inst = 32'h5be00000;
      24800: inst = 32'h244c8000;
      24801: inst = 32'h24428800;
      24802: inst = 32'h8620000;
      24803: inst = 32'h2a0e0003;
      24804: inst = 32'h294f000a;
      24805: inst = 32'h11200000;
      24806: inst = 32'hd2060ea;
      24807: inst = 32'h13e00000;
      24808: inst = 32'hfe0a9ea;
      24809: inst = 32'h5be00000;
      24810: inst = 32'h244c8000;
      24811: inst = 32'h24428800;
      24812: inst = 32'h8620000;
      24813: inst = 32'h13e00000;
      24814: inst = 32'hfe060f4;
      24815: inst = 32'h20200001;
      24816: inst = 32'h5be00000;
      24817: inst = 32'h13e00000;
      24818: inst = 32'hfe060f7;
      24819: inst = 32'h5be00000;
      24820: inst = 32'h13e00000;
      24821: inst = 32'hfe060f7;
      24822: inst = 32'h5be00000;
      24823: inst = 32'h58000000;
      24824: inst = 32'h10408000;
      24825: inst = 32'hc400002;
      24826: inst = 32'h4420000;
      24827: inst = 32'h10600000;
      24828: inst = 32'hc600010;
      24829: inst = 32'h38421800;
      24830: inst = 32'h4042000f;
      24831: inst = 32'h1c40000f;
      24832: inst = 32'h58000000;
      24833: inst = 32'h58200000;
      24834: inst = 32'hc206b50;
      24835: inst = 32'h10408000;
      24836: inst = 32'hc403fe0;
      24837: inst = 32'h8220000;
      24838: inst = 32'h10408000;
      24839: inst = 32'hc403fe1;
      24840: inst = 32'h8220000;
      24841: inst = 32'h10408000;
      24842: inst = 32'hc403fe2;
      24843: inst = 32'h8220000;
      24844: inst = 32'h10408000;
      24845: inst = 32'hc403ff5;
      24846: inst = 32'h8220000;
      24847: inst = 32'h10408000;
      24848: inst = 32'hc403ff8;
      24849: inst = 32'h8220000;
      24850: inst = 32'h10408000;
      24851: inst = 32'hc403ff9;
      24852: inst = 32'h8220000;
      24853: inst = 32'h10408000;
      24854: inst = 32'hc403ffd;
      24855: inst = 32'h8220000;
      24856: inst = 32'h10408000;
      24857: inst = 32'hc403ffe;
      24858: inst = 32'h8220000;
      24859: inst = 32'h10408000;
      24860: inst = 32'hc403fff;
      24861: inst = 32'h8220000;
      24862: inst = 32'h10408000;
      24863: inst = 32'hc404000;
      24864: inst = 32'h8220000;
      24865: inst = 32'h10408000;
      24866: inst = 32'hc404001;
      24867: inst = 32'h8220000;
      24868: inst = 32'h10408000;
      24869: inst = 32'hc404002;
      24870: inst = 32'h8220000;
      24871: inst = 32'h10408000;
      24872: inst = 32'hc404003;
      24873: inst = 32'h8220000;
      24874: inst = 32'h10408000;
      24875: inst = 32'hc404004;
      24876: inst = 32'h8220000;
      24877: inst = 32'h10408000;
      24878: inst = 32'hc404005;
      24879: inst = 32'h8220000;
      24880: inst = 32'h10408000;
      24881: inst = 32'hc404006;
      24882: inst = 32'h8220000;
      24883: inst = 32'h10408000;
      24884: inst = 32'hc404007;
      24885: inst = 32'h8220000;
      24886: inst = 32'h10408000;
      24887: inst = 32'hc404008;
      24888: inst = 32'h8220000;
      24889: inst = 32'h10408000;
      24890: inst = 32'hc404009;
      24891: inst = 32'h8220000;
      24892: inst = 32'h10408000;
      24893: inst = 32'hc40400a;
      24894: inst = 32'h8220000;
      24895: inst = 32'h10408000;
      24896: inst = 32'hc40400b;
      24897: inst = 32'h8220000;
      24898: inst = 32'h10408000;
      24899: inst = 32'hc40400c;
      24900: inst = 32'h8220000;
      24901: inst = 32'h10408000;
      24902: inst = 32'hc40400d;
      24903: inst = 32'h8220000;
      24904: inst = 32'h10408000;
      24905: inst = 32'hc40400e;
      24906: inst = 32'h8220000;
      24907: inst = 32'h10408000;
      24908: inst = 32'hc40400f;
      24909: inst = 32'h8220000;
      24910: inst = 32'h10408000;
      24911: inst = 32'hc404010;
      24912: inst = 32'h8220000;
      24913: inst = 32'h10408000;
      24914: inst = 32'hc404011;
      24915: inst = 32'h8220000;
      24916: inst = 32'h10408000;
      24917: inst = 32'hc404012;
      24918: inst = 32'h8220000;
      24919: inst = 32'h10408000;
      24920: inst = 32'hc404013;
      24921: inst = 32'h8220000;
      24922: inst = 32'h10408000;
      24923: inst = 32'hc404014;
      24924: inst = 32'h8220000;
      24925: inst = 32'h10408000;
      24926: inst = 32'hc404015;
      24927: inst = 32'h8220000;
      24928: inst = 32'h10408000;
      24929: inst = 32'hc404016;
      24930: inst = 32'h8220000;
      24931: inst = 32'h10408000;
      24932: inst = 32'hc404017;
      24933: inst = 32'h8220000;
      24934: inst = 32'h10408000;
      24935: inst = 32'hc404018;
      24936: inst = 32'h8220000;
      24937: inst = 32'h10408000;
      24938: inst = 32'hc404019;
      24939: inst = 32'h8220000;
      24940: inst = 32'h10408000;
      24941: inst = 32'hc40401a;
      24942: inst = 32'h8220000;
      24943: inst = 32'h10408000;
      24944: inst = 32'hc40401b;
      24945: inst = 32'h8220000;
      24946: inst = 32'h10408000;
      24947: inst = 32'hc40401c;
      24948: inst = 32'h8220000;
      24949: inst = 32'h10408000;
      24950: inst = 32'hc40401d;
      24951: inst = 32'h8220000;
      24952: inst = 32'h10408000;
      24953: inst = 32'hc40401e;
      24954: inst = 32'h8220000;
      24955: inst = 32'h10408000;
      24956: inst = 32'hc40401f;
      24957: inst = 32'h8220000;
      24958: inst = 32'h10408000;
      24959: inst = 32'hc404020;
      24960: inst = 32'h8220000;
      24961: inst = 32'h10408000;
      24962: inst = 32'hc404021;
      24963: inst = 32'h8220000;
      24964: inst = 32'h10408000;
      24965: inst = 32'hc404022;
      24966: inst = 32'h8220000;
      24967: inst = 32'h10408000;
      24968: inst = 32'hc404023;
      24969: inst = 32'h8220000;
      24970: inst = 32'h10408000;
      24971: inst = 32'hc404024;
      24972: inst = 32'h8220000;
      24973: inst = 32'h10408000;
      24974: inst = 32'hc404025;
      24975: inst = 32'h8220000;
      24976: inst = 32'h10408000;
      24977: inst = 32'hc404026;
      24978: inst = 32'h8220000;
      24979: inst = 32'h10408000;
      24980: inst = 32'hc404027;
      24981: inst = 32'h8220000;
      24982: inst = 32'h10408000;
      24983: inst = 32'hc404028;
      24984: inst = 32'h8220000;
      24985: inst = 32'h10408000;
      24986: inst = 32'hc404029;
      24987: inst = 32'h8220000;
      24988: inst = 32'h10408000;
      24989: inst = 32'hc40402a;
      24990: inst = 32'h8220000;
      24991: inst = 32'h10408000;
      24992: inst = 32'hc40402b;
      24993: inst = 32'h8220000;
      24994: inst = 32'h10408000;
      24995: inst = 32'hc40402c;
      24996: inst = 32'h8220000;
      24997: inst = 32'h10408000;
      24998: inst = 32'hc40402d;
      24999: inst = 32'h8220000;
      25000: inst = 32'h10408000;
      25001: inst = 32'hc40402e;
      25002: inst = 32'h8220000;
      25003: inst = 32'h10408000;
      25004: inst = 32'hc40402f;
      25005: inst = 32'h8220000;
      25006: inst = 32'h10408000;
      25007: inst = 32'hc404030;
      25008: inst = 32'h8220000;
      25009: inst = 32'h10408000;
      25010: inst = 32'hc404031;
      25011: inst = 32'h8220000;
      25012: inst = 32'h10408000;
      25013: inst = 32'hc404032;
      25014: inst = 32'h8220000;
      25015: inst = 32'h10408000;
      25016: inst = 32'hc404033;
      25017: inst = 32'h8220000;
      25018: inst = 32'h10408000;
      25019: inst = 32'hc404034;
      25020: inst = 32'h8220000;
      25021: inst = 32'h10408000;
      25022: inst = 32'hc404035;
      25023: inst = 32'h8220000;
      25024: inst = 32'h10408000;
      25025: inst = 32'hc404036;
      25026: inst = 32'h8220000;
      25027: inst = 32'h10408000;
      25028: inst = 32'hc404037;
      25029: inst = 32'h8220000;
      25030: inst = 32'h10408000;
      25031: inst = 32'hc404038;
      25032: inst = 32'h8220000;
      25033: inst = 32'h10408000;
      25034: inst = 32'hc404039;
      25035: inst = 32'h8220000;
      25036: inst = 32'h10408000;
      25037: inst = 32'hc40403a;
      25038: inst = 32'h8220000;
      25039: inst = 32'h10408000;
      25040: inst = 32'hc40403b;
      25041: inst = 32'h8220000;
      25042: inst = 32'h10408000;
      25043: inst = 32'hc40403c;
      25044: inst = 32'h8220000;
      25045: inst = 32'h10408000;
      25046: inst = 32'hc40403d;
      25047: inst = 32'h8220000;
      25048: inst = 32'h10408000;
      25049: inst = 32'hc40403e;
      25050: inst = 32'h8220000;
      25051: inst = 32'h10408000;
      25052: inst = 32'hc40403f;
      25053: inst = 32'h8220000;
      25054: inst = 32'h10408000;
      25055: inst = 32'hc404040;
      25056: inst = 32'h8220000;
      25057: inst = 32'h10408000;
      25058: inst = 32'hc404041;
      25059: inst = 32'h8220000;
      25060: inst = 32'h10408000;
      25061: inst = 32'hc404042;
      25062: inst = 32'h8220000;
      25063: inst = 32'h10408000;
      25064: inst = 32'hc404054;
      25065: inst = 32'h8220000;
      25066: inst = 32'h10408000;
      25067: inst = 32'hc404057;
      25068: inst = 32'h8220000;
      25069: inst = 32'h10408000;
      25070: inst = 32'hc404058;
      25071: inst = 32'h8220000;
      25072: inst = 32'h10408000;
      25073: inst = 32'hc40405c;
      25074: inst = 32'h8220000;
      25075: inst = 32'h10408000;
      25076: inst = 32'hc40405d;
      25077: inst = 32'h8220000;
      25078: inst = 32'h10408000;
      25079: inst = 32'hc40405e;
      25080: inst = 32'h8220000;
      25081: inst = 32'h10408000;
      25082: inst = 32'hc40405f;
      25083: inst = 32'h8220000;
      25084: inst = 32'h10408000;
      25085: inst = 32'hc404060;
      25086: inst = 32'h8220000;
      25087: inst = 32'h10408000;
      25088: inst = 32'hc404061;
      25089: inst = 32'h8220000;
      25090: inst = 32'h10408000;
      25091: inst = 32'hc404062;
      25092: inst = 32'h8220000;
      25093: inst = 32'h10408000;
      25094: inst = 32'hc404063;
      25095: inst = 32'h8220000;
      25096: inst = 32'h10408000;
      25097: inst = 32'hc404064;
      25098: inst = 32'h8220000;
      25099: inst = 32'h10408000;
      25100: inst = 32'hc404065;
      25101: inst = 32'h8220000;
      25102: inst = 32'h10408000;
      25103: inst = 32'hc404066;
      25104: inst = 32'h8220000;
      25105: inst = 32'h10408000;
      25106: inst = 32'hc404067;
      25107: inst = 32'h8220000;
      25108: inst = 32'h10408000;
      25109: inst = 32'hc404068;
      25110: inst = 32'h8220000;
      25111: inst = 32'h10408000;
      25112: inst = 32'hc404069;
      25113: inst = 32'h8220000;
      25114: inst = 32'h10408000;
      25115: inst = 32'hc40406a;
      25116: inst = 32'h8220000;
      25117: inst = 32'h10408000;
      25118: inst = 32'hc40406b;
      25119: inst = 32'h8220000;
      25120: inst = 32'h10408000;
      25121: inst = 32'hc40406c;
      25122: inst = 32'h8220000;
      25123: inst = 32'h10408000;
      25124: inst = 32'hc40406d;
      25125: inst = 32'h8220000;
      25126: inst = 32'h10408000;
      25127: inst = 32'hc40406e;
      25128: inst = 32'h8220000;
      25129: inst = 32'h10408000;
      25130: inst = 32'hc40406f;
      25131: inst = 32'h8220000;
      25132: inst = 32'h10408000;
      25133: inst = 32'hc404070;
      25134: inst = 32'h8220000;
      25135: inst = 32'h10408000;
      25136: inst = 32'hc404071;
      25137: inst = 32'h8220000;
      25138: inst = 32'h10408000;
      25139: inst = 32'hc404072;
      25140: inst = 32'h8220000;
      25141: inst = 32'h10408000;
      25142: inst = 32'hc404073;
      25143: inst = 32'h8220000;
      25144: inst = 32'h10408000;
      25145: inst = 32'hc404074;
      25146: inst = 32'h8220000;
      25147: inst = 32'h10408000;
      25148: inst = 32'hc404075;
      25149: inst = 32'h8220000;
      25150: inst = 32'h10408000;
      25151: inst = 32'hc404076;
      25152: inst = 32'h8220000;
      25153: inst = 32'h10408000;
      25154: inst = 32'hc404077;
      25155: inst = 32'h8220000;
      25156: inst = 32'h10408000;
      25157: inst = 32'hc404078;
      25158: inst = 32'h8220000;
      25159: inst = 32'h10408000;
      25160: inst = 32'hc404079;
      25161: inst = 32'h8220000;
      25162: inst = 32'h10408000;
      25163: inst = 32'hc40407a;
      25164: inst = 32'h8220000;
      25165: inst = 32'h10408000;
      25166: inst = 32'hc40407b;
      25167: inst = 32'h8220000;
      25168: inst = 32'h10408000;
      25169: inst = 32'hc40407c;
      25170: inst = 32'h8220000;
      25171: inst = 32'h10408000;
      25172: inst = 32'hc40407d;
      25173: inst = 32'h8220000;
      25174: inst = 32'h10408000;
      25175: inst = 32'hc40407e;
      25176: inst = 32'h8220000;
      25177: inst = 32'h10408000;
      25178: inst = 32'hc40407f;
      25179: inst = 32'h8220000;
      25180: inst = 32'h10408000;
      25181: inst = 32'hc404080;
      25182: inst = 32'h8220000;
      25183: inst = 32'h10408000;
      25184: inst = 32'hc404081;
      25185: inst = 32'h8220000;
      25186: inst = 32'h10408000;
      25187: inst = 32'hc404082;
      25188: inst = 32'h8220000;
      25189: inst = 32'h10408000;
      25190: inst = 32'hc404083;
      25191: inst = 32'h8220000;
      25192: inst = 32'h10408000;
      25193: inst = 32'hc404084;
      25194: inst = 32'h8220000;
      25195: inst = 32'h10408000;
      25196: inst = 32'hc404085;
      25197: inst = 32'h8220000;
      25198: inst = 32'h10408000;
      25199: inst = 32'hc404086;
      25200: inst = 32'h8220000;
      25201: inst = 32'h10408000;
      25202: inst = 32'hc404087;
      25203: inst = 32'h8220000;
      25204: inst = 32'h10408000;
      25205: inst = 32'hc404088;
      25206: inst = 32'h8220000;
      25207: inst = 32'h10408000;
      25208: inst = 32'hc404089;
      25209: inst = 32'h8220000;
      25210: inst = 32'h10408000;
      25211: inst = 32'hc40408a;
      25212: inst = 32'h8220000;
      25213: inst = 32'h10408000;
      25214: inst = 32'hc40408b;
      25215: inst = 32'h8220000;
      25216: inst = 32'h10408000;
      25217: inst = 32'hc40408c;
      25218: inst = 32'h8220000;
      25219: inst = 32'h10408000;
      25220: inst = 32'hc40408d;
      25221: inst = 32'h8220000;
      25222: inst = 32'h10408000;
      25223: inst = 32'hc40408e;
      25224: inst = 32'h8220000;
      25225: inst = 32'h10408000;
      25226: inst = 32'hc40408f;
      25227: inst = 32'h8220000;
      25228: inst = 32'h10408000;
      25229: inst = 32'hc404090;
      25230: inst = 32'h8220000;
      25231: inst = 32'h10408000;
      25232: inst = 32'hc404091;
      25233: inst = 32'h8220000;
      25234: inst = 32'h10408000;
      25235: inst = 32'hc404092;
      25236: inst = 32'h8220000;
      25237: inst = 32'h10408000;
      25238: inst = 32'hc404093;
      25239: inst = 32'h8220000;
      25240: inst = 32'h10408000;
      25241: inst = 32'hc404094;
      25242: inst = 32'h8220000;
      25243: inst = 32'h10408000;
      25244: inst = 32'hc404095;
      25245: inst = 32'h8220000;
      25246: inst = 32'h10408000;
      25247: inst = 32'hc404096;
      25248: inst = 32'h8220000;
      25249: inst = 32'h10408000;
      25250: inst = 32'hc404097;
      25251: inst = 32'h8220000;
      25252: inst = 32'h10408000;
      25253: inst = 32'hc404098;
      25254: inst = 32'h8220000;
      25255: inst = 32'h10408000;
      25256: inst = 32'hc404099;
      25257: inst = 32'h8220000;
      25258: inst = 32'h10408000;
      25259: inst = 32'hc40409a;
      25260: inst = 32'h8220000;
      25261: inst = 32'h10408000;
      25262: inst = 32'hc40409b;
      25263: inst = 32'h8220000;
      25264: inst = 32'h10408000;
      25265: inst = 32'hc40409c;
      25266: inst = 32'h8220000;
      25267: inst = 32'h10408000;
      25268: inst = 32'hc40409d;
      25269: inst = 32'h8220000;
      25270: inst = 32'h10408000;
      25271: inst = 32'hc40409e;
      25272: inst = 32'h8220000;
      25273: inst = 32'h10408000;
      25274: inst = 32'hc40409f;
      25275: inst = 32'h8220000;
      25276: inst = 32'h10408000;
      25277: inst = 32'hc4040a0;
      25278: inst = 32'h8220000;
      25279: inst = 32'h10408000;
      25280: inst = 32'hc4040a1;
      25281: inst = 32'h8220000;
      25282: inst = 32'h10408000;
      25283: inst = 32'hc4040a2;
      25284: inst = 32'h8220000;
      25285: inst = 32'h10408000;
      25286: inst = 32'hc4040af;
      25287: inst = 32'h8220000;
      25288: inst = 32'h10408000;
      25289: inst = 32'hc4040b2;
      25290: inst = 32'h8220000;
      25291: inst = 32'h10408000;
      25292: inst = 32'hc4040b7;
      25293: inst = 32'h8220000;
      25294: inst = 32'h10408000;
      25295: inst = 32'hc4040b8;
      25296: inst = 32'h8220000;
      25297: inst = 32'h10408000;
      25298: inst = 32'hc4040bb;
      25299: inst = 32'h8220000;
      25300: inst = 32'h10408000;
      25301: inst = 32'hc4040bc;
      25302: inst = 32'h8220000;
      25303: inst = 32'h10408000;
      25304: inst = 32'hc4040bd;
      25305: inst = 32'h8220000;
      25306: inst = 32'h10408000;
      25307: inst = 32'hc4040be;
      25308: inst = 32'h8220000;
      25309: inst = 32'h10408000;
      25310: inst = 32'hc4040bf;
      25311: inst = 32'h8220000;
      25312: inst = 32'h10408000;
      25313: inst = 32'hc4040c0;
      25314: inst = 32'h8220000;
      25315: inst = 32'h10408000;
      25316: inst = 32'hc4040c1;
      25317: inst = 32'h8220000;
      25318: inst = 32'h10408000;
      25319: inst = 32'hc4040c2;
      25320: inst = 32'h8220000;
      25321: inst = 32'h10408000;
      25322: inst = 32'hc4040c3;
      25323: inst = 32'h8220000;
      25324: inst = 32'h10408000;
      25325: inst = 32'hc4040c4;
      25326: inst = 32'h8220000;
      25327: inst = 32'h10408000;
      25328: inst = 32'hc4040c5;
      25329: inst = 32'h8220000;
      25330: inst = 32'h10408000;
      25331: inst = 32'hc4040c6;
      25332: inst = 32'h8220000;
      25333: inst = 32'h10408000;
      25334: inst = 32'hc4040c7;
      25335: inst = 32'h8220000;
      25336: inst = 32'h10408000;
      25337: inst = 32'hc4040c8;
      25338: inst = 32'h8220000;
      25339: inst = 32'h10408000;
      25340: inst = 32'hc4040c9;
      25341: inst = 32'h8220000;
      25342: inst = 32'h10408000;
      25343: inst = 32'hc4040ca;
      25344: inst = 32'h8220000;
      25345: inst = 32'h10408000;
      25346: inst = 32'hc4040cb;
      25347: inst = 32'h8220000;
      25348: inst = 32'h10408000;
      25349: inst = 32'hc4040cc;
      25350: inst = 32'h8220000;
      25351: inst = 32'h10408000;
      25352: inst = 32'hc4040cd;
      25353: inst = 32'h8220000;
      25354: inst = 32'h10408000;
      25355: inst = 32'hc4040ce;
      25356: inst = 32'h8220000;
      25357: inst = 32'h10408000;
      25358: inst = 32'hc4040cf;
      25359: inst = 32'h8220000;
      25360: inst = 32'h10408000;
      25361: inst = 32'hc4040d0;
      25362: inst = 32'h8220000;
      25363: inst = 32'h10408000;
      25364: inst = 32'hc4040d1;
      25365: inst = 32'h8220000;
      25366: inst = 32'h10408000;
      25367: inst = 32'hc4040d2;
      25368: inst = 32'h8220000;
      25369: inst = 32'h10408000;
      25370: inst = 32'hc4040d3;
      25371: inst = 32'h8220000;
      25372: inst = 32'h10408000;
      25373: inst = 32'hc4040d4;
      25374: inst = 32'h8220000;
      25375: inst = 32'h10408000;
      25376: inst = 32'hc4040d5;
      25377: inst = 32'h8220000;
      25378: inst = 32'h10408000;
      25379: inst = 32'hc4040d6;
      25380: inst = 32'h8220000;
      25381: inst = 32'h10408000;
      25382: inst = 32'hc4040d7;
      25383: inst = 32'h8220000;
      25384: inst = 32'h10408000;
      25385: inst = 32'hc4040d8;
      25386: inst = 32'h8220000;
      25387: inst = 32'h10408000;
      25388: inst = 32'hc4040d9;
      25389: inst = 32'h8220000;
      25390: inst = 32'h10408000;
      25391: inst = 32'hc4040da;
      25392: inst = 32'h8220000;
      25393: inst = 32'h10408000;
      25394: inst = 32'hc4040db;
      25395: inst = 32'h8220000;
      25396: inst = 32'h10408000;
      25397: inst = 32'hc4040dc;
      25398: inst = 32'h8220000;
      25399: inst = 32'h10408000;
      25400: inst = 32'hc4040dd;
      25401: inst = 32'h8220000;
      25402: inst = 32'h10408000;
      25403: inst = 32'hc4040de;
      25404: inst = 32'h8220000;
      25405: inst = 32'h10408000;
      25406: inst = 32'hc4040df;
      25407: inst = 32'h8220000;
      25408: inst = 32'h10408000;
      25409: inst = 32'hc4040e0;
      25410: inst = 32'h8220000;
      25411: inst = 32'h10408000;
      25412: inst = 32'hc4040e1;
      25413: inst = 32'h8220000;
      25414: inst = 32'h10408000;
      25415: inst = 32'hc4040e2;
      25416: inst = 32'h8220000;
      25417: inst = 32'h10408000;
      25418: inst = 32'hc4040e3;
      25419: inst = 32'h8220000;
      25420: inst = 32'h10408000;
      25421: inst = 32'hc4040e4;
      25422: inst = 32'h8220000;
      25423: inst = 32'h10408000;
      25424: inst = 32'hc4040e5;
      25425: inst = 32'h8220000;
      25426: inst = 32'h10408000;
      25427: inst = 32'hc4040e6;
      25428: inst = 32'h8220000;
      25429: inst = 32'h10408000;
      25430: inst = 32'hc4040e7;
      25431: inst = 32'h8220000;
      25432: inst = 32'h10408000;
      25433: inst = 32'hc4040e8;
      25434: inst = 32'h8220000;
      25435: inst = 32'h10408000;
      25436: inst = 32'hc4040e9;
      25437: inst = 32'h8220000;
      25438: inst = 32'h10408000;
      25439: inst = 32'hc4040ea;
      25440: inst = 32'h8220000;
      25441: inst = 32'h10408000;
      25442: inst = 32'hc4040eb;
      25443: inst = 32'h8220000;
      25444: inst = 32'h10408000;
      25445: inst = 32'hc4040ec;
      25446: inst = 32'h8220000;
      25447: inst = 32'h10408000;
      25448: inst = 32'hc4040ed;
      25449: inst = 32'h8220000;
      25450: inst = 32'h10408000;
      25451: inst = 32'hc4040ee;
      25452: inst = 32'h8220000;
      25453: inst = 32'h10408000;
      25454: inst = 32'hc4040ef;
      25455: inst = 32'h8220000;
      25456: inst = 32'h10408000;
      25457: inst = 32'hc4040f0;
      25458: inst = 32'h8220000;
      25459: inst = 32'h10408000;
      25460: inst = 32'hc4040f1;
      25461: inst = 32'h8220000;
      25462: inst = 32'h10408000;
      25463: inst = 32'hc4040f2;
      25464: inst = 32'h8220000;
      25465: inst = 32'h10408000;
      25466: inst = 32'hc4040f3;
      25467: inst = 32'h8220000;
      25468: inst = 32'h10408000;
      25469: inst = 32'hc4040f4;
      25470: inst = 32'h8220000;
      25471: inst = 32'h10408000;
      25472: inst = 32'hc4040f5;
      25473: inst = 32'h8220000;
      25474: inst = 32'h10408000;
      25475: inst = 32'hc4040f6;
      25476: inst = 32'h8220000;
      25477: inst = 32'h10408000;
      25478: inst = 32'hc4040f7;
      25479: inst = 32'h8220000;
      25480: inst = 32'h10408000;
      25481: inst = 32'hc4040f8;
      25482: inst = 32'h8220000;
      25483: inst = 32'h10408000;
      25484: inst = 32'hc4040f9;
      25485: inst = 32'h8220000;
      25486: inst = 32'h10408000;
      25487: inst = 32'hc4040fa;
      25488: inst = 32'h8220000;
      25489: inst = 32'h10408000;
      25490: inst = 32'hc4040fb;
      25491: inst = 32'h8220000;
      25492: inst = 32'h10408000;
      25493: inst = 32'hc4040fc;
      25494: inst = 32'h8220000;
      25495: inst = 32'h10408000;
      25496: inst = 32'hc4040fd;
      25497: inst = 32'h8220000;
      25498: inst = 32'h10408000;
      25499: inst = 32'hc4040fe;
      25500: inst = 32'h8220000;
      25501: inst = 32'h10408000;
      25502: inst = 32'hc4040ff;
      25503: inst = 32'h8220000;
      25504: inst = 32'h10408000;
      25505: inst = 32'hc404100;
      25506: inst = 32'h8220000;
      25507: inst = 32'h10408000;
      25508: inst = 32'hc404101;
      25509: inst = 32'h8220000;
      25510: inst = 32'h10408000;
      25511: inst = 32'hc404102;
      25512: inst = 32'h8220000;
      25513: inst = 32'h10408000;
      25514: inst = 32'hc40414c;
      25515: inst = 32'h8220000;
      25516: inst = 32'h10408000;
      25517: inst = 32'hc40414d;
      25518: inst = 32'h8220000;
      25519: inst = 32'h10408000;
      25520: inst = 32'hc40414e;
      25521: inst = 32'h8220000;
      25522: inst = 32'h10408000;
      25523: inst = 32'hc40415d;
      25524: inst = 32'h8220000;
      25525: inst = 32'h10408000;
      25526: inst = 32'hc40415e;
      25527: inst = 32'h8220000;
      25528: inst = 32'h10408000;
      25529: inst = 32'hc40415f;
      25530: inst = 32'h8220000;
      25531: inst = 32'h10408000;
      25532: inst = 32'hc404160;
      25533: inst = 32'h8220000;
      25534: inst = 32'h10408000;
      25535: inst = 32'hc404161;
      25536: inst = 32'h8220000;
      25537: inst = 32'h10408000;
      25538: inst = 32'hc404162;
      25539: inst = 32'h8220000;
      25540: inst = 32'h10408000;
      25541: inst = 32'hc4041ac;
      25542: inst = 32'h8220000;
      25543: inst = 32'h10408000;
      25544: inst = 32'hc4041ad;
      25545: inst = 32'h8220000;
      25546: inst = 32'h10408000;
      25547: inst = 32'hc4041ae;
      25548: inst = 32'h8220000;
      25549: inst = 32'h10408000;
      25550: inst = 32'hc4041bd;
      25551: inst = 32'h8220000;
      25552: inst = 32'h10408000;
      25553: inst = 32'hc4041be;
      25554: inst = 32'h8220000;
      25555: inst = 32'h10408000;
      25556: inst = 32'hc4041bf;
      25557: inst = 32'h8220000;
      25558: inst = 32'h10408000;
      25559: inst = 32'hc4041c0;
      25560: inst = 32'h8220000;
      25561: inst = 32'h10408000;
      25562: inst = 32'hc4041c1;
      25563: inst = 32'h8220000;
      25564: inst = 32'h10408000;
      25565: inst = 32'hc4041c2;
      25566: inst = 32'h8220000;
      25567: inst = 32'h10408000;
      25568: inst = 32'hc40420c;
      25569: inst = 32'h8220000;
      25570: inst = 32'h10408000;
      25571: inst = 32'hc40420d;
      25572: inst = 32'h8220000;
      25573: inst = 32'h10408000;
      25574: inst = 32'hc40420e;
      25575: inst = 32'h8220000;
      25576: inst = 32'h10408000;
      25577: inst = 32'hc40421d;
      25578: inst = 32'h8220000;
      25579: inst = 32'h10408000;
      25580: inst = 32'hc40421e;
      25581: inst = 32'h8220000;
      25582: inst = 32'h10408000;
      25583: inst = 32'hc40421f;
      25584: inst = 32'h8220000;
      25585: inst = 32'h10408000;
      25586: inst = 32'hc404220;
      25587: inst = 32'h8220000;
      25588: inst = 32'h10408000;
      25589: inst = 32'hc404221;
      25590: inst = 32'h8220000;
      25591: inst = 32'h10408000;
      25592: inst = 32'hc404222;
      25593: inst = 32'h8220000;
      25594: inst = 32'h10408000;
      25595: inst = 32'hc40426c;
      25596: inst = 32'h8220000;
      25597: inst = 32'h10408000;
      25598: inst = 32'hc40426d;
      25599: inst = 32'h8220000;
      25600: inst = 32'h10408000;
      25601: inst = 32'hc40426e;
      25602: inst = 32'h8220000;
      25603: inst = 32'h10408000;
      25604: inst = 32'hc40427d;
      25605: inst = 32'h8220000;
      25606: inst = 32'h10408000;
      25607: inst = 32'hc40427e;
      25608: inst = 32'h8220000;
      25609: inst = 32'h10408000;
      25610: inst = 32'hc40427f;
      25611: inst = 32'h8220000;
      25612: inst = 32'h10408000;
      25613: inst = 32'hc404280;
      25614: inst = 32'h8220000;
      25615: inst = 32'h10408000;
      25616: inst = 32'hc404281;
      25617: inst = 32'h8220000;
      25618: inst = 32'h10408000;
      25619: inst = 32'hc404282;
      25620: inst = 32'h8220000;
      25621: inst = 32'h10408000;
      25622: inst = 32'hc4042cc;
      25623: inst = 32'h8220000;
      25624: inst = 32'h10408000;
      25625: inst = 32'hc4042cd;
      25626: inst = 32'h8220000;
      25627: inst = 32'h10408000;
      25628: inst = 32'hc4042ce;
      25629: inst = 32'h8220000;
      25630: inst = 32'h10408000;
      25631: inst = 32'hc4042dd;
      25632: inst = 32'h8220000;
      25633: inst = 32'h10408000;
      25634: inst = 32'hc4042de;
      25635: inst = 32'h8220000;
      25636: inst = 32'h10408000;
      25637: inst = 32'hc4042df;
      25638: inst = 32'h8220000;
      25639: inst = 32'h10408000;
      25640: inst = 32'hc4042e0;
      25641: inst = 32'h8220000;
      25642: inst = 32'h10408000;
      25643: inst = 32'hc4042e1;
      25644: inst = 32'h8220000;
      25645: inst = 32'h10408000;
      25646: inst = 32'hc4042e2;
      25647: inst = 32'h8220000;
      25648: inst = 32'h10408000;
      25649: inst = 32'hc40432c;
      25650: inst = 32'h8220000;
      25651: inst = 32'h10408000;
      25652: inst = 32'hc40432d;
      25653: inst = 32'h8220000;
      25654: inst = 32'h10408000;
      25655: inst = 32'hc40432e;
      25656: inst = 32'h8220000;
      25657: inst = 32'h10408000;
      25658: inst = 32'hc40433d;
      25659: inst = 32'h8220000;
      25660: inst = 32'h10408000;
      25661: inst = 32'hc40433e;
      25662: inst = 32'h8220000;
      25663: inst = 32'h10408000;
      25664: inst = 32'hc40433f;
      25665: inst = 32'h8220000;
      25666: inst = 32'h10408000;
      25667: inst = 32'hc404340;
      25668: inst = 32'h8220000;
      25669: inst = 32'h10408000;
      25670: inst = 32'hc404341;
      25671: inst = 32'h8220000;
      25672: inst = 32'h10408000;
      25673: inst = 32'hc404342;
      25674: inst = 32'h8220000;
      25675: inst = 32'h10408000;
      25676: inst = 32'hc40438c;
      25677: inst = 32'h8220000;
      25678: inst = 32'h10408000;
      25679: inst = 32'hc40438d;
      25680: inst = 32'h8220000;
      25681: inst = 32'h10408000;
      25682: inst = 32'hc40438e;
      25683: inst = 32'h8220000;
      25684: inst = 32'h10408000;
      25685: inst = 32'hc40439d;
      25686: inst = 32'h8220000;
      25687: inst = 32'h10408000;
      25688: inst = 32'hc40439e;
      25689: inst = 32'h8220000;
      25690: inst = 32'h10408000;
      25691: inst = 32'hc40439f;
      25692: inst = 32'h8220000;
      25693: inst = 32'h10408000;
      25694: inst = 32'hc4043a0;
      25695: inst = 32'h8220000;
      25696: inst = 32'h10408000;
      25697: inst = 32'hc4043a1;
      25698: inst = 32'h8220000;
      25699: inst = 32'h10408000;
      25700: inst = 32'hc4043a2;
      25701: inst = 32'h8220000;
      25702: inst = 32'h10408000;
      25703: inst = 32'hc4043ec;
      25704: inst = 32'h8220000;
      25705: inst = 32'h10408000;
      25706: inst = 32'hc4043ed;
      25707: inst = 32'h8220000;
      25708: inst = 32'h10408000;
      25709: inst = 32'hc4043ee;
      25710: inst = 32'h8220000;
      25711: inst = 32'h10408000;
      25712: inst = 32'hc4043fd;
      25713: inst = 32'h8220000;
      25714: inst = 32'h10408000;
      25715: inst = 32'hc4043fe;
      25716: inst = 32'h8220000;
      25717: inst = 32'h10408000;
      25718: inst = 32'hc4043ff;
      25719: inst = 32'h8220000;
      25720: inst = 32'h10408000;
      25721: inst = 32'hc404400;
      25722: inst = 32'h8220000;
      25723: inst = 32'h10408000;
      25724: inst = 32'hc404401;
      25725: inst = 32'h8220000;
      25726: inst = 32'h10408000;
      25727: inst = 32'hc404402;
      25728: inst = 32'h8220000;
      25729: inst = 32'h10408000;
      25730: inst = 32'hc40444c;
      25731: inst = 32'h8220000;
      25732: inst = 32'h10408000;
      25733: inst = 32'hc40444d;
      25734: inst = 32'h8220000;
      25735: inst = 32'h10408000;
      25736: inst = 32'hc40444e;
      25737: inst = 32'h8220000;
      25738: inst = 32'h10408000;
      25739: inst = 32'hc40445d;
      25740: inst = 32'h8220000;
      25741: inst = 32'h10408000;
      25742: inst = 32'hc40445e;
      25743: inst = 32'h8220000;
      25744: inst = 32'h10408000;
      25745: inst = 32'hc40445f;
      25746: inst = 32'h8220000;
      25747: inst = 32'h10408000;
      25748: inst = 32'hc404460;
      25749: inst = 32'h8220000;
      25750: inst = 32'h10408000;
      25751: inst = 32'hc404461;
      25752: inst = 32'h8220000;
      25753: inst = 32'h10408000;
      25754: inst = 32'hc404462;
      25755: inst = 32'h8220000;
      25756: inst = 32'h10408000;
      25757: inst = 32'hc4044ac;
      25758: inst = 32'h8220000;
      25759: inst = 32'h10408000;
      25760: inst = 32'hc4044ad;
      25761: inst = 32'h8220000;
      25762: inst = 32'h10408000;
      25763: inst = 32'hc4044ae;
      25764: inst = 32'h8220000;
      25765: inst = 32'h10408000;
      25766: inst = 32'hc4044bd;
      25767: inst = 32'h8220000;
      25768: inst = 32'h10408000;
      25769: inst = 32'hc4044be;
      25770: inst = 32'h8220000;
      25771: inst = 32'h10408000;
      25772: inst = 32'hc4044bf;
      25773: inst = 32'h8220000;
      25774: inst = 32'h10408000;
      25775: inst = 32'hc4044c0;
      25776: inst = 32'h8220000;
      25777: inst = 32'h10408000;
      25778: inst = 32'hc4044c1;
      25779: inst = 32'h8220000;
      25780: inst = 32'h10408000;
      25781: inst = 32'hc4044c2;
      25782: inst = 32'h8220000;
      25783: inst = 32'h10408000;
      25784: inst = 32'hc40450c;
      25785: inst = 32'h8220000;
      25786: inst = 32'h10408000;
      25787: inst = 32'hc40450d;
      25788: inst = 32'h8220000;
      25789: inst = 32'h10408000;
      25790: inst = 32'hc40450e;
      25791: inst = 32'h8220000;
      25792: inst = 32'h10408000;
      25793: inst = 32'hc40451d;
      25794: inst = 32'h8220000;
      25795: inst = 32'h10408000;
      25796: inst = 32'hc40451e;
      25797: inst = 32'h8220000;
      25798: inst = 32'h10408000;
      25799: inst = 32'hc40451f;
      25800: inst = 32'h8220000;
      25801: inst = 32'h10408000;
      25802: inst = 32'hc404520;
      25803: inst = 32'h8220000;
      25804: inst = 32'h10408000;
      25805: inst = 32'hc404521;
      25806: inst = 32'h8220000;
      25807: inst = 32'h10408000;
      25808: inst = 32'hc404522;
      25809: inst = 32'h8220000;
      25810: inst = 32'h10408000;
      25811: inst = 32'hc40456c;
      25812: inst = 32'h8220000;
      25813: inst = 32'h10408000;
      25814: inst = 32'hc40456d;
      25815: inst = 32'h8220000;
      25816: inst = 32'h10408000;
      25817: inst = 32'hc40456e;
      25818: inst = 32'h8220000;
      25819: inst = 32'h10408000;
      25820: inst = 32'hc40457d;
      25821: inst = 32'h8220000;
      25822: inst = 32'h10408000;
      25823: inst = 32'hc40457e;
      25824: inst = 32'h8220000;
      25825: inst = 32'h10408000;
      25826: inst = 32'hc40457f;
      25827: inst = 32'h8220000;
      25828: inst = 32'h10408000;
      25829: inst = 32'hc404580;
      25830: inst = 32'h8220000;
      25831: inst = 32'h10408000;
      25832: inst = 32'hc404581;
      25833: inst = 32'h8220000;
      25834: inst = 32'h10408000;
      25835: inst = 32'hc404582;
      25836: inst = 32'h8220000;
      25837: inst = 32'h10408000;
      25838: inst = 32'hc4045cc;
      25839: inst = 32'h8220000;
      25840: inst = 32'h10408000;
      25841: inst = 32'hc4045cd;
      25842: inst = 32'h8220000;
      25843: inst = 32'h10408000;
      25844: inst = 32'hc4045ce;
      25845: inst = 32'h8220000;
      25846: inst = 32'h10408000;
      25847: inst = 32'hc4045dd;
      25848: inst = 32'h8220000;
      25849: inst = 32'h10408000;
      25850: inst = 32'hc4045de;
      25851: inst = 32'h8220000;
      25852: inst = 32'h10408000;
      25853: inst = 32'hc4045df;
      25854: inst = 32'h8220000;
      25855: inst = 32'h10408000;
      25856: inst = 32'hc4045e0;
      25857: inst = 32'h8220000;
      25858: inst = 32'h10408000;
      25859: inst = 32'hc4045e1;
      25860: inst = 32'h8220000;
      25861: inst = 32'h10408000;
      25862: inst = 32'hc4045e2;
      25863: inst = 32'h8220000;
      25864: inst = 32'h10408000;
      25865: inst = 32'hc40462c;
      25866: inst = 32'h8220000;
      25867: inst = 32'h10408000;
      25868: inst = 32'hc40462d;
      25869: inst = 32'h8220000;
      25870: inst = 32'h10408000;
      25871: inst = 32'hc40462e;
      25872: inst = 32'h8220000;
      25873: inst = 32'h10408000;
      25874: inst = 32'hc40463d;
      25875: inst = 32'h8220000;
      25876: inst = 32'h10408000;
      25877: inst = 32'hc40463e;
      25878: inst = 32'h8220000;
      25879: inst = 32'h10408000;
      25880: inst = 32'hc40463f;
      25881: inst = 32'h8220000;
      25882: inst = 32'h10408000;
      25883: inst = 32'hc404640;
      25884: inst = 32'h8220000;
      25885: inst = 32'h10408000;
      25886: inst = 32'hc404641;
      25887: inst = 32'h8220000;
      25888: inst = 32'h10408000;
      25889: inst = 32'hc404642;
      25890: inst = 32'h8220000;
      25891: inst = 32'h10408000;
      25892: inst = 32'hc40464e;
      25893: inst = 32'h8220000;
      25894: inst = 32'h10408000;
      25895: inst = 32'hc40464f;
      25896: inst = 32'h8220000;
      25897: inst = 32'h10408000;
      25898: inst = 32'hc404650;
      25899: inst = 32'h8220000;
      25900: inst = 32'h10408000;
      25901: inst = 32'hc404651;
      25902: inst = 32'h8220000;
      25903: inst = 32'h10408000;
      25904: inst = 32'hc404652;
      25905: inst = 32'h8220000;
      25906: inst = 32'h10408000;
      25907: inst = 32'hc404653;
      25908: inst = 32'h8220000;
      25909: inst = 32'h10408000;
      25910: inst = 32'hc404654;
      25911: inst = 32'h8220000;
      25912: inst = 32'h10408000;
      25913: inst = 32'hc404655;
      25914: inst = 32'h8220000;
      25915: inst = 32'h10408000;
      25916: inst = 32'hc404656;
      25917: inst = 32'h8220000;
      25918: inst = 32'h10408000;
      25919: inst = 32'hc404657;
      25920: inst = 32'h8220000;
      25921: inst = 32'h10408000;
      25922: inst = 32'hc404658;
      25923: inst = 32'h8220000;
      25924: inst = 32'h10408000;
      25925: inst = 32'hc404659;
      25926: inst = 32'h8220000;
      25927: inst = 32'h10408000;
      25928: inst = 32'hc40465a;
      25929: inst = 32'h8220000;
      25930: inst = 32'h10408000;
      25931: inst = 32'hc40465b;
      25932: inst = 32'h8220000;
      25933: inst = 32'h10408000;
      25934: inst = 32'hc40465c;
      25935: inst = 32'h8220000;
      25936: inst = 32'h10408000;
      25937: inst = 32'hc40465d;
      25938: inst = 32'h8220000;
      25939: inst = 32'h10408000;
      25940: inst = 32'hc40465e;
      25941: inst = 32'h8220000;
      25942: inst = 32'h10408000;
      25943: inst = 32'hc40465f;
      25944: inst = 32'h8220000;
      25945: inst = 32'h10408000;
      25946: inst = 32'hc404660;
      25947: inst = 32'h8220000;
      25948: inst = 32'h10408000;
      25949: inst = 32'hc404661;
      25950: inst = 32'h8220000;
      25951: inst = 32'h10408000;
      25952: inst = 32'hc404662;
      25953: inst = 32'h8220000;
      25954: inst = 32'h10408000;
      25955: inst = 32'hc404663;
      25956: inst = 32'h8220000;
      25957: inst = 32'h10408000;
      25958: inst = 32'hc404664;
      25959: inst = 32'h8220000;
      25960: inst = 32'h10408000;
      25961: inst = 32'hc404665;
      25962: inst = 32'h8220000;
      25963: inst = 32'h10408000;
      25964: inst = 32'hc404666;
      25965: inst = 32'h8220000;
      25966: inst = 32'h10408000;
      25967: inst = 32'hc404667;
      25968: inst = 32'h8220000;
      25969: inst = 32'h10408000;
      25970: inst = 32'hc404668;
      25971: inst = 32'h8220000;
      25972: inst = 32'h10408000;
      25973: inst = 32'hc404669;
      25974: inst = 32'h8220000;
      25975: inst = 32'h10408000;
      25976: inst = 32'hc40466e;
      25977: inst = 32'h8220000;
      25978: inst = 32'h10408000;
      25979: inst = 32'hc40466f;
      25980: inst = 32'h8220000;
      25981: inst = 32'h10408000;
      25982: inst = 32'hc404673;
      25983: inst = 32'h8220000;
      25984: inst = 32'h10408000;
      25985: inst = 32'hc404676;
      25986: inst = 32'h8220000;
      25987: inst = 32'h10408000;
      25988: inst = 32'hc40468c;
      25989: inst = 32'h8220000;
      25990: inst = 32'h10408000;
      25991: inst = 32'hc40468d;
      25992: inst = 32'h8220000;
      25993: inst = 32'h10408000;
      25994: inst = 32'hc40468e;
      25995: inst = 32'h8220000;
      25996: inst = 32'h10408000;
      25997: inst = 32'hc40469d;
      25998: inst = 32'h8220000;
      25999: inst = 32'h10408000;
      26000: inst = 32'hc40469e;
      26001: inst = 32'h8220000;
      26002: inst = 32'h10408000;
      26003: inst = 32'hc40469f;
      26004: inst = 32'h8220000;
      26005: inst = 32'h10408000;
      26006: inst = 32'hc4046a0;
      26007: inst = 32'h8220000;
      26008: inst = 32'h10408000;
      26009: inst = 32'hc4046a1;
      26010: inst = 32'h8220000;
      26011: inst = 32'h10408000;
      26012: inst = 32'hc4046a2;
      26013: inst = 32'h8220000;
      26014: inst = 32'h10408000;
      26015: inst = 32'hc4046ae;
      26016: inst = 32'h8220000;
      26017: inst = 32'h10408000;
      26018: inst = 32'hc4046af;
      26019: inst = 32'h8220000;
      26020: inst = 32'h10408000;
      26021: inst = 32'hc4046b0;
      26022: inst = 32'h8220000;
      26023: inst = 32'h10408000;
      26024: inst = 32'hc4046b1;
      26025: inst = 32'h8220000;
      26026: inst = 32'h10408000;
      26027: inst = 32'hc4046b2;
      26028: inst = 32'h8220000;
      26029: inst = 32'h10408000;
      26030: inst = 32'hc4046b3;
      26031: inst = 32'h8220000;
      26032: inst = 32'h10408000;
      26033: inst = 32'hc4046b4;
      26034: inst = 32'h8220000;
      26035: inst = 32'h10408000;
      26036: inst = 32'hc4046b5;
      26037: inst = 32'h8220000;
      26038: inst = 32'h10408000;
      26039: inst = 32'hc4046b6;
      26040: inst = 32'h8220000;
      26041: inst = 32'h10408000;
      26042: inst = 32'hc4046b7;
      26043: inst = 32'h8220000;
      26044: inst = 32'h10408000;
      26045: inst = 32'hc4046b8;
      26046: inst = 32'h8220000;
      26047: inst = 32'h10408000;
      26048: inst = 32'hc4046b9;
      26049: inst = 32'h8220000;
      26050: inst = 32'h10408000;
      26051: inst = 32'hc4046ba;
      26052: inst = 32'h8220000;
      26053: inst = 32'h10408000;
      26054: inst = 32'hc4046bb;
      26055: inst = 32'h8220000;
      26056: inst = 32'h10408000;
      26057: inst = 32'hc4046bc;
      26058: inst = 32'h8220000;
      26059: inst = 32'h10408000;
      26060: inst = 32'hc4046bd;
      26061: inst = 32'h8220000;
      26062: inst = 32'h10408000;
      26063: inst = 32'hc4046be;
      26064: inst = 32'h8220000;
      26065: inst = 32'h10408000;
      26066: inst = 32'hc4046bf;
      26067: inst = 32'h8220000;
      26068: inst = 32'h10408000;
      26069: inst = 32'hc4046c0;
      26070: inst = 32'h8220000;
      26071: inst = 32'h10408000;
      26072: inst = 32'hc4046c1;
      26073: inst = 32'h8220000;
      26074: inst = 32'h10408000;
      26075: inst = 32'hc4046c2;
      26076: inst = 32'h8220000;
      26077: inst = 32'h10408000;
      26078: inst = 32'hc4046c3;
      26079: inst = 32'h8220000;
      26080: inst = 32'h10408000;
      26081: inst = 32'hc4046c4;
      26082: inst = 32'h8220000;
      26083: inst = 32'h10408000;
      26084: inst = 32'hc4046c5;
      26085: inst = 32'h8220000;
      26086: inst = 32'h10408000;
      26087: inst = 32'hc4046c6;
      26088: inst = 32'h8220000;
      26089: inst = 32'h10408000;
      26090: inst = 32'hc4046c7;
      26091: inst = 32'h8220000;
      26092: inst = 32'h10408000;
      26093: inst = 32'hc4046c8;
      26094: inst = 32'h8220000;
      26095: inst = 32'h10408000;
      26096: inst = 32'hc4046c9;
      26097: inst = 32'h8220000;
      26098: inst = 32'h10408000;
      26099: inst = 32'hc4046ce;
      26100: inst = 32'h8220000;
      26101: inst = 32'h10408000;
      26102: inst = 32'hc4046cf;
      26103: inst = 32'h8220000;
      26104: inst = 32'h10408000;
      26105: inst = 32'hc4046d0;
      26106: inst = 32'h8220000;
      26107: inst = 32'h10408000;
      26108: inst = 32'hc4046d1;
      26109: inst = 32'h8220000;
      26110: inst = 32'h10408000;
      26111: inst = 32'hc4046d6;
      26112: inst = 32'h8220000;
      26113: inst = 32'h10408000;
      26114: inst = 32'hc4046ec;
      26115: inst = 32'h8220000;
      26116: inst = 32'h10408000;
      26117: inst = 32'hc4046ed;
      26118: inst = 32'h8220000;
      26119: inst = 32'h10408000;
      26120: inst = 32'hc4046ee;
      26121: inst = 32'h8220000;
      26122: inst = 32'h10408000;
      26123: inst = 32'hc4046fd;
      26124: inst = 32'h8220000;
      26125: inst = 32'h10408000;
      26126: inst = 32'hc4046fe;
      26127: inst = 32'h8220000;
      26128: inst = 32'h10408000;
      26129: inst = 32'hc4046ff;
      26130: inst = 32'h8220000;
      26131: inst = 32'h10408000;
      26132: inst = 32'hc404700;
      26133: inst = 32'h8220000;
      26134: inst = 32'h10408000;
      26135: inst = 32'hc404701;
      26136: inst = 32'h8220000;
      26137: inst = 32'h10408000;
      26138: inst = 32'hc404702;
      26139: inst = 32'h8220000;
      26140: inst = 32'h10408000;
      26141: inst = 32'hc40470e;
      26142: inst = 32'h8220000;
      26143: inst = 32'h10408000;
      26144: inst = 32'hc40470f;
      26145: inst = 32'h8220000;
      26146: inst = 32'h10408000;
      26147: inst = 32'hc404710;
      26148: inst = 32'h8220000;
      26149: inst = 32'h10408000;
      26150: inst = 32'hc404711;
      26151: inst = 32'h8220000;
      26152: inst = 32'h10408000;
      26153: inst = 32'hc404712;
      26154: inst = 32'h8220000;
      26155: inst = 32'h10408000;
      26156: inst = 32'hc404713;
      26157: inst = 32'h8220000;
      26158: inst = 32'h10408000;
      26159: inst = 32'hc404714;
      26160: inst = 32'h8220000;
      26161: inst = 32'h10408000;
      26162: inst = 32'hc404715;
      26163: inst = 32'h8220000;
      26164: inst = 32'h10408000;
      26165: inst = 32'hc404716;
      26166: inst = 32'h8220000;
      26167: inst = 32'h10408000;
      26168: inst = 32'hc404717;
      26169: inst = 32'h8220000;
      26170: inst = 32'h10408000;
      26171: inst = 32'hc404718;
      26172: inst = 32'h8220000;
      26173: inst = 32'h10408000;
      26174: inst = 32'hc404719;
      26175: inst = 32'h8220000;
      26176: inst = 32'h10408000;
      26177: inst = 32'hc40471a;
      26178: inst = 32'h8220000;
      26179: inst = 32'h10408000;
      26180: inst = 32'hc40471b;
      26181: inst = 32'h8220000;
      26182: inst = 32'h10408000;
      26183: inst = 32'hc40471c;
      26184: inst = 32'h8220000;
      26185: inst = 32'h10408000;
      26186: inst = 32'hc40471d;
      26187: inst = 32'h8220000;
      26188: inst = 32'h10408000;
      26189: inst = 32'hc40471e;
      26190: inst = 32'h8220000;
      26191: inst = 32'h10408000;
      26192: inst = 32'hc40471f;
      26193: inst = 32'h8220000;
      26194: inst = 32'h10408000;
      26195: inst = 32'hc404720;
      26196: inst = 32'h8220000;
      26197: inst = 32'h10408000;
      26198: inst = 32'hc404721;
      26199: inst = 32'h8220000;
      26200: inst = 32'h10408000;
      26201: inst = 32'hc404722;
      26202: inst = 32'h8220000;
      26203: inst = 32'h10408000;
      26204: inst = 32'hc404723;
      26205: inst = 32'h8220000;
      26206: inst = 32'h10408000;
      26207: inst = 32'hc404724;
      26208: inst = 32'h8220000;
      26209: inst = 32'h10408000;
      26210: inst = 32'hc404725;
      26211: inst = 32'h8220000;
      26212: inst = 32'h10408000;
      26213: inst = 32'hc404726;
      26214: inst = 32'h8220000;
      26215: inst = 32'h10408000;
      26216: inst = 32'hc404727;
      26217: inst = 32'h8220000;
      26218: inst = 32'h10408000;
      26219: inst = 32'hc404728;
      26220: inst = 32'h8220000;
      26221: inst = 32'h10408000;
      26222: inst = 32'hc404729;
      26223: inst = 32'h8220000;
      26224: inst = 32'h10408000;
      26225: inst = 32'hc40472a;
      26226: inst = 32'h8220000;
      26227: inst = 32'h10408000;
      26228: inst = 32'hc40472f;
      26229: inst = 32'h8220000;
      26230: inst = 32'h10408000;
      26231: inst = 32'hc404736;
      26232: inst = 32'h8220000;
      26233: inst = 32'h10408000;
      26234: inst = 32'hc404737;
      26235: inst = 32'h8220000;
      26236: inst = 32'h10408000;
      26237: inst = 32'hc404738;
      26238: inst = 32'h8220000;
      26239: inst = 32'h10408000;
      26240: inst = 32'hc40474c;
      26241: inst = 32'h8220000;
      26242: inst = 32'h10408000;
      26243: inst = 32'hc40474d;
      26244: inst = 32'h8220000;
      26245: inst = 32'h10408000;
      26246: inst = 32'hc40474e;
      26247: inst = 32'h8220000;
      26248: inst = 32'h10408000;
      26249: inst = 32'hc40475d;
      26250: inst = 32'h8220000;
      26251: inst = 32'h10408000;
      26252: inst = 32'hc40475e;
      26253: inst = 32'h8220000;
      26254: inst = 32'h10408000;
      26255: inst = 32'hc40475f;
      26256: inst = 32'h8220000;
      26257: inst = 32'h10408000;
      26258: inst = 32'hc404760;
      26259: inst = 32'h8220000;
      26260: inst = 32'h10408000;
      26261: inst = 32'hc404761;
      26262: inst = 32'h8220000;
      26263: inst = 32'h10408000;
      26264: inst = 32'hc404762;
      26265: inst = 32'h8220000;
      26266: inst = 32'h10408000;
      26267: inst = 32'hc40476e;
      26268: inst = 32'h8220000;
      26269: inst = 32'h10408000;
      26270: inst = 32'hc40476f;
      26271: inst = 32'h8220000;
      26272: inst = 32'h10408000;
      26273: inst = 32'hc404770;
      26274: inst = 32'h8220000;
      26275: inst = 32'h10408000;
      26276: inst = 32'hc4047ac;
      26277: inst = 32'h8220000;
      26278: inst = 32'h10408000;
      26279: inst = 32'hc4047ad;
      26280: inst = 32'h8220000;
      26281: inst = 32'h10408000;
      26282: inst = 32'hc4047ae;
      26283: inst = 32'h8220000;
      26284: inst = 32'h10408000;
      26285: inst = 32'hc4047bd;
      26286: inst = 32'h8220000;
      26287: inst = 32'h10408000;
      26288: inst = 32'hc4047be;
      26289: inst = 32'h8220000;
      26290: inst = 32'h10408000;
      26291: inst = 32'hc4047bf;
      26292: inst = 32'h8220000;
      26293: inst = 32'h10408000;
      26294: inst = 32'hc4047c0;
      26295: inst = 32'h8220000;
      26296: inst = 32'h10408000;
      26297: inst = 32'hc4047c1;
      26298: inst = 32'h8220000;
      26299: inst = 32'h10408000;
      26300: inst = 32'hc4047c2;
      26301: inst = 32'h8220000;
      26302: inst = 32'h10408000;
      26303: inst = 32'hc4047ce;
      26304: inst = 32'h8220000;
      26305: inst = 32'h10408000;
      26306: inst = 32'hc4047cf;
      26307: inst = 32'h8220000;
      26308: inst = 32'h10408000;
      26309: inst = 32'hc4047d0;
      26310: inst = 32'h8220000;
      26311: inst = 32'h10408000;
      26312: inst = 32'hc40480c;
      26313: inst = 32'h8220000;
      26314: inst = 32'h10408000;
      26315: inst = 32'hc40480d;
      26316: inst = 32'h8220000;
      26317: inst = 32'h10408000;
      26318: inst = 32'hc40480e;
      26319: inst = 32'h8220000;
      26320: inst = 32'h10408000;
      26321: inst = 32'hc40481d;
      26322: inst = 32'h8220000;
      26323: inst = 32'h10408000;
      26324: inst = 32'hc40481e;
      26325: inst = 32'h8220000;
      26326: inst = 32'h10408000;
      26327: inst = 32'hc40481f;
      26328: inst = 32'h8220000;
      26329: inst = 32'h10408000;
      26330: inst = 32'hc404820;
      26331: inst = 32'h8220000;
      26332: inst = 32'h10408000;
      26333: inst = 32'hc404821;
      26334: inst = 32'h8220000;
      26335: inst = 32'h10408000;
      26336: inst = 32'hc404822;
      26337: inst = 32'h8220000;
      26338: inst = 32'h10408000;
      26339: inst = 32'hc40482e;
      26340: inst = 32'h8220000;
      26341: inst = 32'h10408000;
      26342: inst = 32'hc40482f;
      26343: inst = 32'h8220000;
      26344: inst = 32'h10408000;
      26345: inst = 32'hc404830;
      26346: inst = 32'h8220000;
      26347: inst = 32'h10408000;
      26348: inst = 32'hc40486c;
      26349: inst = 32'h8220000;
      26350: inst = 32'h10408000;
      26351: inst = 32'hc40486d;
      26352: inst = 32'h8220000;
      26353: inst = 32'h10408000;
      26354: inst = 32'hc40486e;
      26355: inst = 32'h8220000;
      26356: inst = 32'h10408000;
      26357: inst = 32'hc40487d;
      26358: inst = 32'h8220000;
      26359: inst = 32'h10408000;
      26360: inst = 32'hc40487e;
      26361: inst = 32'h8220000;
      26362: inst = 32'h10408000;
      26363: inst = 32'hc40487f;
      26364: inst = 32'h8220000;
      26365: inst = 32'h10408000;
      26366: inst = 32'hc404880;
      26367: inst = 32'h8220000;
      26368: inst = 32'h10408000;
      26369: inst = 32'hc404881;
      26370: inst = 32'h8220000;
      26371: inst = 32'h10408000;
      26372: inst = 32'hc404882;
      26373: inst = 32'h8220000;
      26374: inst = 32'h10408000;
      26375: inst = 32'hc40488e;
      26376: inst = 32'h8220000;
      26377: inst = 32'h10408000;
      26378: inst = 32'hc40488f;
      26379: inst = 32'h8220000;
      26380: inst = 32'h10408000;
      26381: inst = 32'hc404890;
      26382: inst = 32'h8220000;
      26383: inst = 32'h10408000;
      26384: inst = 32'hc4048cc;
      26385: inst = 32'h8220000;
      26386: inst = 32'h10408000;
      26387: inst = 32'hc4048cd;
      26388: inst = 32'h8220000;
      26389: inst = 32'h10408000;
      26390: inst = 32'hc4048ce;
      26391: inst = 32'h8220000;
      26392: inst = 32'h10408000;
      26393: inst = 32'hc4048dd;
      26394: inst = 32'h8220000;
      26395: inst = 32'h10408000;
      26396: inst = 32'hc4048de;
      26397: inst = 32'h8220000;
      26398: inst = 32'h10408000;
      26399: inst = 32'hc4048df;
      26400: inst = 32'h8220000;
      26401: inst = 32'h10408000;
      26402: inst = 32'hc4048e0;
      26403: inst = 32'h8220000;
      26404: inst = 32'h10408000;
      26405: inst = 32'hc4048e1;
      26406: inst = 32'h8220000;
      26407: inst = 32'h10408000;
      26408: inst = 32'hc4048e2;
      26409: inst = 32'h8220000;
      26410: inst = 32'h10408000;
      26411: inst = 32'hc4048ee;
      26412: inst = 32'h8220000;
      26413: inst = 32'h10408000;
      26414: inst = 32'hc4048ef;
      26415: inst = 32'h8220000;
      26416: inst = 32'h10408000;
      26417: inst = 32'hc4048f0;
      26418: inst = 32'h8220000;
      26419: inst = 32'h10408000;
      26420: inst = 32'hc40492c;
      26421: inst = 32'h8220000;
      26422: inst = 32'h10408000;
      26423: inst = 32'hc40492d;
      26424: inst = 32'h8220000;
      26425: inst = 32'h10408000;
      26426: inst = 32'hc40492e;
      26427: inst = 32'h8220000;
      26428: inst = 32'h10408000;
      26429: inst = 32'hc40493d;
      26430: inst = 32'h8220000;
      26431: inst = 32'h10408000;
      26432: inst = 32'hc40493e;
      26433: inst = 32'h8220000;
      26434: inst = 32'h10408000;
      26435: inst = 32'hc40493f;
      26436: inst = 32'h8220000;
      26437: inst = 32'h10408000;
      26438: inst = 32'hc404940;
      26439: inst = 32'h8220000;
      26440: inst = 32'h10408000;
      26441: inst = 32'hc404941;
      26442: inst = 32'h8220000;
      26443: inst = 32'h10408000;
      26444: inst = 32'hc404942;
      26445: inst = 32'h8220000;
      26446: inst = 32'h10408000;
      26447: inst = 32'hc40494e;
      26448: inst = 32'h8220000;
      26449: inst = 32'h10408000;
      26450: inst = 32'hc40494f;
      26451: inst = 32'h8220000;
      26452: inst = 32'h10408000;
      26453: inst = 32'hc404950;
      26454: inst = 32'h8220000;
      26455: inst = 32'h10408000;
      26456: inst = 32'hc404986;
      26457: inst = 32'h8220000;
      26458: inst = 32'h10408000;
      26459: inst = 32'hc404987;
      26460: inst = 32'h8220000;
      26461: inst = 32'h10408000;
      26462: inst = 32'hc404988;
      26463: inst = 32'h8220000;
      26464: inst = 32'h10408000;
      26465: inst = 32'hc404989;
      26466: inst = 32'h8220000;
      26467: inst = 32'h10408000;
      26468: inst = 32'hc40498a;
      26469: inst = 32'h8220000;
      26470: inst = 32'h10408000;
      26471: inst = 32'hc40498b;
      26472: inst = 32'h8220000;
      26473: inst = 32'h10408000;
      26474: inst = 32'hc40498c;
      26475: inst = 32'h8220000;
      26476: inst = 32'h10408000;
      26477: inst = 32'hc40498d;
      26478: inst = 32'h8220000;
      26479: inst = 32'h10408000;
      26480: inst = 32'hc40498e;
      26481: inst = 32'h8220000;
      26482: inst = 32'h10408000;
      26483: inst = 32'hc40499d;
      26484: inst = 32'h8220000;
      26485: inst = 32'h10408000;
      26486: inst = 32'hc40499e;
      26487: inst = 32'h8220000;
      26488: inst = 32'h10408000;
      26489: inst = 32'hc40499f;
      26490: inst = 32'h8220000;
      26491: inst = 32'h10408000;
      26492: inst = 32'hc4049a0;
      26493: inst = 32'h8220000;
      26494: inst = 32'h10408000;
      26495: inst = 32'hc4049a1;
      26496: inst = 32'h8220000;
      26497: inst = 32'h10408000;
      26498: inst = 32'hc4049a2;
      26499: inst = 32'h8220000;
      26500: inst = 32'h10408000;
      26501: inst = 32'hc4049ae;
      26502: inst = 32'h8220000;
      26503: inst = 32'h10408000;
      26504: inst = 32'hc4049af;
      26505: inst = 32'h8220000;
      26506: inst = 32'h10408000;
      26507: inst = 32'hc4049b0;
      26508: inst = 32'h8220000;
      26509: inst = 32'h10408000;
      26510: inst = 32'hc4049e6;
      26511: inst = 32'h8220000;
      26512: inst = 32'h10408000;
      26513: inst = 32'hc4049e7;
      26514: inst = 32'h8220000;
      26515: inst = 32'h10408000;
      26516: inst = 32'hc4049e8;
      26517: inst = 32'h8220000;
      26518: inst = 32'h10408000;
      26519: inst = 32'hc4049e9;
      26520: inst = 32'h8220000;
      26521: inst = 32'h10408000;
      26522: inst = 32'hc4049ea;
      26523: inst = 32'h8220000;
      26524: inst = 32'h10408000;
      26525: inst = 32'hc4049eb;
      26526: inst = 32'h8220000;
      26527: inst = 32'h10408000;
      26528: inst = 32'hc4049ec;
      26529: inst = 32'h8220000;
      26530: inst = 32'h10408000;
      26531: inst = 32'hc4049ed;
      26532: inst = 32'h8220000;
      26533: inst = 32'h10408000;
      26534: inst = 32'hc4049ee;
      26535: inst = 32'h8220000;
      26536: inst = 32'h10408000;
      26537: inst = 32'hc4049fd;
      26538: inst = 32'h8220000;
      26539: inst = 32'h10408000;
      26540: inst = 32'hc4049fe;
      26541: inst = 32'h8220000;
      26542: inst = 32'h10408000;
      26543: inst = 32'hc4049ff;
      26544: inst = 32'h8220000;
      26545: inst = 32'h10408000;
      26546: inst = 32'hc404a00;
      26547: inst = 32'h8220000;
      26548: inst = 32'h10408000;
      26549: inst = 32'hc404a01;
      26550: inst = 32'h8220000;
      26551: inst = 32'h10408000;
      26552: inst = 32'hc404a02;
      26553: inst = 32'h8220000;
      26554: inst = 32'h10408000;
      26555: inst = 32'hc404a0e;
      26556: inst = 32'h8220000;
      26557: inst = 32'h10408000;
      26558: inst = 32'hc404a0f;
      26559: inst = 32'h8220000;
      26560: inst = 32'h10408000;
      26561: inst = 32'hc404a10;
      26562: inst = 32'h8220000;
      26563: inst = 32'h10408000;
      26564: inst = 32'hc404a46;
      26565: inst = 32'h8220000;
      26566: inst = 32'h10408000;
      26567: inst = 32'hc404a47;
      26568: inst = 32'h8220000;
      26569: inst = 32'h10408000;
      26570: inst = 32'hc404a48;
      26571: inst = 32'h8220000;
      26572: inst = 32'h10408000;
      26573: inst = 32'hc404a49;
      26574: inst = 32'h8220000;
      26575: inst = 32'h10408000;
      26576: inst = 32'hc404a4a;
      26577: inst = 32'h8220000;
      26578: inst = 32'h10408000;
      26579: inst = 32'hc404a4b;
      26580: inst = 32'h8220000;
      26581: inst = 32'h10408000;
      26582: inst = 32'hc404a4c;
      26583: inst = 32'h8220000;
      26584: inst = 32'h10408000;
      26585: inst = 32'hc404a4d;
      26586: inst = 32'h8220000;
      26587: inst = 32'h10408000;
      26588: inst = 32'hc404a4e;
      26589: inst = 32'h8220000;
      26590: inst = 32'h10408000;
      26591: inst = 32'hc404a5d;
      26592: inst = 32'h8220000;
      26593: inst = 32'h10408000;
      26594: inst = 32'hc404a5e;
      26595: inst = 32'h8220000;
      26596: inst = 32'h10408000;
      26597: inst = 32'hc404a5f;
      26598: inst = 32'h8220000;
      26599: inst = 32'h10408000;
      26600: inst = 32'hc404a60;
      26601: inst = 32'h8220000;
      26602: inst = 32'h10408000;
      26603: inst = 32'hc404a61;
      26604: inst = 32'h8220000;
      26605: inst = 32'h10408000;
      26606: inst = 32'hc404a62;
      26607: inst = 32'h8220000;
      26608: inst = 32'h10408000;
      26609: inst = 32'hc404a6e;
      26610: inst = 32'h8220000;
      26611: inst = 32'h10408000;
      26612: inst = 32'hc404a6f;
      26613: inst = 32'h8220000;
      26614: inst = 32'h10408000;
      26615: inst = 32'hc404a70;
      26616: inst = 32'h8220000;
      26617: inst = 32'h10408000;
      26618: inst = 32'hc404abd;
      26619: inst = 32'h8220000;
      26620: inst = 32'h10408000;
      26621: inst = 32'hc404abe;
      26622: inst = 32'h8220000;
      26623: inst = 32'h10408000;
      26624: inst = 32'hc404abf;
      26625: inst = 32'h8220000;
      26626: inst = 32'h10408000;
      26627: inst = 32'hc404ac0;
      26628: inst = 32'h8220000;
      26629: inst = 32'h10408000;
      26630: inst = 32'hc404ac1;
      26631: inst = 32'h8220000;
      26632: inst = 32'h10408000;
      26633: inst = 32'hc404ac2;
      26634: inst = 32'h8220000;
      26635: inst = 32'h10408000;
      26636: inst = 32'hc404ace;
      26637: inst = 32'h8220000;
      26638: inst = 32'h10408000;
      26639: inst = 32'hc404acf;
      26640: inst = 32'h8220000;
      26641: inst = 32'h10408000;
      26642: inst = 32'hc404ad0;
      26643: inst = 32'h8220000;
      26644: inst = 32'h10408000;
      26645: inst = 32'hc404b1d;
      26646: inst = 32'h8220000;
      26647: inst = 32'h10408000;
      26648: inst = 32'hc404b1e;
      26649: inst = 32'h8220000;
      26650: inst = 32'h10408000;
      26651: inst = 32'hc404b1f;
      26652: inst = 32'h8220000;
      26653: inst = 32'h10408000;
      26654: inst = 32'hc404b20;
      26655: inst = 32'h8220000;
      26656: inst = 32'h10408000;
      26657: inst = 32'hc404b21;
      26658: inst = 32'h8220000;
      26659: inst = 32'h10408000;
      26660: inst = 32'hc404b22;
      26661: inst = 32'h8220000;
      26662: inst = 32'h10408000;
      26663: inst = 32'hc404b23;
      26664: inst = 32'h8220000;
      26665: inst = 32'h10408000;
      26666: inst = 32'hc404b24;
      26667: inst = 32'h8220000;
      26668: inst = 32'h10408000;
      26669: inst = 32'hc404b25;
      26670: inst = 32'h8220000;
      26671: inst = 32'h10408000;
      26672: inst = 32'hc404b26;
      26673: inst = 32'h8220000;
      26674: inst = 32'h10408000;
      26675: inst = 32'hc404b27;
      26676: inst = 32'h8220000;
      26677: inst = 32'h10408000;
      26678: inst = 32'hc404b28;
      26679: inst = 32'h8220000;
      26680: inst = 32'h10408000;
      26681: inst = 32'hc404b29;
      26682: inst = 32'h8220000;
      26683: inst = 32'h10408000;
      26684: inst = 32'hc404b2a;
      26685: inst = 32'h8220000;
      26686: inst = 32'h10408000;
      26687: inst = 32'hc404b2b;
      26688: inst = 32'h8220000;
      26689: inst = 32'h10408000;
      26690: inst = 32'hc404b2c;
      26691: inst = 32'h8220000;
      26692: inst = 32'h10408000;
      26693: inst = 32'hc404b2d;
      26694: inst = 32'h8220000;
      26695: inst = 32'h10408000;
      26696: inst = 32'hc404b2e;
      26697: inst = 32'h8220000;
      26698: inst = 32'h10408000;
      26699: inst = 32'hc404b2f;
      26700: inst = 32'h8220000;
      26701: inst = 32'h10408000;
      26702: inst = 32'hc404b30;
      26703: inst = 32'h8220000;
      26704: inst = 32'h10408000;
      26705: inst = 32'hc404b7d;
      26706: inst = 32'h8220000;
      26707: inst = 32'h10408000;
      26708: inst = 32'hc404b7e;
      26709: inst = 32'h8220000;
      26710: inst = 32'h10408000;
      26711: inst = 32'hc404b7f;
      26712: inst = 32'h8220000;
      26713: inst = 32'h10408000;
      26714: inst = 32'hc404b80;
      26715: inst = 32'h8220000;
      26716: inst = 32'h10408000;
      26717: inst = 32'hc404b81;
      26718: inst = 32'h8220000;
      26719: inst = 32'h10408000;
      26720: inst = 32'hc404b82;
      26721: inst = 32'h8220000;
      26722: inst = 32'h10408000;
      26723: inst = 32'hc404b83;
      26724: inst = 32'h8220000;
      26725: inst = 32'h10408000;
      26726: inst = 32'hc404b84;
      26727: inst = 32'h8220000;
      26728: inst = 32'h10408000;
      26729: inst = 32'hc404b85;
      26730: inst = 32'h8220000;
      26731: inst = 32'h10408000;
      26732: inst = 32'hc404b86;
      26733: inst = 32'h8220000;
      26734: inst = 32'h10408000;
      26735: inst = 32'hc404b87;
      26736: inst = 32'h8220000;
      26737: inst = 32'h10408000;
      26738: inst = 32'hc404b88;
      26739: inst = 32'h8220000;
      26740: inst = 32'h10408000;
      26741: inst = 32'hc404b89;
      26742: inst = 32'h8220000;
      26743: inst = 32'h10408000;
      26744: inst = 32'hc404b8a;
      26745: inst = 32'h8220000;
      26746: inst = 32'h10408000;
      26747: inst = 32'hc404b8b;
      26748: inst = 32'h8220000;
      26749: inst = 32'h10408000;
      26750: inst = 32'hc404b8c;
      26751: inst = 32'h8220000;
      26752: inst = 32'h10408000;
      26753: inst = 32'hc404b8d;
      26754: inst = 32'h8220000;
      26755: inst = 32'h10408000;
      26756: inst = 32'hc404b8e;
      26757: inst = 32'h8220000;
      26758: inst = 32'h10408000;
      26759: inst = 32'hc404b8f;
      26760: inst = 32'h8220000;
      26761: inst = 32'h10408000;
      26762: inst = 32'hc404b90;
      26763: inst = 32'h8220000;
      26764: inst = 32'h10408000;
      26765: inst = 32'hc404bdd;
      26766: inst = 32'h8220000;
      26767: inst = 32'h10408000;
      26768: inst = 32'hc404bde;
      26769: inst = 32'h8220000;
      26770: inst = 32'h10408000;
      26771: inst = 32'hc404bdf;
      26772: inst = 32'h8220000;
      26773: inst = 32'h10408000;
      26774: inst = 32'hc404be0;
      26775: inst = 32'h8220000;
      26776: inst = 32'h10408000;
      26777: inst = 32'hc404be1;
      26778: inst = 32'h8220000;
      26779: inst = 32'h10408000;
      26780: inst = 32'hc404be2;
      26781: inst = 32'h8220000;
      26782: inst = 32'h10408000;
      26783: inst = 32'hc404be3;
      26784: inst = 32'h8220000;
      26785: inst = 32'h10408000;
      26786: inst = 32'hc404be4;
      26787: inst = 32'h8220000;
      26788: inst = 32'h10408000;
      26789: inst = 32'hc404be5;
      26790: inst = 32'h8220000;
      26791: inst = 32'h10408000;
      26792: inst = 32'hc404be6;
      26793: inst = 32'h8220000;
      26794: inst = 32'h10408000;
      26795: inst = 32'hc404be7;
      26796: inst = 32'h8220000;
      26797: inst = 32'h10408000;
      26798: inst = 32'hc404be8;
      26799: inst = 32'h8220000;
      26800: inst = 32'h10408000;
      26801: inst = 32'hc404be9;
      26802: inst = 32'h8220000;
      26803: inst = 32'h10408000;
      26804: inst = 32'hc404bea;
      26805: inst = 32'h8220000;
      26806: inst = 32'h10408000;
      26807: inst = 32'hc404beb;
      26808: inst = 32'h8220000;
      26809: inst = 32'h10408000;
      26810: inst = 32'hc404bec;
      26811: inst = 32'h8220000;
      26812: inst = 32'h10408000;
      26813: inst = 32'hc404bed;
      26814: inst = 32'h8220000;
      26815: inst = 32'h10408000;
      26816: inst = 32'hc404bee;
      26817: inst = 32'h8220000;
      26818: inst = 32'h10408000;
      26819: inst = 32'hc404bef;
      26820: inst = 32'h8220000;
      26821: inst = 32'h10408000;
      26822: inst = 32'hc404bf0;
      26823: inst = 32'h8220000;
      26824: inst = 32'h10408000;
      26825: inst = 32'hc404c3d;
      26826: inst = 32'h8220000;
      26827: inst = 32'h10408000;
      26828: inst = 32'hc404c3e;
      26829: inst = 32'h8220000;
      26830: inst = 32'h10408000;
      26831: inst = 32'hc404c3f;
      26832: inst = 32'h8220000;
      26833: inst = 32'h10408000;
      26834: inst = 32'hc404c40;
      26835: inst = 32'h8220000;
      26836: inst = 32'h10408000;
      26837: inst = 32'hc404c41;
      26838: inst = 32'h8220000;
      26839: inst = 32'h10408000;
      26840: inst = 32'hc404c42;
      26841: inst = 32'h8220000;
      26842: inst = 32'h10408000;
      26843: inst = 32'hc404c9d;
      26844: inst = 32'h8220000;
      26845: inst = 32'h10408000;
      26846: inst = 32'hc404c9e;
      26847: inst = 32'h8220000;
      26848: inst = 32'h10408000;
      26849: inst = 32'hc404c9f;
      26850: inst = 32'h8220000;
      26851: inst = 32'h10408000;
      26852: inst = 32'hc404ca0;
      26853: inst = 32'h8220000;
      26854: inst = 32'h10408000;
      26855: inst = 32'hc404ca1;
      26856: inst = 32'h8220000;
      26857: inst = 32'h10408000;
      26858: inst = 32'hc404ca2;
      26859: inst = 32'h8220000;
      26860: inst = 32'h10408000;
      26861: inst = 32'hc404cfd;
      26862: inst = 32'h8220000;
      26863: inst = 32'h10408000;
      26864: inst = 32'hc404cfe;
      26865: inst = 32'h8220000;
      26866: inst = 32'h10408000;
      26867: inst = 32'hc404cff;
      26868: inst = 32'h8220000;
      26869: inst = 32'h10408000;
      26870: inst = 32'hc404d00;
      26871: inst = 32'h8220000;
      26872: inst = 32'h10408000;
      26873: inst = 32'hc404d01;
      26874: inst = 32'h8220000;
      26875: inst = 32'h10408000;
      26876: inst = 32'hc404d02;
      26877: inst = 32'h8220000;
      26878: inst = 32'h10408000;
      26879: inst = 32'hc404d25;
      26880: inst = 32'h8220000;
      26881: inst = 32'h10408000;
      26882: inst = 32'hc404d26;
      26883: inst = 32'h8220000;
      26884: inst = 32'h10408000;
      26885: inst = 32'hc404d27;
      26886: inst = 32'h8220000;
      26887: inst = 32'h10408000;
      26888: inst = 32'hc404d28;
      26889: inst = 32'h8220000;
      26890: inst = 32'h10408000;
      26891: inst = 32'hc404d29;
      26892: inst = 32'h8220000;
      26893: inst = 32'h10408000;
      26894: inst = 32'hc404d2a;
      26895: inst = 32'h8220000;
      26896: inst = 32'h10408000;
      26897: inst = 32'hc404d2b;
      26898: inst = 32'h8220000;
      26899: inst = 32'h10408000;
      26900: inst = 32'hc404d2c;
      26901: inst = 32'h8220000;
      26902: inst = 32'h10408000;
      26903: inst = 32'hc404d2d;
      26904: inst = 32'h8220000;
      26905: inst = 32'h10408000;
      26906: inst = 32'hc404d2e;
      26907: inst = 32'h8220000;
      26908: inst = 32'h10408000;
      26909: inst = 32'hc404d2f;
      26910: inst = 32'h8220000;
      26911: inst = 32'h10408000;
      26912: inst = 32'hc404d30;
      26913: inst = 32'h8220000;
      26914: inst = 32'h10408000;
      26915: inst = 32'hc404d31;
      26916: inst = 32'h8220000;
      26917: inst = 32'h10408000;
      26918: inst = 32'hc404d32;
      26919: inst = 32'h8220000;
      26920: inst = 32'h10408000;
      26921: inst = 32'hc404d33;
      26922: inst = 32'h8220000;
      26923: inst = 32'h10408000;
      26924: inst = 32'hc404d34;
      26925: inst = 32'h8220000;
      26926: inst = 32'h10408000;
      26927: inst = 32'hc404d35;
      26928: inst = 32'h8220000;
      26929: inst = 32'h10408000;
      26930: inst = 32'hc404d36;
      26931: inst = 32'h8220000;
      26932: inst = 32'h10408000;
      26933: inst = 32'hc404d37;
      26934: inst = 32'h8220000;
      26935: inst = 32'h10408000;
      26936: inst = 32'hc404d38;
      26937: inst = 32'h8220000;
      26938: inst = 32'h10408000;
      26939: inst = 32'hc404d39;
      26940: inst = 32'h8220000;
      26941: inst = 32'h10408000;
      26942: inst = 32'hc404d3a;
      26943: inst = 32'h8220000;
      26944: inst = 32'h10408000;
      26945: inst = 32'hc404d5d;
      26946: inst = 32'h8220000;
      26947: inst = 32'h10408000;
      26948: inst = 32'hc404d5e;
      26949: inst = 32'h8220000;
      26950: inst = 32'h10408000;
      26951: inst = 32'hc404d5f;
      26952: inst = 32'h8220000;
      26953: inst = 32'h10408000;
      26954: inst = 32'hc404d60;
      26955: inst = 32'h8220000;
      26956: inst = 32'h10408000;
      26957: inst = 32'hc404d61;
      26958: inst = 32'h8220000;
      26959: inst = 32'h10408000;
      26960: inst = 32'hc404d62;
      26961: inst = 32'h8220000;
      26962: inst = 32'h10408000;
      26963: inst = 32'hc404d85;
      26964: inst = 32'h8220000;
      26965: inst = 32'h10408000;
      26966: inst = 32'hc404d86;
      26967: inst = 32'h8220000;
      26968: inst = 32'h10408000;
      26969: inst = 32'hc404d87;
      26970: inst = 32'h8220000;
      26971: inst = 32'h10408000;
      26972: inst = 32'hc404d88;
      26973: inst = 32'h8220000;
      26974: inst = 32'h10408000;
      26975: inst = 32'hc404d89;
      26976: inst = 32'h8220000;
      26977: inst = 32'h10408000;
      26978: inst = 32'hc404d8a;
      26979: inst = 32'h8220000;
      26980: inst = 32'h10408000;
      26981: inst = 32'hc404d8b;
      26982: inst = 32'h8220000;
      26983: inst = 32'h10408000;
      26984: inst = 32'hc404d8c;
      26985: inst = 32'h8220000;
      26986: inst = 32'h10408000;
      26987: inst = 32'hc404d8d;
      26988: inst = 32'h8220000;
      26989: inst = 32'h10408000;
      26990: inst = 32'hc404d8e;
      26991: inst = 32'h8220000;
      26992: inst = 32'h10408000;
      26993: inst = 32'hc404d8f;
      26994: inst = 32'h8220000;
      26995: inst = 32'h10408000;
      26996: inst = 32'hc404d90;
      26997: inst = 32'h8220000;
      26998: inst = 32'h10408000;
      26999: inst = 32'hc404d91;
      27000: inst = 32'h8220000;
      27001: inst = 32'h10408000;
      27002: inst = 32'hc404d92;
      27003: inst = 32'h8220000;
      27004: inst = 32'h10408000;
      27005: inst = 32'hc404d93;
      27006: inst = 32'h8220000;
      27007: inst = 32'h10408000;
      27008: inst = 32'hc404d94;
      27009: inst = 32'h8220000;
      27010: inst = 32'h10408000;
      27011: inst = 32'hc404d95;
      27012: inst = 32'h8220000;
      27013: inst = 32'h10408000;
      27014: inst = 32'hc404d96;
      27015: inst = 32'h8220000;
      27016: inst = 32'h10408000;
      27017: inst = 32'hc404d97;
      27018: inst = 32'h8220000;
      27019: inst = 32'h10408000;
      27020: inst = 32'hc404d98;
      27021: inst = 32'h8220000;
      27022: inst = 32'h10408000;
      27023: inst = 32'hc404d99;
      27024: inst = 32'h8220000;
      27025: inst = 32'h10408000;
      27026: inst = 32'hc404d9a;
      27027: inst = 32'h8220000;
      27028: inst = 32'h10408000;
      27029: inst = 32'hc404dbd;
      27030: inst = 32'h8220000;
      27031: inst = 32'h10408000;
      27032: inst = 32'hc404dbe;
      27033: inst = 32'h8220000;
      27034: inst = 32'h10408000;
      27035: inst = 32'hc404dbf;
      27036: inst = 32'h8220000;
      27037: inst = 32'h10408000;
      27038: inst = 32'hc404dc0;
      27039: inst = 32'h8220000;
      27040: inst = 32'h10408000;
      27041: inst = 32'hc404dc1;
      27042: inst = 32'h8220000;
      27043: inst = 32'h10408000;
      27044: inst = 32'hc404dc2;
      27045: inst = 32'h8220000;
      27046: inst = 32'h10408000;
      27047: inst = 32'hc404de5;
      27048: inst = 32'h8220000;
      27049: inst = 32'h10408000;
      27050: inst = 32'hc404de6;
      27051: inst = 32'h8220000;
      27052: inst = 32'h10408000;
      27053: inst = 32'hc404de7;
      27054: inst = 32'h8220000;
      27055: inst = 32'h10408000;
      27056: inst = 32'hc404de8;
      27057: inst = 32'h8220000;
      27058: inst = 32'h10408000;
      27059: inst = 32'hc404de9;
      27060: inst = 32'h8220000;
      27061: inst = 32'h10408000;
      27062: inst = 32'hc404dea;
      27063: inst = 32'h8220000;
      27064: inst = 32'h10408000;
      27065: inst = 32'hc404deb;
      27066: inst = 32'h8220000;
      27067: inst = 32'h10408000;
      27068: inst = 32'hc404dec;
      27069: inst = 32'h8220000;
      27070: inst = 32'h10408000;
      27071: inst = 32'hc404ded;
      27072: inst = 32'h8220000;
      27073: inst = 32'h10408000;
      27074: inst = 32'hc404dee;
      27075: inst = 32'h8220000;
      27076: inst = 32'h10408000;
      27077: inst = 32'hc404def;
      27078: inst = 32'h8220000;
      27079: inst = 32'h10408000;
      27080: inst = 32'hc404df0;
      27081: inst = 32'h8220000;
      27082: inst = 32'h10408000;
      27083: inst = 32'hc404df1;
      27084: inst = 32'h8220000;
      27085: inst = 32'h10408000;
      27086: inst = 32'hc404df2;
      27087: inst = 32'h8220000;
      27088: inst = 32'h10408000;
      27089: inst = 32'hc404df3;
      27090: inst = 32'h8220000;
      27091: inst = 32'h10408000;
      27092: inst = 32'hc404df4;
      27093: inst = 32'h8220000;
      27094: inst = 32'h10408000;
      27095: inst = 32'hc404df5;
      27096: inst = 32'h8220000;
      27097: inst = 32'h10408000;
      27098: inst = 32'hc404df6;
      27099: inst = 32'h8220000;
      27100: inst = 32'h10408000;
      27101: inst = 32'hc404df7;
      27102: inst = 32'h8220000;
      27103: inst = 32'h10408000;
      27104: inst = 32'hc404df8;
      27105: inst = 32'h8220000;
      27106: inst = 32'h10408000;
      27107: inst = 32'hc404df9;
      27108: inst = 32'h8220000;
      27109: inst = 32'h10408000;
      27110: inst = 32'hc404dfa;
      27111: inst = 32'h8220000;
      27112: inst = 32'h10408000;
      27113: inst = 32'hc404e1d;
      27114: inst = 32'h8220000;
      27115: inst = 32'h10408000;
      27116: inst = 32'hc404e1e;
      27117: inst = 32'h8220000;
      27118: inst = 32'h10408000;
      27119: inst = 32'hc404e1f;
      27120: inst = 32'h8220000;
      27121: inst = 32'h10408000;
      27122: inst = 32'hc404e20;
      27123: inst = 32'h8220000;
      27124: inst = 32'h10408000;
      27125: inst = 32'hc404e21;
      27126: inst = 32'h8220000;
      27127: inst = 32'h10408000;
      27128: inst = 32'hc404e22;
      27129: inst = 32'h8220000;
      27130: inst = 32'h10408000;
      27131: inst = 32'hc404e58;
      27132: inst = 32'h8220000;
      27133: inst = 32'h10408000;
      27134: inst = 32'hc404e59;
      27135: inst = 32'h8220000;
      27136: inst = 32'h10408000;
      27137: inst = 32'hc404e5a;
      27138: inst = 32'h8220000;
      27139: inst = 32'h10408000;
      27140: inst = 32'hc404e7d;
      27141: inst = 32'h8220000;
      27142: inst = 32'h10408000;
      27143: inst = 32'hc404e7e;
      27144: inst = 32'h8220000;
      27145: inst = 32'h10408000;
      27146: inst = 32'hc404e7f;
      27147: inst = 32'h8220000;
      27148: inst = 32'h10408000;
      27149: inst = 32'hc404e80;
      27150: inst = 32'h8220000;
      27151: inst = 32'h10408000;
      27152: inst = 32'hc404e81;
      27153: inst = 32'h8220000;
      27154: inst = 32'h10408000;
      27155: inst = 32'hc404e82;
      27156: inst = 32'h8220000;
      27157: inst = 32'h10408000;
      27158: inst = 32'hc404eb8;
      27159: inst = 32'h8220000;
      27160: inst = 32'h10408000;
      27161: inst = 32'hc404eb9;
      27162: inst = 32'h8220000;
      27163: inst = 32'h10408000;
      27164: inst = 32'hc404eba;
      27165: inst = 32'h8220000;
      27166: inst = 32'h10408000;
      27167: inst = 32'hc404edd;
      27168: inst = 32'h8220000;
      27169: inst = 32'h10408000;
      27170: inst = 32'hc404ede;
      27171: inst = 32'h8220000;
      27172: inst = 32'h10408000;
      27173: inst = 32'hc404edf;
      27174: inst = 32'h8220000;
      27175: inst = 32'h10408000;
      27176: inst = 32'hc404ee0;
      27177: inst = 32'h8220000;
      27178: inst = 32'h10408000;
      27179: inst = 32'hc404ee1;
      27180: inst = 32'h8220000;
      27181: inst = 32'h10408000;
      27182: inst = 32'hc404ee2;
      27183: inst = 32'h8220000;
      27184: inst = 32'h10408000;
      27185: inst = 32'hc404f18;
      27186: inst = 32'h8220000;
      27187: inst = 32'h10408000;
      27188: inst = 32'hc404f19;
      27189: inst = 32'h8220000;
      27190: inst = 32'h10408000;
      27191: inst = 32'hc404f1a;
      27192: inst = 32'h8220000;
      27193: inst = 32'h10408000;
      27194: inst = 32'hc404f3d;
      27195: inst = 32'h8220000;
      27196: inst = 32'h10408000;
      27197: inst = 32'hc404f3e;
      27198: inst = 32'h8220000;
      27199: inst = 32'h10408000;
      27200: inst = 32'hc404f3f;
      27201: inst = 32'h8220000;
      27202: inst = 32'h10408000;
      27203: inst = 32'hc404f40;
      27204: inst = 32'h8220000;
      27205: inst = 32'h10408000;
      27206: inst = 32'hc404f41;
      27207: inst = 32'h8220000;
      27208: inst = 32'h10408000;
      27209: inst = 32'hc404f42;
      27210: inst = 32'h8220000;
      27211: inst = 32'h10408000;
      27212: inst = 32'hc404f78;
      27213: inst = 32'h8220000;
      27214: inst = 32'h10408000;
      27215: inst = 32'hc404f79;
      27216: inst = 32'h8220000;
      27217: inst = 32'h10408000;
      27218: inst = 32'hc404f7a;
      27219: inst = 32'h8220000;
      27220: inst = 32'h10408000;
      27221: inst = 32'hc404f9d;
      27222: inst = 32'h8220000;
      27223: inst = 32'h10408000;
      27224: inst = 32'hc404f9e;
      27225: inst = 32'h8220000;
      27226: inst = 32'h10408000;
      27227: inst = 32'hc404f9f;
      27228: inst = 32'h8220000;
      27229: inst = 32'h10408000;
      27230: inst = 32'hc404fa0;
      27231: inst = 32'h8220000;
      27232: inst = 32'h10408000;
      27233: inst = 32'hc404fa1;
      27234: inst = 32'h8220000;
      27235: inst = 32'h10408000;
      27236: inst = 32'hc404fa2;
      27237: inst = 32'h8220000;
      27238: inst = 32'h10408000;
      27239: inst = 32'hc404fd8;
      27240: inst = 32'h8220000;
      27241: inst = 32'h10408000;
      27242: inst = 32'hc404fd9;
      27243: inst = 32'h8220000;
      27244: inst = 32'h10408000;
      27245: inst = 32'hc404fda;
      27246: inst = 32'h8220000;
      27247: inst = 32'h10408000;
      27248: inst = 32'hc404ffd;
      27249: inst = 32'h8220000;
      27250: inst = 32'h10408000;
      27251: inst = 32'hc404ffe;
      27252: inst = 32'h8220000;
      27253: inst = 32'h10408000;
      27254: inst = 32'hc404fff;
      27255: inst = 32'h8220000;
      27256: inst = 32'h10408000;
      27257: inst = 32'hc405000;
      27258: inst = 32'h8220000;
      27259: inst = 32'h10408000;
      27260: inst = 32'hc405001;
      27261: inst = 32'h8220000;
      27262: inst = 32'h10408000;
      27263: inst = 32'hc405002;
      27264: inst = 32'h8220000;
      27265: inst = 32'h10408000;
      27266: inst = 32'hc405038;
      27267: inst = 32'h8220000;
      27268: inst = 32'h10408000;
      27269: inst = 32'hc405039;
      27270: inst = 32'h8220000;
      27271: inst = 32'h10408000;
      27272: inst = 32'hc40503a;
      27273: inst = 32'h8220000;
      27274: inst = 32'h10408000;
      27275: inst = 32'hc40505d;
      27276: inst = 32'h8220000;
      27277: inst = 32'h10408000;
      27278: inst = 32'hc40505e;
      27279: inst = 32'h8220000;
      27280: inst = 32'h10408000;
      27281: inst = 32'hc40505f;
      27282: inst = 32'h8220000;
      27283: inst = 32'h10408000;
      27284: inst = 32'hc405060;
      27285: inst = 32'h8220000;
      27286: inst = 32'h10408000;
      27287: inst = 32'hc405061;
      27288: inst = 32'h8220000;
      27289: inst = 32'h10408000;
      27290: inst = 32'hc405062;
      27291: inst = 32'h8220000;
      27292: inst = 32'h10408000;
      27293: inst = 32'hc405098;
      27294: inst = 32'h8220000;
      27295: inst = 32'h10408000;
      27296: inst = 32'hc405099;
      27297: inst = 32'h8220000;
      27298: inst = 32'h10408000;
      27299: inst = 32'hc40509a;
      27300: inst = 32'h8220000;
      27301: inst = 32'h10408000;
      27302: inst = 32'hc40509b;
      27303: inst = 32'h8220000;
      27304: inst = 32'h10408000;
      27305: inst = 32'hc40509c;
      27306: inst = 32'h8220000;
      27307: inst = 32'h10408000;
      27308: inst = 32'hc40509d;
      27309: inst = 32'h8220000;
      27310: inst = 32'h10408000;
      27311: inst = 32'hc40509e;
      27312: inst = 32'h8220000;
      27313: inst = 32'h10408000;
      27314: inst = 32'hc40509f;
      27315: inst = 32'h8220000;
      27316: inst = 32'h10408000;
      27317: inst = 32'hc4050a0;
      27318: inst = 32'h8220000;
      27319: inst = 32'h10408000;
      27320: inst = 32'hc4050a1;
      27321: inst = 32'h8220000;
      27322: inst = 32'h10408000;
      27323: inst = 32'hc4050a2;
      27324: inst = 32'h8220000;
      27325: inst = 32'h10408000;
      27326: inst = 32'hc4050a3;
      27327: inst = 32'h8220000;
      27328: inst = 32'h10408000;
      27329: inst = 32'hc4050a4;
      27330: inst = 32'h8220000;
      27331: inst = 32'h10408000;
      27332: inst = 32'hc4050a5;
      27333: inst = 32'h8220000;
      27334: inst = 32'h10408000;
      27335: inst = 32'hc4050a6;
      27336: inst = 32'h8220000;
      27337: inst = 32'h10408000;
      27338: inst = 32'hc4050a7;
      27339: inst = 32'h8220000;
      27340: inst = 32'h10408000;
      27341: inst = 32'hc4050a8;
      27342: inst = 32'h8220000;
      27343: inst = 32'h10408000;
      27344: inst = 32'hc4050a9;
      27345: inst = 32'h8220000;
      27346: inst = 32'h10408000;
      27347: inst = 32'hc4050aa;
      27348: inst = 32'h8220000;
      27349: inst = 32'h10408000;
      27350: inst = 32'hc4050ab;
      27351: inst = 32'h8220000;
      27352: inst = 32'h10408000;
      27353: inst = 32'hc4050ac;
      27354: inst = 32'h8220000;
      27355: inst = 32'h10408000;
      27356: inst = 32'hc4050ad;
      27357: inst = 32'h8220000;
      27358: inst = 32'h10408000;
      27359: inst = 32'hc4050ae;
      27360: inst = 32'h8220000;
      27361: inst = 32'h10408000;
      27362: inst = 32'hc4050af;
      27363: inst = 32'h8220000;
      27364: inst = 32'h10408000;
      27365: inst = 32'hc4050b0;
      27366: inst = 32'h8220000;
      27367: inst = 32'h10408000;
      27368: inst = 32'hc4050b1;
      27369: inst = 32'h8220000;
      27370: inst = 32'h10408000;
      27371: inst = 32'hc4050b2;
      27372: inst = 32'h8220000;
      27373: inst = 32'h10408000;
      27374: inst = 32'hc4050b3;
      27375: inst = 32'h8220000;
      27376: inst = 32'h10408000;
      27377: inst = 32'hc4050b4;
      27378: inst = 32'h8220000;
      27379: inst = 32'h10408000;
      27380: inst = 32'hc4050b5;
      27381: inst = 32'h8220000;
      27382: inst = 32'h10408000;
      27383: inst = 32'hc4050b6;
      27384: inst = 32'h8220000;
      27385: inst = 32'h10408000;
      27386: inst = 32'hc4050b7;
      27387: inst = 32'h8220000;
      27388: inst = 32'h10408000;
      27389: inst = 32'hc4050b8;
      27390: inst = 32'h8220000;
      27391: inst = 32'h10408000;
      27392: inst = 32'hc4050b9;
      27393: inst = 32'h8220000;
      27394: inst = 32'h10408000;
      27395: inst = 32'hc4050ba;
      27396: inst = 32'h8220000;
      27397: inst = 32'h10408000;
      27398: inst = 32'hc4050bb;
      27399: inst = 32'h8220000;
      27400: inst = 32'h10408000;
      27401: inst = 32'hc4050bc;
      27402: inst = 32'h8220000;
      27403: inst = 32'h10408000;
      27404: inst = 32'hc4050bd;
      27405: inst = 32'h8220000;
      27406: inst = 32'h10408000;
      27407: inst = 32'hc4050be;
      27408: inst = 32'h8220000;
      27409: inst = 32'h10408000;
      27410: inst = 32'hc4050bf;
      27411: inst = 32'h8220000;
      27412: inst = 32'h10408000;
      27413: inst = 32'hc4050c0;
      27414: inst = 32'h8220000;
      27415: inst = 32'h10408000;
      27416: inst = 32'hc4050c1;
      27417: inst = 32'h8220000;
      27418: inst = 32'h10408000;
      27419: inst = 32'hc4050c2;
      27420: inst = 32'h8220000;
      27421: inst = 32'h10408000;
      27422: inst = 32'hc4050f8;
      27423: inst = 32'h8220000;
      27424: inst = 32'h10408000;
      27425: inst = 32'hc4050f9;
      27426: inst = 32'h8220000;
      27427: inst = 32'h10408000;
      27428: inst = 32'hc4050fa;
      27429: inst = 32'h8220000;
      27430: inst = 32'h10408000;
      27431: inst = 32'hc4050fb;
      27432: inst = 32'h8220000;
      27433: inst = 32'h10408000;
      27434: inst = 32'hc4050fc;
      27435: inst = 32'h8220000;
      27436: inst = 32'h10408000;
      27437: inst = 32'hc4050fd;
      27438: inst = 32'h8220000;
      27439: inst = 32'h10408000;
      27440: inst = 32'hc4050fe;
      27441: inst = 32'h8220000;
      27442: inst = 32'h10408000;
      27443: inst = 32'hc4050ff;
      27444: inst = 32'h8220000;
      27445: inst = 32'h10408000;
      27446: inst = 32'hc405100;
      27447: inst = 32'h8220000;
      27448: inst = 32'h10408000;
      27449: inst = 32'hc405101;
      27450: inst = 32'h8220000;
      27451: inst = 32'h10408000;
      27452: inst = 32'hc405102;
      27453: inst = 32'h8220000;
      27454: inst = 32'h10408000;
      27455: inst = 32'hc405103;
      27456: inst = 32'h8220000;
      27457: inst = 32'h10408000;
      27458: inst = 32'hc405104;
      27459: inst = 32'h8220000;
      27460: inst = 32'h10408000;
      27461: inst = 32'hc405105;
      27462: inst = 32'h8220000;
      27463: inst = 32'h10408000;
      27464: inst = 32'hc405106;
      27465: inst = 32'h8220000;
      27466: inst = 32'h10408000;
      27467: inst = 32'hc405107;
      27468: inst = 32'h8220000;
      27469: inst = 32'h10408000;
      27470: inst = 32'hc405108;
      27471: inst = 32'h8220000;
      27472: inst = 32'h10408000;
      27473: inst = 32'hc405109;
      27474: inst = 32'h8220000;
      27475: inst = 32'h10408000;
      27476: inst = 32'hc40510a;
      27477: inst = 32'h8220000;
      27478: inst = 32'h10408000;
      27479: inst = 32'hc40510b;
      27480: inst = 32'h8220000;
      27481: inst = 32'h10408000;
      27482: inst = 32'hc40510c;
      27483: inst = 32'h8220000;
      27484: inst = 32'h10408000;
      27485: inst = 32'hc40510d;
      27486: inst = 32'h8220000;
      27487: inst = 32'h10408000;
      27488: inst = 32'hc40510e;
      27489: inst = 32'h8220000;
      27490: inst = 32'h10408000;
      27491: inst = 32'hc40510f;
      27492: inst = 32'h8220000;
      27493: inst = 32'h10408000;
      27494: inst = 32'hc405110;
      27495: inst = 32'h8220000;
      27496: inst = 32'h10408000;
      27497: inst = 32'hc405111;
      27498: inst = 32'h8220000;
      27499: inst = 32'h10408000;
      27500: inst = 32'hc405112;
      27501: inst = 32'h8220000;
      27502: inst = 32'h10408000;
      27503: inst = 32'hc405113;
      27504: inst = 32'h8220000;
      27505: inst = 32'h10408000;
      27506: inst = 32'hc405114;
      27507: inst = 32'h8220000;
      27508: inst = 32'h10408000;
      27509: inst = 32'hc405115;
      27510: inst = 32'h8220000;
      27511: inst = 32'h10408000;
      27512: inst = 32'hc405116;
      27513: inst = 32'h8220000;
      27514: inst = 32'h10408000;
      27515: inst = 32'hc405117;
      27516: inst = 32'h8220000;
      27517: inst = 32'h10408000;
      27518: inst = 32'hc405118;
      27519: inst = 32'h8220000;
      27520: inst = 32'h10408000;
      27521: inst = 32'hc405119;
      27522: inst = 32'h8220000;
      27523: inst = 32'h10408000;
      27524: inst = 32'hc40511a;
      27525: inst = 32'h8220000;
      27526: inst = 32'h10408000;
      27527: inst = 32'hc40511b;
      27528: inst = 32'h8220000;
      27529: inst = 32'h10408000;
      27530: inst = 32'hc40511c;
      27531: inst = 32'h8220000;
      27532: inst = 32'h10408000;
      27533: inst = 32'hc40511d;
      27534: inst = 32'h8220000;
      27535: inst = 32'h10408000;
      27536: inst = 32'hc40511e;
      27537: inst = 32'h8220000;
      27538: inst = 32'h10408000;
      27539: inst = 32'hc40511f;
      27540: inst = 32'h8220000;
      27541: inst = 32'h10408000;
      27542: inst = 32'hc405120;
      27543: inst = 32'h8220000;
      27544: inst = 32'h10408000;
      27545: inst = 32'hc405121;
      27546: inst = 32'h8220000;
      27547: inst = 32'h10408000;
      27548: inst = 32'hc405122;
      27549: inst = 32'h8220000;
      27550: inst = 32'h10408000;
      27551: inst = 32'hc405136;
      27552: inst = 32'h8220000;
      27553: inst = 32'h10408000;
      27554: inst = 32'hc405137;
      27555: inst = 32'h8220000;
      27556: inst = 32'h10408000;
      27557: inst = 32'hc405138;
      27558: inst = 32'h8220000;
      27559: inst = 32'h10408000;
      27560: inst = 32'hc405158;
      27561: inst = 32'h8220000;
      27562: inst = 32'h10408000;
      27563: inst = 32'hc405159;
      27564: inst = 32'h8220000;
      27565: inst = 32'h10408000;
      27566: inst = 32'hc40515a;
      27567: inst = 32'h8220000;
      27568: inst = 32'h10408000;
      27569: inst = 32'hc40515b;
      27570: inst = 32'h8220000;
      27571: inst = 32'h10408000;
      27572: inst = 32'hc40515c;
      27573: inst = 32'h8220000;
      27574: inst = 32'h10408000;
      27575: inst = 32'hc40515d;
      27576: inst = 32'h8220000;
      27577: inst = 32'h10408000;
      27578: inst = 32'hc40515e;
      27579: inst = 32'h8220000;
      27580: inst = 32'h10408000;
      27581: inst = 32'hc40515f;
      27582: inst = 32'h8220000;
      27583: inst = 32'h10408000;
      27584: inst = 32'hc405160;
      27585: inst = 32'h8220000;
      27586: inst = 32'h10408000;
      27587: inst = 32'hc405161;
      27588: inst = 32'h8220000;
      27589: inst = 32'h10408000;
      27590: inst = 32'hc405162;
      27591: inst = 32'h8220000;
      27592: inst = 32'h10408000;
      27593: inst = 32'hc405163;
      27594: inst = 32'h8220000;
      27595: inst = 32'h10408000;
      27596: inst = 32'hc405164;
      27597: inst = 32'h8220000;
      27598: inst = 32'h10408000;
      27599: inst = 32'hc405165;
      27600: inst = 32'h8220000;
      27601: inst = 32'h10408000;
      27602: inst = 32'hc405166;
      27603: inst = 32'h8220000;
      27604: inst = 32'h10408000;
      27605: inst = 32'hc405167;
      27606: inst = 32'h8220000;
      27607: inst = 32'h10408000;
      27608: inst = 32'hc405168;
      27609: inst = 32'h8220000;
      27610: inst = 32'h10408000;
      27611: inst = 32'hc405169;
      27612: inst = 32'h8220000;
      27613: inst = 32'h10408000;
      27614: inst = 32'hc40516a;
      27615: inst = 32'h8220000;
      27616: inst = 32'h10408000;
      27617: inst = 32'hc40516b;
      27618: inst = 32'h8220000;
      27619: inst = 32'h10408000;
      27620: inst = 32'hc40516c;
      27621: inst = 32'h8220000;
      27622: inst = 32'h10408000;
      27623: inst = 32'hc40516d;
      27624: inst = 32'h8220000;
      27625: inst = 32'h10408000;
      27626: inst = 32'hc40516e;
      27627: inst = 32'h8220000;
      27628: inst = 32'h10408000;
      27629: inst = 32'hc40516f;
      27630: inst = 32'h8220000;
      27631: inst = 32'h10408000;
      27632: inst = 32'hc405170;
      27633: inst = 32'h8220000;
      27634: inst = 32'h10408000;
      27635: inst = 32'hc405171;
      27636: inst = 32'h8220000;
      27637: inst = 32'h10408000;
      27638: inst = 32'hc405172;
      27639: inst = 32'h8220000;
      27640: inst = 32'h10408000;
      27641: inst = 32'hc405173;
      27642: inst = 32'h8220000;
      27643: inst = 32'h10408000;
      27644: inst = 32'hc405174;
      27645: inst = 32'h8220000;
      27646: inst = 32'h10408000;
      27647: inst = 32'hc405175;
      27648: inst = 32'h8220000;
      27649: inst = 32'h10408000;
      27650: inst = 32'hc405176;
      27651: inst = 32'h8220000;
      27652: inst = 32'h10408000;
      27653: inst = 32'hc405177;
      27654: inst = 32'h8220000;
      27655: inst = 32'h10408000;
      27656: inst = 32'hc405178;
      27657: inst = 32'h8220000;
      27658: inst = 32'h10408000;
      27659: inst = 32'hc405179;
      27660: inst = 32'h8220000;
      27661: inst = 32'h10408000;
      27662: inst = 32'hc40517a;
      27663: inst = 32'h8220000;
      27664: inst = 32'h10408000;
      27665: inst = 32'hc40517b;
      27666: inst = 32'h8220000;
      27667: inst = 32'h10408000;
      27668: inst = 32'hc40517c;
      27669: inst = 32'h8220000;
      27670: inst = 32'h10408000;
      27671: inst = 32'hc40517d;
      27672: inst = 32'h8220000;
      27673: inst = 32'h10408000;
      27674: inst = 32'hc40517e;
      27675: inst = 32'h8220000;
      27676: inst = 32'h10408000;
      27677: inst = 32'hc40517f;
      27678: inst = 32'h8220000;
      27679: inst = 32'h10408000;
      27680: inst = 32'hc405180;
      27681: inst = 32'h8220000;
      27682: inst = 32'h10408000;
      27683: inst = 32'hc405181;
      27684: inst = 32'h8220000;
      27685: inst = 32'h10408000;
      27686: inst = 32'hc405182;
      27687: inst = 32'h8220000;
      27688: inst = 32'h10408000;
      27689: inst = 32'hc405196;
      27690: inst = 32'h8220000;
      27691: inst = 32'h10408000;
      27692: inst = 32'hc405197;
      27693: inst = 32'h8220000;
      27694: inst = 32'h10408000;
      27695: inst = 32'hc405198;
      27696: inst = 32'h8220000;
      27697: inst = 32'h10408000;
      27698: inst = 32'hc4051dd;
      27699: inst = 32'h8220000;
      27700: inst = 32'h10408000;
      27701: inst = 32'hc4051de;
      27702: inst = 32'h8220000;
      27703: inst = 32'h10408000;
      27704: inst = 32'hc4051df;
      27705: inst = 32'h8220000;
      27706: inst = 32'h10408000;
      27707: inst = 32'hc4051e0;
      27708: inst = 32'h8220000;
      27709: inst = 32'h10408000;
      27710: inst = 32'hc4051e1;
      27711: inst = 32'h8220000;
      27712: inst = 32'h10408000;
      27713: inst = 32'hc4051e2;
      27714: inst = 32'h8220000;
      27715: inst = 32'h10408000;
      27716: inst = 32'hc4051f6;
      27717: inst = 32'h8220000;
      27718: inst = 32'h10408000;
      27719: inst = 32'hc4051f7;
      27720: inst = 32'h8220000;
      27721: inst = 32'h10408000;
      27722: inst = 32'hc4051f8;
      27723: inst = 32'h8220000;
      27724: inst = 32'h10408000;
      27725: inst = 32'hc40523d;
      27726: inst = 32'h8220000;
      27727: inst = 32'h10408000;
      27728: inst = 32'hc40523e;
      27729: inst = 32'h8220000;
      27730: inst = 32'h10408000;
      27731: inst = 32'hc40523f;
      27732: inst = 32'h8220000;
      27733: inst = 32'h10408000;
      27734: inst = 32'hc405240;
      27735: inst = 32'h8220000;
      27736: inst = 32'h10408000;
      27737: inst = 32'hc405241;
      27738: inst = 32'h8220000;
      27739: inst = 32'h10408000;
      27740: inst = 32'hc405242;
      27741: inst = 32'h8220000;
      27742: inst = 32'h10408000;
      27743: inst = 32'hc405256;
      27744: inst = 32'h8220000;
      27745: inst = 32'h10408000;
      27746: inst = 32'hc405257;
      27747: inst = 32'h8220000;
      27748: inst = 32'h10408000;
      27749: inst = 32'hc405258;
      27750: inst = 32'h8220000;
      27751: inst = 32'h10408000;
      27752: inst = 32'hc40529d;
      27753: inst = 32'h8220000;
      27754: inst = 32'h10408000;
      27755: inst = 32'hc40529e;
      27756: inst = 32'h8220000;
      27757: inst = 32'h10408000;
      27758: inst = 32'hc40529f;
      27759: inst = 32'h8220000;
      27760: inst = 32'h10408000;
      27761: inst = 32'hc4052a0;
      27762: inst = 32'h8220000;
      27763: inst = 32'h10408000;
      27764: inst = 32'hc4052a1;
      27765: inst = 32'h8220000;
      27766: inst = 32'h10408000;
      27767: inst = 32'hc4052a2;
      27768: inst = 32'h8220000;
      27769: inst = 32'h10408000;
      27770: inst = 32'hc4052b6;
      27771: inst = 32'h8220000;
      27772: inst = 32'h10408000;
      27773: inst = 32'hc4052b7;
      27774: inst = 32'h8220000;
      27775: inst = 32'h10408000;
      27776: inst = 32'hc4052b8;
      27777: inst = 32'h8220000;
      27778: inst = 32'h10408000;
      27779: inst = 32'hc4052fd;
      27780: inst = 32'h8220000;
      27781: inst = 32'h10408000;
      27782: inst = 32'hc4052fe;
      27783: inst = 32'h8220000;
      27784: inst = 32'h10408000;
      27785: inst = 32'hc4052ff;
      27786: inst = 32'h8220000;
      27787: inst = 32'h10408000;
      27788: inst = 32'hc405300;
      27789: inst = 32'h8220000;
      27790: inst = 32'h10408000;
      27791: inst = 32'hc405301;
      27792: inst = 32'h8220000;
      27793: inst = 32'h10408000;
      27794: inst = 32'hc405302;
      27795: inst = 32'h8220000;
      27796: inst = 32'h10408000;
      27797: inst = 32'hc405316;
      27798: inst = 32'h8220000;
      27799: inst = 32'h10408000;
      27800: inst = 32'hc405317;
      27801: inst = 32'h8220000;
      27802: inst = 32'h10408000;
      27803: inst = 32'hc405318;
      27804: inst = 32'h8220000;
      27805: inst = 32'h10408000;
      27806: inst = 32'hc40535d;
      27807: inst = 32'h8220000;
      27808: inst = 32'h10408000;
      27809: inst = 32'hc40535e;
      27810: inst = 32'h8220000;
      27811: inst = 32'h10408000;
      27812: inst = 32'hc40535f;
      27813: inst = 32'h8220000;
      27814: inst = 32'h10408000;
      27815: inst = 32'hc405360;
      27816: inst = 32'h8220000;
      27817: inst = 32'h10408000;
      27818: inst = 32'hc405361;
      27819: inst = 32'h8220000;
      27820: inst = 32'h10408000;
      27821: inst = 32'hc405362;
      27822: inst = 32'h8220000;
      27823: inst = 32'h10408000;
      27824: inst = 32'hc405376;
      27825: inst = 32'h8220000;
      27826: inst = 32'h10408000;
      27827: inst = 32'hc405377;
      27828: inst = 32'h8220000;
      27829: inst = 32'h10408000;
      27830: inst = 32'hc405378;
      27831: inst = 32'h8220000;
      27832: inst = 32'h10408000;
      27833: inst = 32'hc4053bd;
      27834: inst = 32'h8220000;
      27835: inst = 32'h10408000;
      27836: inst = 32'hc4053be;
      27837: inst = 32'h8220000;
      27838: inst = 32'h10408000;
      27839: inst = 32'hc4053bf;
      27840: inst = 32'h8220000;
      27841: inst = 32'h10408000;
      27842: inst = 32'hc4053c0;
      27843: inst = 32'h8220000;
      27844: inst = 32'h10408000;
      27845: inst = 32'hc4053c1;
      27846: inst = 32'h8220000;
      27847: inst = 32'h10408000;
      27848: inst = 32'hc4053c2;
      27849: inst = 32'h8220000;
      27850: inst = 32'h10408000;
      27851: inst = 32'hc4053d6;
      27852: inst = 32'h8220000;
      27853: inst = 32'h10408000;
      27854: inst = 32'hc4053d7;
      27855: inst = 32'h8220000;
      27856: inst = 32'h10408000;
      27857: inst = 32'hc4053d8;
      27858: inst = 32'h8220000;
      27859: inst = 32'h10408000;
      27860: inst = 32'hc40541d;
      27861: inst = 32'h8220000;
      27862: inst = 32'h10408000;
      27863: inst = 32'hc40541e;
      27864: inst = 32'h8220000;
      27865: inst = 32'h10408000;
      27866: inst = 32'hc40541f;
      27867: inst = 32'h8220000;
      27868: inst = 32'h10408000;
      27869: inst = 32'hc405420;
      27870: inst = 32'h8220000;
      27871: inst = 32'h10408000;
      27872: inst = 32'hc405421;
      27873: inst = 32'h8220000;
      27874: inst = 32'h10408000;
      27875: inst = 32'hc405422;
      27876: inst = 32'h8220000;
      27877: inst = 32'h10408000;
      27878: inst = 32'hc405436;
      27879: inst = 32'h8220000;
      27880: inst = 32'h10408000;
      27881: inst = 32'hc405437;
      27882: inst = 32'h8220000;
      27883: inst = 32'h10408000;
      27884: inst = 32'hc405438;
      27885: inst = 32'h8220000;
      27886: inst = 32'h10408000;
      27887: inst = 32'hc405439;
      27888: inst = 32'h8220000;
      27889: inst = 32'h10408000;
      27890: inst = 32'hc40543a;
      27891: inst = 32'h8220000;
      27892: inst = 32'h10408000;
      27893: inst = 32'hc40543b;
      27894: inst = 32'h8220000;
      27895: inst = 32'h10408000;
      27896: inst = 32'hc40543c;
      27897: inst = 32'h8220000;
      27898: inst = 32'h10408000;
      27899: inst = 32'hc40543d;
      27900: inst = 32'h8220000;
      27901: inst = 32'h10408000;
      27902: inst = 32'hc40543e;
      27903: inst = 32'h8220000;
      27904: inst = 32'h10408000;
      27905: inst = 32'hc40543f;
      27906: inst = 32'h8220000;
      27907: inst = 32'h10408000;
      27908: inst = 32'hc405440;
      27909: inst = 32'h8220000;
      27910: inst = 32'h10408000;
      27911: inst = 32'hc405441;
      27912: inst = 32'h8220000;
      27913: inst = 32'h10408000;
      27914: inst = 32'hc405442;
      27915: inst = 32'h8220000;
      27916: inst = 32'h10408000;
      27917: inst = 32'hc405443;
      27918: inst = 32'h8220000;
      27919: inst = 32'h10408000;
      27920: inst = 32'hc405444;
      27921: inst = 32'h8220000;
      27922: inst = 32'h10408000;
      27923: inst = 32'hc405445;
      27924: inst = 32'h8220000;
      27925: inst = 32'h10408000;
      27926: inst = 32'hc405446;
      27927: inst = 32'h8220000;
      27928: inst = 32'h10408000;
      27929: inst = 32'hc405447;
      27930: inst = 32'h8220000;
      27931: inst = 32'h10408000;
      27932: inst = 32'hc405448;
      27933: inst = 32'h8220000;
      27934: inst = 32'h10408000;
      27935: inst = 32'hc405449;
      27936: inst = 32'h8220000;
      27937: inst = 32'h10408000;
      27938: inst = 32'hc40547d;
      27939: inst = 32'h8220000;
      27940: inst = 32'h10408000;
      27941: inst = 32'hc40547e;
      27942: inst = 32'h8220000;
      27943: inst = 32'h10408000;
      27944: inst = 32'hc40547f;
      27945: inst = 32'h8220000;
      27946: inst = 32'h10408000;
      27947: inst = 32'hc405480;
      27948: inst = 32'h8220000;
      27949: inst = 32'h10408000;
      27950: inst = 32'hc405481;
      27951: inst = 32'h8220000;
      27952: inst = 32'h10408000;
      27953: inst = 32'hc405482;
      27954: inst = 32'h8220000;
      27955: inst = 32'h10408000;
      27956: inst = 32'hc405496;
      27957: inst = 32'h8220000;
      27958: inst = 32'h10408000;
      27959: inst = 32'hc405497;
      27960: inst = 32'h8220000;
      27961: inst = 32'h10408000;
      27962: inst = 32'hc405498;
      27963: inst = 32'h8220000;
      27964: inst = 32'h10408000;
      27965: inst = 32'hc405499;
      27966: inst = 32'h8220000;
      27967: inst = 32'h10408000;
      27968: inst = 32'hc40549a;
      27969: inst = 32'h8220000;
      27970: inst = 32'h10408000;
      27971: inst = 32'hc40549b;
      27972: inst = 32'h8220000;
      27973: inst = 32'h10408000;
      27974: inst = 32'hc40549c;
      27975: inst = 32'h8220000;
      27976: inst = 32'h10408000;
      27977: inst = 32'hc40549d;
      27978: inst = 32'h8220000;
      27979: inst = 32'h10408000;
      27980: inst = 32'hc40549e;
      27981: inst = 32'h8220000;
      27982: inst = 32'h10408000;
      27983: inst = 32'hc40549f;
      27984: inst = 32'h8220000;
      27985: inst = 32'h10408000;
      27986: inst = 32'hc4054a0;
      27987: inst = 32'h8220000;
      27988: inst = 32'h10408000;
      27989: inst = 32'hc4054a1;
      27990: inst = 32'h8220000;
      27991: inst = 32'h10408000;
      27992: inst = 32'hc4054a2;
      27993: inst = 32'h8220000;
      27994: inst = 32'h10408000;
      27995: inst = 32'hc4054a3;
      27996: inst = 32'h8220000;
      27997: inst = 32'h10408000;
      27998: inst = 32'hc4054a4;
      27999: inst = 32'h8220000;
      28000: inst = 32'h10408000;
      28001: inst = 32'hc4054a5;
      28002: inst = 32'h8220000;
      28003: inst = 32'h10408000;
      28004: inst = 32'hc4054a6;
      28005: inst = 32'h8220000;
      28006: inst = 32'h10408000;
      28007: inst = 32'hc4054a7;
      28008: inst = 32'h8220000;
      28009: inst = 32'h10408000;
      28010: inst = 32'hc4054a8;
      28011: inst = 32'h8220000;
      28012: inst = 32'h10408000;
      28013: inst = 32'hc4054a9;
      28014: inst = 32'h8220000;
      28015: inst = 32'h10408000;
      28016: inst = 32'hc4054dd;
      28017: inst = 32'h8220000;
      28018: inst = 32'h10408000;
      28019: inst = 32'hc4054de;
      28020: inst = 32'h8220000;
      28021: inst = 32'h10408000;
      28022: inst = 32'hc4054df;
      28023: inst = 32'h8220000;
      28024: inst = 32'h10408000;
      28025: inst = 32'hc4054e0;
      28026: inst = 32'h8220000;
      28027: inst = 32'h10408000;
      28028: inst = 32'hc4054e1;
      28029: inst = 32'h8220000;
      28030: inst = 32'h10408000;
      28031: inst = 32'hc4054e2;
      28032: inst = 32'h8220000;
      28033: inst = 32'h10408000;
      28034: inst = 32'hc4054f6;
      28035: inst = 32'h8220000;
      28036: inst = 32'h10408000;
      28037: inst = 32'hc4054f7;
      28038: inst = 32'h8220000;
      28039: inst = 32'h10408000;
      28040: inst = 32'hc4054f8;
      28041: inst = 32'h8220000;
      28042: inst = 32'h10408000;
      28043: inst = 32'hc4054f9;
      28044: inst = 32'h8220000;
      28045: inst = 32'h10408000;
      28046: inst = 32'hc4054fa;
      28047: inst = 32'h8220000;
      28048: inst = 32'h10408000;
      28049: inst = 32'hc4054fb;
      28050: inst = 32'h8220000;
      28051: inst = 32'h10408000;
      28052: inst = 32'hc4054fc;
      28053: inst = 32'h8220000;
      28054: inst = 32'h10408000;
      28055: inst = 32'hc4054fd;
      28056: inst = 32'h8220000;
      28057: inst = 32'h10408000;
      28058: inst = 32'hc4054fe;
      28059: inst = 32'h8220000;
      28060: inst = 32'h10408000;
      28061: inst = 32'hc4054ff;
      28062: inst = 32'h8220000;
      28063: inst = 32'h10408000;
      28064: inst = 32'hc405500;
      28065: inst = 32'h8220000;
      28066: inst = 32'h10408000;
      28067: inst = 32'hc405501;
      28068: inst = 32'h8220000;
      28069: inst = 32'h10408000;
      28070: inst = 32'hc405502;
      28071: inst = 32'h8220000;
      28072: inst = 32'h10408000;
      28073: inst = 32'hc405503;
      28074: inst = 32'h8220000;
      28075: inst = 32'h10408000;
      28076: inst = 32'hc405504;
      28077: inst = 32'h8220000;
      28078: inst = 32'h10408000;
      28079: inst = 32'hc405505;
      28080: inst = 32'h8220000;
      28081: inst = 32'h10408000;
      28082: inst = 32'hc405506;
      28083: inst = 32'h8220000;
      28084: inst = 32'h10408000;
      28085: inst = 32'hc405507;
      28086: inst = 32'h8220000;
      28087: inst = 32'h10408000;
      28088: inst = 32'hc405508;
      28089: inst = 32'h8220000;
      28090: inst = 32'h10408000;
      28091: inst = 32'hc405509;
      28092: inst = 32'h8220000;
      28093: inst = 32'h10408000;
      28094: inst = 32'hc40553d;
      28095: inst = 32'h8220000;
      28096: inst = 32'h10408000;
      28097: inst = 32'hc40553e;
      28098: inst = 32'h8220000;
      28099: inst = 32'h10408000;
      28100: inst = 32'hc40553f;
      28101: inst = 32'h8220000;
      28102: inst = 32'h10408000;
      28103: inst = 32'hc405540;
      28104: inst = 32'h8220000;
      28105: inst = 32'h10408000;
      28106: inst = 32'hc405541;
      28107: inst = 32'h8220000;
      28108: inst = 32'h10408000;
      28109: inst = 32'hc405542;
      28110: inst = 32'h8220000;
      28111: inst = 32'h10408000;
      28112: inst = 32'hc405556;
      28113: inst = 32'h8220000;
      28114: inst = 32'h10408000;
      28115: inst = 32'hc405557;
      28116: inst = 32'h8220000;
      28117: inst = 32'h10408000;
      28118: inst = 32'hc405558;
      28119: inst = 32'h8220000;
      28120: inst = 32'h10408000;
      28121: inst = 32'hc40559d;
      28122: inst = 32'h8220000;
      28123: inst = 32'h10408000;
      28124: inst = 32'hc40559e;
      28125: inst = 32'h8220000;
      28126: inst = 32'h10408000;
      28127: inst = 32'hc40559f;
      28128: inst = 32'h8220000;
      28129: inst = 32'h10408000;
      28130: inst = 32'hc4055a0;
      28131: inst = 32'h8220000;
      28132: inst = 32'h10408000;
      28133: inst = 32'hc4055a1;
      28134: inst = 32'h8220000;
      28135: inst = 32'h10408000;
      28136: inst = 32'hc4055a2;
      28137: inst = 32'h8220000;
      28138: inst = 32'h10408000;
      28139: inst = 32'hc4055b6;
      28140: inst = 32'h8220000;
      28141: inst = 32'h10408000;
      28142: inst = 32'hc4055b7;
      28143: inst = 32'h8220000;
      28144: inst = 32'h10408000;
      28145: inst = 32'hc4055b8;
      28146: inst = 32'h8220000;
      28147: inst = 32'h10408000;
      28148: inst = 32'hc4055fd;
      28149: inst = 32'h8220000;
      28150: inst = 32'h10408000;
      28151: inst = 32'hc4055fe;
      28152: inst = 32'h8220000;
      28153: inst = 32'h10408000;
      28154: inst = 32'hc4055ff;
      28155: inst = 32'h8220000;
      28156: inst = 32'h10408000;
      28157: inst = 32'hc405600;
      28158: inst = 32'h8220000;
      28159: inst = 32'h10408000;
      28160: inst = 32'hc405601;
      28161: inst = 32'h8220000;
      28162: inst = 32'h10408000;
      28163: inst = 32'hc405602;
      28164: inst = 32'h8220000;
      28165: inst = 32'h10408000;
      28166: inst = 32'hc405616;
      28167: inst = 32'h8220000;
      28168: inst = 32'h10408000;
      28169: inst = 32'hc405617;
      28170: inst = 32'h8220000;
      28171: inst = 32'h10408000;
      28172: inst = 32'hc405618;
      28173: inst = 32'h8220000;
      28174: inst = 32'h10408000;
      28175: inst = 32'hc40565d;
      28176: inst = 32'h8220000;
      28177: inst = 32'h10408000;
      28178: inst = 32'hc40565e;
      28179: inst = 32'h8220000;
      28180: inst = 32'h10408000;
      28181: inst = 32'hc40565f;
      28182: inst = 32'h8220000;
      28183: inst = 32'h10408000;
      28184: inst = 32'hc405660;
      28185: inst = 32'h8220000;
      28186: inst = 32'h10408000;
      28187: inst = 32'hc405661;
      28188: inst = 32'h8220000;
      28189: inst = 32'h10408000;
      28190: inst = 32'hc405662;
      28191: inst = 32'h8220000;
      28192: inst = 32'h10408000;
      28193: inst = 32'hc405676;
      28194: inst = 32'h8220000;
      28195: inst = 32'h10408000;
      28196: inst = 32'hc405677;
      28197: inst = 32'h8220000;
      28198: inst = 32'h10408000;
      28199: inst = 32'hc405678;
      28200: inst = 32'h8220000;
      28201: inst = 32'h10408000;
      28202: inst = 32'hc4056b7;
      28203: inst = 32'h8220000;
      28204: inst = 32'h10408000;
      28205: inst = 32'hc4056b8;
      28206: inst = 32'h8220000;
      28207: inst = 32'h10408000;
      28208: inst = 32'hc4056b9;
      28209: inst = 32'h8220000;
      28210: inst = 32'h10408000;
      28211: inst = 32'hc4056bd;
      28212: inst = 32'h8220000;
      28213: inst = 32'h10408000;
      28214: inst = 32'hc4056be;
      28215: inst = 32'h8220000;
      28216: inst = 32'h10408000;
      28217: inst = 32'hc4056bf;
      28218: inst = 32'h8220000;
      28219: inst = 32'h10408000;
      28220: inst = 32'hc4056c0;
      28221: inst = 32'h8220000;
      28222: inst = 32'h10408000;
      28223: inst = 32'hc4056c1;
      28224: inst = 32'h8220000;
      28225: inst = 32'h10408000;
      28226: inst = 32'hc4056c2;
      28227: inst = 32'h8220000;
      28228: inst = 32'h10408000;
      28229: inst = 32'hc4056c3;
      28230: inst = 32'h8220000;
      28231: inst = 32'h10408000;
      28232: inst = 32'hc4056c4;
      28233: inst = 32'h8220000;
      28234: inst = 32'h10408000;
      28235: inst = 32'hc4056c5;
      28236: inst = 32'h8220000;
      28237: inst = 32'h10408000;
      28238: inst = 32'hc4056c6;
      28239: inst = 32'h8220000;
      28240: inst = 32'h10408000;
      28241: inst = 32'hc4056c7;
      28242: inst = 32'h8220000;
      28243: inst = 32'h10408000;
      28244: inst = 32'hc4056c8;
      28245: inst = 32'h8220000;
      28246: inst = 32'h10408000;
      28247: inst = 32'hc4056c9;
      28248: inst = 32'h8220000;
      28249: inst = 32'h10408000;
      28250: inst = 32'hc4056d4;
      28251: inst = 32'h8220000;
      28252: inst = 32'h10408000;
      28253: inst = 32'hc4056d5;
      28254: inst = 32'h8220000;
      28255: inst = 32'h10408000;
      28256: inst = 32'hc4056d6;
      28257: inst = 32'h8220000;
      28258: inst = 32'h10408000;
      28259: inst = 32'hc4056d7;
      28260: inst = 32'h8220000;
      28261: inst = 32'h10408000;
      28262: inst = 32'hc4056d8;
      28263: inst = 32'h8220000;
      28264: inst = 32'h10408000;
      28265: inst = 32'hc4056d9;
      28266: inst = 32'h8220000;
      28267: inst = 32'h10408000;
      28268: inst = 32'hc4056da;
      28269: inst = 32'h8220000;
      28270: inst = 32'h10408000;
      28271: inst = 32'hc4056db;
      28272: inst = 32'h8220000;
      28273: inst = 32'h10408000;
      28274: inst = 32'hc4056dc;
      28275: inst = 32'h8220000;
      28276: inst = 32'h10408000;
      28277: inst = 32'hc4056dd;
      28278: inst = 32'h8220000;
      28279: inst = 32'h10408000;
      28280: inst = 32'hc4056de;
      28281: inst = 32'h8220000;
      28282: inst = 32'h10408000;
      28283: inst = 32'hc4056df;
      28284: inst = 32'h8220000;
      28285: inst = 32'h10408000;
      28286: inst = 32'hc4056e0;
      28287: inst = 32'h8220000;
      28288: inst = 32'h10408000;
      28289: inst = 32'hc4056e1;
      28290: inst = 32'h8220000;
      28291: inst = 32'h10408000;
      28292: inst = 32'hc4056e2;
      28293: inst = 32'h8220000;
      28294: inst = 32'h10408000;
      28295: inst = 32'hc4056e3;
      28296: inst = 32'h8220000;
      28297: inst = 32'h10408000;
      28298: inst = 32'hc4056e4;
      28299: inst = 32'h8220000;
      28300: inst = 32'h10408000;
      28301: inst = 32'hc4056e5;
      28302: inst = 32'h8220000;
      28303: inst = 32'h10408000;
      28304: inst = 32'hc4056e6;
      28305: inst = 32'h8220000;
      28306: inst = 32'h10408000;
      28307: inst = 32'hc4056e7;
      28308: inst = 32'h8220000;
      28309: inst = 32'h10408000;
      28310: inst = 32'hc4056e8;
      28311: inst = 32'h8220000;
      28312: inst = 32'h10408000;
      28313: inst = 32'hc4056e9;
      28314: inst = 32'h8220000;
      28315: inst = 32'h10408000;
      28316: inst = 32'hc4056ea;
      28317: inst = 32'h8220000;
      28318: inst = 32'h10408000;
      28319: inst = 32'hc4056eb;
      28320: inst = 32'h8220000;
      28321: inst = 32'h10408000;
      28322: inst = 32'hc4056ec;
      28323: inst = 32'h8220000;
      28324: inst = 32'h10408000;
      28325: inst = 32'hc4056ed;
      28326: inst = 32'h8220000;
      28327: inst = 32'h10408000;
      28328: inst = 32'hc4056ee;
      28329: inst = 32'h8220000;
      28330: inst = 32'h10408000;
      28331: inst = 32'hc4056ef;
      28332: inst = 32'h8220000;
      28333: inst = 32'h10408000;
      28334: inst = 32'hc4056f0;
      28335: inst = 32'h8220000;
      28336: inst = 32'h10408000;
      28337: inst = 32'hc4056f1;
      28338: inst = 32'h8220000;
      28339: inst = 32'h10408000;
      28340: inst = 32'hc4056f2;
      28341: inst = 32'h8220000;
      28342: inst = 32'h10408000;
      28343: inst = 32'hc4056f3;
      28344: inst = 32'h8220000;
      28345: inst = 32'h10408000;
      28346: inst = 32'hc4056f4;
      28347: inst = 32'h8220000;
      28348: inst = 32'h10408000;
      28349: inst = 32'hc4056f5;
      28350: inst = 32'h8220000;
      28351: inst = 32'h10408000;
      28352: inst = 32'hc4056f6;
      28353: inst = 32'h8220000;
      28354: inst = 32'h10408000;
      28355: inst = 32'hc4056f7;
      28356: inst = 32'h8220000;
      28357: inst = 32'h10408000;
      28358: inst = 32'hc4056f8;
      28359: inst = 32'h8220000;
      28360: inst = 32'h10408000;
      28361: inst = 32'hc4056f9;
      28362: inst = 32'h8220000;
      28363: inst = 32'h10408000;
      28364: inst = 32'hc4056fa;
      28365: inst = 32'h8220000;
      28366: inst = 32'h10408000;
      28367: inst = 32'hc4056fb;
      28368: inst = 32'h8220000;
      28369: inst = 32'h10408000;
      28370: inst = 32'hc4056fc;
      28371: inst = 32'h8220000;
      28372: inst = 32'h10408000;
      28373: inst = 32'hc4056fd;
      28374: inst = 32'h8220000;
      28375: inst = 32'h10408000;
      28376: inst = 32'hc405701;
      28377: inst = 32'h8220000;
      28378: inst = 32'h10408000;
      28379: inst = 32'hc405702;
      28380: inst = 32'h8220000;
      28381: inst = 32'h10408000;
      28382: inst = 32'hc405703;
      28383: inst = 32'h8220000;
      28384: inst = 32'h10408000;
      28385: inst = 32'hc405704;
      28386: inst = 32'h8220000;
      28387: inst = 32'h10408000;
      28388: inst = 32'hc405705;
      28389: inst = 32'h8220000;
      28390: inst = 32'h10408000;
      28391: inst = 32'hc405706;
      28392: inst = 32'h8220000;
      28393: inst = 32'h10408000;
      28394: inst = 32'hc405707;
      28395: inst = 32'h8220000;
      28396: inst = 32'h10408000;
      28397: inst = 32'hc405708;
      28398: inst = 32'h8220000;
      28399: inst = 32'h10408000;
      28400: inst = 32'hc405709;
      28401: inst = 32'h8220000;
      28402: inst = 32'h10408000;
      28403: inst = 32'hc40570a;
      28404: inst = 32'h8220000;
      28405: inst = 32'h10408000;
      28406: inst = 32'hc40570b;
      28407: inst = 32'h8220000;
      28408: inst = 32'h10408000;
      28409: inst = 32'hc40570c;
      28410: inst = 32'h8220000;
      28411: inst = 32'h10408000;
      28412: inst = 32'hc40570d;
      28413: inst = 32'h8220000;
      28414: inst = 32'h10408000;
      28415: inst = 32'hc40570e;
      28416: inst = 32'h8220000;
      28417: inst = 32'h10408000;
      28418: inst = 32'hc40570f;
      28419: inst = 32'h8220000;
      28420: inst = 32'h10408000;
      28421: inst = 32'hc405710;
      28422: inst = 32'h8220000;
      28423: inst = 32'h10408000;
      28424: inst = 32'hc405717;
      28425: inst = 32'h8220000;
      28426: inst = 32'h10408000;
      28427: inst = 32'hc405718;
      28428: inst = 32'h8220000;
      28429: inst = 32'h10408000;
      28430: inst = 32'hc405719;
      28431: inst = 32'h8220000;
      28432: inst = 32'h10408000;
      28433: inst = 32'hc40571d;
      28434: inst = 32'h8220000;
      28435: inst = 32'h10408000;
      28436: inst = 32'hc40571e;
      28437: inst = 32'h8220000;
      28438: inst = 32'h10408000;
      28439: inst = 32'hc40571f;
      28440: inst = 32'h8220000;
      28441: inst = 32'h10408000;
      28442: inst = 32'hc405720;
      28443: inst = 32'h8220000;
      28444: inst = 32'h10408000;
      28445: inst = 32'hc405721;
      28446: inst = 32'h8220000;
      28447: inst = 32'h10408000;
      28448: inst = 32'hc405722;
      28449: inst = 32'h8220000;
      28450: inst = 32'h10408000;
      28451: inst = 32'hc405723;
      28452: inst = 32'h8220000;
      28453: inst = 32'h10408000;
      28454: inst = 32'hc405724;
      28455: inst = 32'h8220000;
      28456: inst = 32'h10408000;
      28457: inst = 32'hc405725;
      28458: inst = 32'h8220000;
      28459: inst = 32'h10408000;
      28460: inst = 32'hc405726;
      28461: inst = 32'h8220000;
      28462: inst = 32'h10408000;
      28463: inst = 32'hc405727;
      28464: inst = 32'h8220000;
      28465: inst = 32'h10408000;
      28466: inst = 32'hc405728;
      28467: inst = 32'h8220000;
      28468: inst = 32'h10408000;
      28469: inst = 32'hc405729;
      28470: inst = 32'h8220000;
      28471: inst = 32'h10408000;
      28472: inst = 32'hc40572a;
      28473: inst = 32'h8220000;
      28474: inst = 32'h10408000;
      28475: inst = 32'hc40572b;
      28476: inst = 32'h8220000;
      28477: inst = 32'h10408000;
      28478: inst = 32'hc40572c;
      28479: inst = 32'h8220000;
      28480: inst = 32'h10408000;
      28481: inst = 32'hc40572d;
      28482: inst = 32'h8220000;
      28483: inst = 32'h10408000;
      28484: inst = 32'hc40572e;
      28485: inst = 32'h8220000;
      28486: inst = 32'h10408000;
      28487: inst = 32'hc40572f;
      28488: inst = 32'h8220000;
      28489: inst = 32'h10408000;
      28490: inst = 32'hc405730;
      28491: inst = 32'h8220000;
      28492: inst = 32'h10408000;
      28493: inst = 32'hc405731;
      28494: inst = 32'h8220000;
      28495: inst = 32'h10408000;
      28496: inst = 32'hc405732;
      28497: inst = 32'h8220000;
      28498: inst = 32'h10408000;
      28499: inst = 32'hc405733;
      28500: inst = 32'h8220000;
      28501: inst = 32'h10408000;
      28502: inst = 32'hc405734;
      28503: inst = 32'h8220000;
      28504: inst = 32'h10408000;
      28505: inst = 32'hc405735;
      28506: inst = 32'h8220000;
      28507: inst = 32'h10408000;
      28508: inst = 32'hc405736;
      28509: inst = 32'h8220000;
      28510: inst = 32'h10408000;
      28511: inst = 32'hc405737;
      28512: inst = 32'h8220000;
      28513: inst = 32'h10408000;
      28514: inst = 32'hc405738;
      28515: inst = 32'h8220000;
      28516: inst = 32'h10408000;
      28517: inst = 32'hc405739;
      28518: inst = 32'h8220000;
      28519: inst = 32'h10408000;
      28520: inst = 32'hc40573a;
      28521: inst = 32'h8220000;
      28522: inst = 32'h10408000;
      28523: inst = 32'hc40573b;
      28524: inst = 32'h8220000;
      28525: inst = 32'h10408000;
      28526: inst = 32'hc40573c;
      28527: inst = 32'h8220000;
      28528: inst = 32'h10408000;
      28529: inst = 32'hc40573d;
      28530: inst = 32'h8220000;
      28531: inst = 32'h10408000;
      28532: inst = 32'hc40573e;
      28533: inst = 32'h8220000;
      28534: inst = 32'h10408000;
      28535: inst = 32'hc40573f;
      28536: inst = 32'h8220000;
      28537: inst = 32'h10408000;
      28538: inst = 32'hc405740;
      28539: inst = 32'h8220000;
      28540: inst = 32'h10408000;
      28541: inst = 32'hc405741;
      28542: inst = 32'h8220000;
      28543: inst = 32'h10408000;
      28544: inst = 32'hc405742;
      28545: inst = 32'h8220000;
      28546: inst = 32'h10408000;
      28547: inst = 32'hc405743;
      28548: inst = 32'h8220000;
      28549: inst = 32'h10408000;
      28550: inst = 32'hc405744;
      28551: inst = 32'h8220000;
      28552: inst = 32'h10408000;
      28553: inst = 32'hc405745;
      28554: inst = 32'h8220000;
      28555: inst = 32'h10408000;
      28556: inst = 32'hc405746;
      28557: inst = 32'h8220000;
      28558: inst = 32'h10408000;
      28559: inst = 32'hc405747;
      28560: inst = 32'h8220000;
      28561: inst = 32'h10408000;
      28562: inst = 32'hc405748;
      28563: inst = 32'h8220000;
      28564: inst = 32'h10408000;
      28565: inst = 32'hc405749;
      28566: inst = 32'h8220000;
      28567: inst = 32'h10408000;
      28568: inst = 32'hc40574a;
      28569: inst = 32'h8220000;
      28570: inst = 32'h10408000;
      28571: inst = 32'hc40574b;
      28572: inst = 32'h8220000;
      28573: inst = 32'h10408000;
      28574: inst = 32'hc40574c;
      28575: inst = 32'h8220000;
      28576: inst = 32'h10408000;
      28577: inst = 32'hc40574d;
      28578: inst = 32'h8220000;
      28579: inst = 32'h10408000;
      28580: inst = 32'hc40574e;
      28581: inst = 32'h8220000;
      28582: inst = 32'h10408000;
      28583: inst = 32'hc40574f;
      28584: inst = 32'h8220000;
      28585: inst = 32'h10408000;
      28586: inst = 32'hc405750;
      28587: inst = 32'h8220000;
      28588: inst = 32'h10408000;
      28589: inst = 32'hc405751;
      28590: inst = 32'h8220000;
      28591: inst = 32'h10408000;
      28592: inst = 32'hc405752;
      28593: inst = 32'h8220000;
      28594: inst = 32'h10408000;
      28595: inst = 32'hc405753;
      28596: inst = 32'h8220000;
      28597: inst = 32'h10408000;
      28598: inst = 32'hc405754;
      28599: inst = 32'h8220000;
      28600: inst = 32'h10408000;
      28601: inst = 32'hc405755;
      28602: inst = 32'h8220000;
      28603: inst = 32'h10408000;
      28604: inst = 32'hc405756;
      28605: inst = 32'h8220000;
      28606: inst = 32'h10408000;
      28607: inst = 32'hc405757;
      28608: inst = 32'h8220000;
      28609: inst = 32'h10408000;
      28610: inst = 32'hc405758;
      28611: inst = 32'h8220000;
      28612: inst = 32'h10408000;
      28613: inst = 32'hc405759;
      28614: inst = 32'h8220000;
      28615: inst = 32'h10408000;
      28616: inst = 32'hc40575a;
      28617: inst = 32'h8220000;
      28618: inst = 32'h10408000;
      28619: inst = 32'hc40575b;
      28620: inst = 32'h8220000;
      28621: inst = 32'h10408000;
      28622: inst = 32'hc40575c;
      28623: inst = 32'h8220000;
      28624: inst = 32'h10408000;
      28625: inst = 32'hc40575d;
      28626: inst = 32'h8220000;
      28627: inst = 32'h10408000;
      28628: inst = 32'hc40575e;
      28629: inst = 32'h8220000;
      28630: inst = 32'h10408000;
      28631: inst = 32'hc405761;
      28632: inst = 32'h8220000;
      28633: inst = 32'h10408000;
      28634: inst = 32'hc405762;
      28635: inst = 32'h8220000;
      28636: inst = 32'h10408000;
      28637: inst = 32'hc405763;
      28638: inst = 32'h8220000;
      28639: inst = 32'h10408000;
      28640: inst = 32'hc405764;
      28641: inst = 32'h8220000;
      28642: inst = 32'h10408000;
      28643: inst = 32'hc405765;
      28644: inst = 32'h8220000;
      28645: inst = 32'h10408000;
      28646: inst = 32'hc405766;
      28647: inst = 32'h8220000;
      28648: inst = 32'h10408000;
      28649: inst = 32'hc405767;
      28650: inst = 32'h8220000;
      28651: inst = 32'h10408000;
      28652: inst = 32'hc405768;
      28653: inst = 32'h8220000;
      28654: inst = 32'h10408000;
      28655: inst = 32'hc405769;
      28656: inst = 32'h8220000;
      28657: inst = 32'h10408000;
      28658: inst = 32'hc40576a;
      28659: inst = 32'h8220000;
      28660: inst = 32'h10408000;
      28661: inst = 32'hc40576b;
      28662: inst = 32'h8220000;
      28663: inst = 32'h10408000;
      28664: inst = 32'hc40576c;
      28665: inst = 32'h8220000;
      28666: inst = 32'h10408000;
      28667: inst = 32'hc40576d;
      28668: inst = 32'h8220000;
      28669: inst = 32'h10408000;
      28670: inst = 32'hc40576e;
      28671: inst = 32'h8220000;
      28672: inst = 32'h10408000;
      28673: inst = 32'hc40576f;
      28674: inst = 32'h8220000;
      28675: inst = 32'h10408000;
      28676: inst = 32'hc405770;
      28677: inst = 32'h8220000;
      28678: inst = 32'h10408000;
      28679: inst = 32'hc40577d;
      28680: inst = 32'h8220000;
      28681: inst = 32'h10408000;
      28682: inst = 32'hc40577e;
      28683: inst = 32'h8220000;
      28684: inst = 32'h10408000;
      28685: inst = 32'hc40577f;
      28686: inst = 32'h8220000;
      28687: inst = 32'h10408000;
      28688: inst = 32'hc405780;
      28689: inst = 32'h8220000;
      28690: inst = 32'h10408000;
      28691: inst = 32'hc405781;
      28692: inst = 32'h8220000;
      28693: inst = 32'h10408000;
      28694: inst = 32'hc405782;
      28695: inst = 32'h8220000;
      28696: inst = 32'h10408000;
      28697: inst = 32'hc405783;
      28698: inst = 32'h8220000;
      28699: inst = 32'h10408000;
      28700: inst = 32'hc405784;
      28701: inst = 32'h8220000;
      28702: inst = 32'h10408000;
      28703: inst = 32'hc405785;
      28704: inst = 32'h8220000;
      28705: inst = 32'h10408000;
      28706: inst = 32'hc405786;
      28707: inst = 32'h8220000;
      28708: inst = 32'h10408000;
      28709: inst = 32'hc405787;
      28710: inst = 32'h8220000;
      28711: inst = 32'h10408000;
      28712: inst = 32'hc405788;
      28713: inst = 32'h8220000;
      28714: inst = 32'h10408000;
      28715: inst = 32'hc405789;
      28716: inst = 32'h8220000;
      28717: inst = 32'h10408000;
      28718: inst = 32'hc40578a;
      28719: inst = 32'h8220000;
      28720: inst = 32'h10408000;
      28721: inst = 32'hc40578b;
      28722: inst = 32'h8220000;
      28723: inst = 32'h10408000;
      28724: inst = 32'hc40578c;
      28725: inst = 32'h8220000;
      28726: inst = 32'h10408000;
      28727: inst = 32'hc40578d;
      28728: inst = 32'h8220000;
      28729: inst = 32'h10408000;
      28730: inst = 32'hc40578e;
      28731: inst = 32'h8220000;
      28732: inst = 32'h10408000;
      28733: inst = 32'hc40578f;
      28734: inst = 32'h8220000;
      28735: inst = 32'h10408000;
      28736: inst = 32'hc405790;
      28737: inst = 32'h8220000;
      28738: inst = 32'h10408000;
      28739: inst = 32'hc405791;
      28740: inst = 32'h8220000;
      28741: inst = 32'h10408000;
      28742: inst = 32'hc405792;
      28743: inst = 32'h8220000;
      28744: inst = 32'h10408000;
      28745: inst = 32'hc405793;
      28746: inst = 32'h8220000;
      28747: inst = 32'h10408000;
      28748: inst = 32'hc405794;
      28749: inst = 32'h8220000;
      28750: inst = 32'h10408000;
      28751: inst = 32'hc405795;
      28752: inst = 32'h8220000;
      28753: inst = 32'h10408000;
      28754: inst = 32'hc405796;
      28755: inst = 32'h8220000;
      28756: inst = 32'h10408000;
      28757: inst = 32'hc405797;
      28758: inst = 32'h8220000;
      28759: inst = 32'h10408000;
      28760: inst = 32'hc405798;
      28761: inst = 32'h8220000;
      28762: inst = 32'h10408000;
      28763: inst = 32'hc405799;
      28764: inst = 32'h8220000;
      28765: inst = 32'h10408000;
      28766: inst = 32'hc40579a;
      28767: inst = 32'h8220000;
      28768: inst = 32'h10408000;
      28769: inst = 32'hc40579b;
      28770: inst = 32'h8220000;
      28771: inst = 32'h10408000;
      28772: inst = 32'hc40579c;
      28773: inst = 32'h8220000;
      28774: inst = 32'h10408000;
      28775: inst = 32'hc40579d;
      28776: inst = 32'h8220000;
      28777: inst = 32'h10408000;
      28778: inst = 32'hc40579e;
      28779: inst = 32'h8220000;
      28780: inst = 32'h10408000;
      28781: inst = 32'hc40579f;
      28782: inst = 32'h8220000;
      28783: inst = 32'h10408000;
      28784: inst = 32'hc4057a0;
      28785: inst = 32'h8220000;
      28786: inst = 32'h10408000;
      28787: inst = 32'hc4057a1;
      28788: inst = 32'h8220000;
      28789: inst = 32'h10408000;
      28790: inst = 32'hc4057a2;
      28791: inst = 32'h8220000;
      28792: inst = 32'h10408000;
      28793: inst = 32'hc4057a3;
      28794: inst = 32'h8220000;
      28795: inst = 32'h10408000;
      28796: inst = 32'hc4057a4;
      28797: inst = 32'h8220000;
      28798: inst = 32'h10408000;
      28799: inst = 32'hc4057a5;
      28800: inst = 32'h8220000;
      28801: inst = 32'h10408000;
      28802: inst = 32'hc4057a6;
      28803: inst = 32'h8220000;
      28804: inst = 32'h10408000;
      28805: inst = 32'hc4057a7;
      28806: inst = 32'h8220000;
      28807: inst = 32'h10408000;
      28808: inst = 32'hc4057a8;
      28809: inst = 32'h8220000;
      28810: inst = 32'h10408000;
      28811: inst = 32'hc4057a9;
      28812: inst = 32'h8220000;
      28813: inst = 32'h10408000;
      28814: inst = 32'hc4057aa;
      28815: inst = 32'h8220000;
      28816: inst = 32'h10408000;
      28817: inst = 32'hc4057ab;
      28818: inst = 32'h8220000;
      28819: inst = 32'h10408000;
      28820: inst = 32'hc4057ac;
      28821: inst = 32'h8220000;
      28822: inst = 32'h10408000;
      28823: inst = 32'hc4057ad;
      28824: inst = 32'h8220000;
      28825: inst = 32'h10408000;
      28826: inst = 32'hc4057ae;
      28827: inst = 32'h8220000;
      28828: inst = 32'h10408000;
      28829: inst = 32'hc4057af;
      28830: inst = 32'h8220000;
      28831: inst = 32'h10408000;
      28832: inst = 32'hc4057b0;
      28833: inst = 32'h8220000;
      28834: inst = 32'h10408000;
      28835: inst = 32'hc4057b1;
      28836: inst = 32'h8220000;
      28837: inst = 32'h10408000;
      28838: inst = 32'hc4057b2;
      28839: inst = 32'h8220000;
      28840: inst = 32'h10408000;
      28841: inst = 32'hc4057b3;
      28842: inst = 32'h8220000;
      28843: inst = 32'h10408000;
      28844: inst = 32'hc4057b4;
      28845: inst = 32'h8220000;
      28846: inst = 32'h10408000;
      28847: inst = 32'hc4057b5;
      28848: inst = 32'h8220000;
      28849: inst = 32'h10408000;
      28850: inst = 32'hc4057b6;
      28851: inst = 32'h8220000;
      28852: inst = 32'h10408000;
      28853: inst = 32'hc4057b7;
      28854: inst = 32'h8220000;
      28855: inst = 32'h10408000;
      28856: inst = 32'hc4057b8;
      28857: inst = 32'h8220000;
      28858: inst = 32'h10408000;
      28859: inst = 32'hc4057b9;
      28860: inst = 32'h8220000;
      28861: inst = 32'h10408000;
      28862: inst = 32'hc4057ba;
      28863: inst = 32'h8220000;
      28864: inst = 32'h10408000;
      28865: inst = 32'hc4057bb;
      28866: inst = 32'h8220000;
      28867: inst = 32'h10408000;
      28868: inst = 32'hc4057bc;
      28869: inst = 32'h8220000;
      28870: inst = 32'h10408000;
      28871: inst = 32'hc4057bd;
      28872: inst = 32'h8220000;
      28873: inst = 32'h10408000;
      28874: inst = 32'hc4057be;
      28875: inst = 32'h8220000;
      28876: inst = 32'h10408000;
      28877: inst = 32'hc4057c1;
      28878: inst = 32'h8220000;
      28879: inst = 32'h10408000;
      28880: inst = 32'hc4057c2;
      28881: inst = 32'h8220000;
      28882: inst = 32'h10408000;
      28883: inst = 32'hc4057c3;
      28884: inst = 32'h8220000;
      28885: inst = 32'h10408000;
      28886: inst = 32'hc4057c4;
      28887: inst = 32'h8220000;
      28888: inst = 32'h10408000;
      28889: inst = 32'hc4057c5;
      28890: inst = 32'h8220000;
      28891: inst = 32'h10408000;
      28892: inst = 32'hc4057c6;
      28893: inst = 32'h8220000;
      28894: inst = 32'h10408000;
      28895: inst = 32'hc4057c7;
      28896: inst = 32'h8220000;
      28897: inst = 32'h10408000;
      28898: inst = 32'hc4057c8;
      28899: inst = 32'h8220000;
      28900: inst = 32'h10408000;
      28901: inst = 32'hc4057c9;
      28902: inst = 32'h8220000;
      28903: inst = 32'h10408000;
      28904: inst = 32'hc4057ca;
      28905: inst = 32'h8220000;
      28906: inst = 32'h10408000;
      28907: inst = 32'hc4057cb;
      28908: inst = 32'h8220000;
      28909: inst = 32'h10408000;
      28910: inst = 32'hc4057cc;
      28911: inst = 32'h8220000;
      28912: inst = 32'h10408000;
      28913: inst = 32'hc4057cd;
      28914: inst = 32'h8220000;
      28915: inst = 32'h10408000;
      28916: inst = 32'hc4057ce;
      28917: inst = 32'h8220000;
      28918: inst = 32'h10408000;
      28919: inst = 32'hc4057cf;
      28920: inst = 32'h8220000;
      28921: inst = 32'h10408000;
      28922: inst = 32'hc4057d0;
      28923: inst = 32'h8220000;
      28924: inst = 32'h10408000;
      28925: inst = 32'hc4057dd;
      28926: inst = 32'h8220000;
      28927: inst = 32'h10408000;
      28928: inst = 32'hc4057de;
      28929: inst = 32'h8220000;
      28930: inst = 32'h10408000;
      28931: inst = 32'hc4057df;
      28932: inst = 32'h8220000;
      28933: inst = 32'hc20eeb6;
      28934: inst = 32'h10408000;
      28935: inst = 32'hc403fe3;
      28936: inst = 32'h8220000;
      28937: inst = 32'h10408000;
      28938: inst = 32'hc404043;
      28939: inst = 32'h8220000;
      28940: inst = 32'h10408000;
      28941: inst = 32'hc4040a3;
      28942: inst = 32'h8220000;
      28943: inst = 32'h10408000;
      28944: inst = 32'hc404103;
      28945: inst = 32'h8220000;
      28946: inst = 32'h10408000;
      28947: inst = 32'hc40410e;
      28948: inst = 32'h8220000;
      28949: inst = 32'h10408000;
      28950: inst = 32'hc40410f;
      28951: inst = 32'h8220000;
      28952: inst = 32'h10408000;
      28953: inst = 32'hc404110;
      28954: inst = 32'h8220000;
      28955: inst = 32'h10408000;
      28956: inst = 32'hc404111;
      28957: inst = 32'h8220000;
      28958: inst = 32'h10408000;
      28959: inst = 32'hc404112;
      28960: inst = 32'h8220000;
      28961: inst = 32'h10408000;
      28962: inst = 32'hc404115;
      28963: inst = 32'h8220000;
      28964: inst = 32'h10408000;
      28965: inst = 32'hc404118;
      28966: inst = 32'h8220000;
      28967: inst = 32'h10408000;
      28968: inst = 32'hc404119;
      28969: inst = 32'h8220000;
      28970: inst = 32'h10408000;
      28971: inst = 32'hc40411a;
      28972: inst = 32'h8220000;
      28973: inst = 32'h10408000;
      28974: inst = 32'hc40411b;
      28975: inst = 32'h8220000;
      28976: inst = 32'h10408000;
      28977: inst = 32'hc40411c;
      28978: inst = 32'h8220000;
      28979: inst = 32'h10408000;
      28980: inst = 32'hc40411d;
      28981: inst = 32'h8220000;
      28982: inst = 32'h10408000;
      28983: inst = 32'hc40411e;
      28984: inst = 32'h8220000;
      28985: inst = 32'h10408000;
      28986: inst = 32'hc40411f;
      28987: inst = 32'h8220000;
      28988: inst = 32'h10408000;
      28989: inst = 32'hc404120;
      28990: inst = 32'h8220000;
      28991: inst = 32'h10408000;
      28992: inst = 32'hc404121;
      28993: inst = 32'h8220000;
      28994: inst = 32'h10408000;
      28995: inst = 32'hc404122;
      28996: inst = 32'h8220000;
      28997: inst = 32'h10408000;
      28998: inst = 32'hc404123;
      28999: inst = 32'h8220000;
      29000: inst = 32'h10408000;
      29001: inst = 32'hc404124;
      29002: inst = 32'h8220000;
      29003: inst = 32'h10408000;
      29004: inst = 32'hc404125;
      29005: inst = 32'h8220000;
      29006: inst = 32'h10408000;
      29007: inst = 32'hc404126;
      29008: inst = 32'h8220000;
      29009: inst = 32'h10408000;
      29010: inst = 32'hc404127;
      29011: inst = 32'h8220000;
      29012: inst = 32'h10408000;
      29013: inst = 32'hc404128;
      29014: inst = 32'h8220000;
      29015: inst = 32'h10408000;
      29016: inst = 32'hc404129;
      29017: inst = 32'h8220000;
      29018: inst = 32'h10408000;
      29019: inst = 32'hc40412a;
      29020: inst = 32'h8220000;
      29021: inst = 32'h10408000;
      29022: inst = 32'hc40412b;
      29023: inst = 32'h8220000;
      29024: inst = 32'h10408000;
      29025: inst = 32'hc40412c;
      29026: inst = 32'h8220000;
      29027: inst = 32'h10408000;
      29028: inst = 32'hc40412d;
      29029: inst = 32'h8220000;
      29030: inst = 32'h10408000;
      29031: inst = 32'hc40412e;
      29032: inst = 32'h8220000;
      29033: inst = 32'h10408000;
      29034: inst = 32'hc40412f;
      29035: inst = 32'h8220000;
      29036: inst = 32'h10408000;
      29037: inst = 32'hc404130;
      29038: inst = 32'h8220000;
      29039: inst = 32'h10408000;
      29040: inst = 32'hc404131;
      29041: inst = 32'h8220000;
      29042: inst = 32'h10408000;
      29043: inst = 32'hc404132;
      29044: inst = 32'h8220000;
      29045: inst = 32'h10408000;
      29046: inst = 32'hc404133;
      29047: inst = 32'h8220000;
      29048: inst = 32'h10408000;
      29049: inst = 32'hc404134;
      29050: inst = 32'h8220000;
      29051: inst = 32'h10408000;
      29052: inst = 32'hc404135;
      29053: inst = 32'h8220000;
      29054: inst = 32'h10408000;
      29055: inst = 32'hc404136;
      29056: inst = 32'h8220000;
      29057: inst = 32'h10408000;
      29058: inst = 32'hc404137;
      29059: inst = 32'h8220000;
      29060: inst = 32'h10408000;
      29061: inst = 32'hc404138;
      29062: inst = 32'h8220000;
      29063: inst = 32'h10408000;
      29064: inst = 32'hc404139;
      29065: inst = 32'h8220000;
      29066: inst = 32'h10408000;
      29067: inst = 32'hc40413a;
      29068: inst = 32'h8220000;
      29069: inst = 32'h10408000;
      29070: inst = 32'hc40413b;
      29071: inst = 32'h8220000;
      29072: inst = 32'h10408000;
      29073: inst = 32'hc40413c;
      29074: inst = 32'h8220000;
      29075: inst = 32'h10408000;
      29076: inst = 32'hc40413d;
      29077: inst = 32'h8220000;
      29078: inst = 32'h10408000;
      29079: inst = 32'hc40413e;
      29080: inst = 32'h8220000;
      29081: inst = 32'h10408000;
      29082: inst = 32'hc40413f;
      29083: inst = 32'h8220000;
      29084: inst = 32'h10408000;
      29085: inst = 32'hc404140;
      29086: inst = 32'h8220000;
      29087: inst = 32'h10408000;
      29088: inst = 32'hc404141;
      29089: inst = 32'h8220000;
      29090: inst = 32'h10408000;
      29091: inst = 32'hc404142;
      29092: inst = 32'h8220000;
      29093: inst = 32'h10408000;
      29094: inst = 32'hc404143;
      29095: inst = 32'h8220000;
      29096: inst = 32'h10408000;
      29097: inst = 32'hc404144;
      29098: inst = 32'h8220000;
      29099: inst = 32'h10408000;
      29100: inst = 32'hc404145;
      29101: inst = 32'h8220000;
      29102: inst = 32'h10408000;
      29103: inst = 32'hc404146;
      29104: inst = 32'h8220000;
      29105: inst = 32'h10408000;
      29106: inst = 32'hc404147;
      29107: inst = 32'h8220000;
      29108: inst = 32'h10408000;
      29109: inst = 32'hc404148;
      29110: inst = 32'h8220000;
      29111: inst = 32'h10408000;
      29112: inst = 32'hc404149;
      29113: inst = 32'h8220000;
      29114: inst = 32'h10408000;
      29115: inst = 32'hc40414a;
      29116: inst = 32'h8220000;
      29117: inst = 32'h10408000;
      29118: inst = 32'hc40414b;
      29119: inst = 32'h8220000;
      29120: inst = 32'h10408000;
      29121: inst = 32'hc40414f;
      29122: inst = 32'h8220000;
      29123: inst = 32'h10408000;
      29124: inst = 32'hc404150;
      29125: inst = 32'h8220000;
      29126: inst = 32'h10408000;
      29127: inst = 32'hc404163;
      29128: inst = 32'h8220000;
      29129: inst = 32'h10408000;
      29130: inst = 32'hc40416e;
      29131: inst = 32'h8220000;
      29132: inst = 32'h10408000;
      29133: inst = 32'hc40416f;
      29134: inst = 32'h8220000;
      29135: inst = 32'h10408000;
      29136: inst = 32'hc404170;
      29137: inst = 32'h8220000;
      29138: inst = 32'h10408000;
      29139: inst = 32'hc404171;
      29140: inst = 32'h8220000;
      29141: inst = 32'h10408000;
      29142: inst = 32'hc404172;
      29143: inst = 32'h8220000;
      29144: inst = 32'h10408000;
      29145: inst = 32'hc404173;
      29146: inst = 32'h8220000;
      29147: inst = 32'h10408000;
      29148: inst = 32'hc404174;
      29149: inst = 32'h8220000;
      29150: inst = 32'h10408000;
      29151: inst = 32'hc404175;
      29152: inst = 32'h8220000;
      29153: inst = 32'h10408000;
      29154: inst = 32'hc404178;
      29155: inst = 32'h8220000;
      29156: inst = 32'h10408000;
      29157: inst = 32'hc404179;
      29158: inst = 32'h8220000;
      29159: inst = 32'h10408000;
      29160: inst = 32'hc40417a;
      29161: inst = 32'h8220000;
      29162: inst = 32'h10408000;
      29163: inst = 32'hc40417c;
      29164: inst = 32'h8220000;
      29165: inst = 32'h10408000;
      29166: inst = 32'hc40417d;
      29167: inst = 32'h8220000;
      29168: inst = 32'h10408000;
      29169: inst = 32'hc40417e;
      29170: inst = 32'h8220000;
      29171: inst = 32'h10408000;
      29172: inst = 32'hc40417f;
      29173: inst = 32'h8220000;
      29174: inst = 32'h10408000;
      29175: inst = 32'hc404180;
      29176: inst = 32'h8220000;
      29177: inst = 32'h10408000;
      29178: inst = 32'hc404181;
      29179: inst = 32'h8220000;
      29180: inst = 32'h10408000;
      29181: inst = 32'hc404182;
      29182: inst = 32'h8220000;
      29183: inst = 32'h10408000;
      29184: inst = 32'hc404183;
      29185: inst = 32'h8220000;
      29186: inst = 32'h10408000;
      29187: inst = 32'hc404184;
      29188: inst = 32'h8220000;
      29189: inst = 32'h10408000;
      29190: inst = 32'hc404185;
      29191: inst = 32'h8220000;
      29192: inst = 32'h10408000;
      29193: inst = 32'hc404186;
      29194: inst = 32'h8220000;
      29195: inst = 32'h10408000;
      29196: inst = 32'hc404187;
      29197: inst = 32'h8220000;
      29198: inst = 32'h10408000;
      29199: inst = 32'hc404188;
      29200: inst = 32'h8220000;
      29201: inst = 32'h10408000;
      29202: inst = 32'hc404189;
      29203: inst = 32'h8220000;
      29204: inst = 32'h10408000;
      29205: inst = 32'hc40418a;
      29206: inst = 32'h8220000;
      29207: inst = 32'h10408000;
      29208: inst = 32'hc40418b;
      29209: inst = 32'h8220000;
      29210: inst = 32'h10408000;
      29211: inst = 32'hc40418c;
      29212: inst = 32'h8220000;
      29213: inst = 32'h10408000;
      29214: inst = 32'hc40418d;
      29215: inst = 32'h8220000;
      29216: inst = 32'h10408000;
      29217: inst = 32'hc40418e;
      29218: inst = 32'h8220000;
      29219: inst = 32'h10408000;
      29220: inst = 32'hc40418f;
      29221: inst = 32'h8220000;
      29222: inst = 32'h10408000;
      29223: inst = 32'hc404190;
      29224: inst = 32'h8220000;
      29225: inst = 32'h10408000;
      29226: inst = 32'hc404191;
      29227: inst = 32'h8220000;
      29228: inst = 32'h10408000;
      29229: inst = 32'hc404192;
      29230: inst = 32'h8220000;
      29231: inst = 32'h10408000;
      29232: inst = 32'hc404193;
      29233: inst = 32'h8220000;
      29234: inst = 32'h10408000;
      29235: inst = 32'hc404194;
      29236: inst = 32'h8220000;
      29237: inst = 32'h10408000;
      29238: inst = 32'hc404195;
      29239: inst = 32'h8220000;
      29240: inst = 32'h10408000;
      29241: inst = 32'hc404196;
      29242: inst = 32'h8220000;
      29243: inst = 32'h10408000;
      29244: inst = 32'hc404197;
      29245: inst = 32'h8220000;
      29246: inst = 32'h10408000;
      29247: inst = 32'hc404198;
      29248: inst = 32'h8220000;
      29249: inst = 32'h10408000;
      29250: inst = 32'hc404199;
      29251: inst = 32'h8220000;
      29252: inst = 32'h10408000;
      29253: inst = 32'hc40419a;
      29254: inst = 32'h8220000;
      29255: inst = 32'h10408000;
      29256: inst = 32'hc40419b;
      29257: inst = 32'h8220000;
      29258: inst = 32'h10408000;
      29259: inst = 32'hc40419c;
      29260: inst = 32'h8220000;
      29261: inst = 32'h10408000;
      29262: inst = 32'hc40419d;
      29263: inst = 32'h8220000;
      29264: inst = 32'h10408000;
      29265: inst = 32'hc40419e;
      29266: inst = 32'h8220000;
      29267: inst = 32'h10408000;
      29268: inst = 32'hc40419f;
      29269: inst = 32'h8220000;
      29270: inst = 32'h10408000;
      29271: inst = 32'hc4041a0;
      29272: inst = 32'h8220000;
      29273: inst = 32'h10408000;
      29274: inst = 32'hc4041a1;
      29275: inst = 32'h8220000;
      29276: inst = 32'h10408000;
      29277: inst = 32'hc4041a2;
      29278: inst = 32'h8220000;
      29279: inst = 32'h10408000;
      29280: inst = 32'hc4041a3;
      29281: inst = 32'h8220000;
      29282: inst = 32'h10408000;
      29283: inst = 32'hc4041a4;
      29284: inst = 32'h8220000;
      29285: inst = 32'h10408000;
      29286: inst = 32'hc4041a5;
      29287: inst = 32'h8220000;
      29288: inst = 32'h10408000;
      29289: inst = 32'hc4041a6;
      29290: inst = 32'h8220000;
      29291: inst = 32'h10408000;
      29292: inst = 32'hc4041a7;
      29293: inst = 32'h8220000;
      29294: inst = 32'h10408000;
      29295: inst = 32'hc4041a8;
      29296: inst = 32'h8220000;
      29297: inst = 32'h10408000;
      29298: inst = 32'hc4041a9;
      29299: inst = 32'h8220000;
      29300: inst = 32'h10408000;
      29301: inst = 32'hc4041aa;
      29302: inst = 32'h8220000;
      29303: inst = 32'h10408000;
      29304: inst = 32'hc4041ab;
      29305: inst = 32'h8220000;
      29306: inst = 32'h10408000;
      29307: inst = 32'hc4041af;
      29308: inst = 32'h8220000;
      29309: inst = 32'h10408000;
      29310: inst = 32'hc4041b5;
      29311: inst = 32'h8220000;
      29312: inst = 32'h10408000;
      29313: inst = 32'hc4041c3;
      29314: inst = 32'h8220000;
      29315: inst = 32'h10408000;
      29316: inst = 32'hc4041cd;
      29317: inst = 32'h8220000;
      29318: inst = 32'h10408000;
      29319: inst = 32'hc4041ce;
      29320: inst = 32'h8220000;
      29321: inst = 32'h10408000;
      29322: inst = 32'hc4041cf;
      29323: inst = 32'h8220000;
      29324: inst = 32'h10408000;
      29325: inst = 32'hc4041d2;
      29326: inst = 32'h8220000;
      29327: inst = 32'h10408000;
      29328: inst = 32'hc4041d3;
      29329: inst = 32'h8220000;
      29330: inst = 32'h10408000;
      29331: inst = 32'hc4041d4;
      29332: inst = 32'h8220000;
      29333: inst = 32'h10408000;
      29334: inst = 32'hc4041d5;
      29335: inst = 32'h8220000;
      29336: inst = 32'h10408000;
      29337: inst = 32'hc4041d9;
      29338: inst = 32'h8220000;
      29339: inst = 32'h10408000;
      29340: inst = 32'hc4041da;
      29341: inst = 32'h8220000;
      29342: inst = 32'h10408000;
      29343: inst = 32'hc4041dd;
      29344: inst = 32'h8220000;
      29345: inst = 32'h10408000;
      29346: inst = 32'hc4041de;
      29347: inst = 32'h8220000;
      29348: inst = 32'h10408000;
      29349: inst = 32'hc4041df;
      29350: inst = 32'h8220000;
      29351: inst = 32'h10408000;
      29352: inst = 32'hc4041e0;
      29353: inst = 32'h8220000;
      29354: inst = 32'h10408000;
      29355: inst = 32'hc4041e1;
      29356: inst = 32'h8220000;
      29357: inst = 32'h10408000;
      29358: inst = 32'hc4041e2;
      29359: inst = 32'h8220000;
      29360: inst = 32'h10408000;
      29361: inst = 32'hc4041e3;
      29362: inst = 32'h8220000;
      29363: inst = 32'h10408000;
      29364: inst = 32'hc4041e4;
      29365: inst = 32'h8220000;
      29366: inst = 32'h10408000;
      29367: inst = 32'hc4041e5;
      29368: inst = 32'h8220000;
      29369: inst = 32'h10408000;
      29370: inst = 32'hc4041e6;
      29371: inst = 32'h8220000;
      29372: inst = 32'h10408000;
      29373: inst = 32'hc4041e7;
      29374: inst = 32'h8220000;
      29375: inst = 32'h10408000;
      29376: inst = 32'hc4041e8;
      29377: inst = 32'h8220000;
      29378: inst = 32'h10408000;
      29379: inst = 32'hc4041e9;
      29380: inst = 32'h8220000;
      29381: inst = 32'h10408000;
      29382: inst = 32'hc4041ea;
      29383: inst = 32'h8220000;
      29384: inst = 32'h10408000;
      29385: inst = 32'hc4041eb;
      29386: inst = 32'h8220000;
      29387: inst = 32'h10408000;
      29388: inst = 32'hc4041ec;
      29389: inst = 32'h8220000;
      29390: inst = 32'h10408000;
      29391: inst = 32'hc4041ed;
      29392: inst = 32'h8220000;
      29393: inst = 32'h10408000;
      29394: inst = 32'hc4041ee;
      29395: inst = 32'h8220000;
      29396: inst = 32'h10408000;
      29397: inst = 32'hc4041ef;
      29398: inst = 32'h8220000;
      29399: inst = 32'h10408000;
      29400: inst = 32'hc4041f0;
      29401: inst = 32'h8220000;
      29402: inst = 32'h10408000;
      29403: inst = 32'hc4041f1;
      29404: inst = 32'h8220000;
      29405: inst = 32'h10408000;
      29406: inst = 32'hc4041f2;
      29407: inst = 32'h8220000;
      29408: inst = 32'h10408000;
      29409: inst = 32'hc4041f3;
      29410: inst = 32'h8220000;
      29411: inst = 32'h10408000;
      29412: inst = 32'hc4041f4;
      29413: inst = 32'h8220000;
      29414: inst = 32'h10408000;
      29415: inst = 32'hc4041f5;
      29416: inst = 32'h8220000;
      29417: inst = 32'h10408000;
      29418: inst = 32'hc4041f6;
      29419: inst = 32'h8220000;
      29420: inst = 32'h10408000;
      29421: inst = 32'hc4041f7;
      29422: inst = 32'h8220000;
      29423: inst = 32'h10408000;
      29424: inst = 32'hc4041f8;
      29425: inst = 32'h8220000;
      29426: inst = 32'h10408000;
      29427: inst = 32'hc4041f9;
      29428: inst = 32'h8220000;
      29429: inst = 32'h10408000;
      29430: inst = 32'hc4041fa;
      29431: inst = 32'h8220000;
      29432: inst = 32'h10408000;
      29433: inst = 32'hc4041fb;
      29434: inst = 32'h8220000;
      29435: inst = 32'h10408000;
      29436: inst = 32'hc4041fc;
      29437: inst = 32'h8220000;
      29438: inst = 32'h10408000;
      29439: inst = 32'hc4041fd;
      29440: inst = 32'h8220000;
      29441: inst = 32'h10408000;
      29442: inst = 32'hc4041fe;
      29443: inst = 32'h8220000;
      29444: inst = 32'h10408000;
      29445: inst = 32'hc4041ff;
      29446: inst = 32'h8220000;
      29447: inst = 32'h10408000;
      29448: inst = 32'hc404200;
      29449: inst = 32'h8220000;
      29450: inst = 32'h10408000;
      29451: inst = 32'hc404201;
      29452: inst = 32'h8220000;
      29453: inst = 32'h10408000;
      29454: inst = 32'hc404202;
      29455: inst = 32'h8220000;
      29456: inst = 32'h10408000;
      29457: inst = 32'hc404203;
      29458: inst = 32'h8220000;
      29459: inst = 32'h10408000;
      29460: inst = 32'hc404204;
      29461: inst = 32'h8220000;
      29462: inst = 32'h10408000;
      29463: inst = 32'hc404205;
      29464: inst = 32'h8220000;
      29465: inst = 32'h10408000;
      29466: inst = 32'hc404206;
      29467: inst = 32'h8220000;
      29468: inst = 32'h10408000;
      29469: inst = 32'hc404207;
      29470: inst = 32'h8220000;
      29471: inst = 32'h10408000;
      29472: inst = 32'hc404208;
      29473: inst = 32'h8220000;
      29474: inst = 32'h10408000;
      29475: inst = 32'hc404209;
      29476: inst = 32'h8220000;
      29477: inst = 32'h10408000;
      29478: inst = 32'hc40420a;
      29479: inst = 32'h8220000;
      29480: inst = 32'h10408000;
      29481: inst = 32'hc40420b;
      29482: inst = 32'h8220000;
      29483: inst = 32'h10408000;
      29484: inst = 32'hc40420f;
      29485: inst = 32'h8220000;
      29486: inst = 32'h10408000;
      29487: inst = 32'hc404214;
      29488: inst = 32'h8220000;
      29489: inst = 32'h10408000;
      29490: inst = 32'hc404223;
      29491: inst = 32'h8220000;
      29492: inst = 32'h10408000;
      29493: inst = 32'hc40422d;
      29494: inst = 32'h8220000;
      29495: inst = 32'h10408000;
      29496: inst = 32'hc40422e;
      29497: inst = 32'h8220000;
      29498: inst = 32'h10408000;
      29499: inst = 32'hc404232;
      29500: inst = 32'h8220000;
      29501: inst = 32'h10408000;
      29502: inst = 32'hc404233;
      29503: inst = 32'h8220000;
      29504: inst = 32'h10408000;
      29505: inst = 32'hc404234;
      29506: inst = 32'h8220000;
      29507: inst = 32'h10408000;
      29508: inst = 32'hc404235;
      29509: inst = 32'h8220000;
      29510: inst = 32'h10408000;
      29511: inst = 32'hc404236;
      29512: inst = 32'h8220000;
      29513: inst = 32'h10408000;
      29514: inst = 32'hc404237;
      29515: inst = 32'h8220000;
      29516: inst = 32'h10408000;
      29517: inst = 32'hc404238;
      29518: inst = 32'h8220000;
      29519: inst = 32'h10408000;
      29520: inst = 32'hc404239;
      29521: inst = 32'h8220000;
      29522: inst = 32'h10408000;
      29523: inst = 32'hc40423a;
      29524: inst = 32'h8220000;
      29525: inst = 32'h10408000;
      29526: inst = 32'hc40423d;
      29527: inst = 32'h8220000;
      29528: inst = 32'h10408000;
      29529: inst = 32'hc40423e;
      29530: inst = 32'h8220000;
      29531: inst = 32'h10408000;
      29532: inst = 32'hc40423f;
      29533: inst = 32'h8220000;
      29534: inst = 32'h10408000;
      29535: inst = 32'hc404240;
      29536: inst = 32'h8220000;
      29537: inst = 32'h10408000;
      29538: inst = 32'hc404241;
      29539: inst = 32'h8220000;
      29540: inst = 32'h10408000;
      29541: inst = 32'hc404242;
      29542: inst = 32'h8220000;
      29543: inst = 32'h10408000;
      29544: inst = 32'hc404243;
      29545: inst = 32'h8220000;
      29546: inst = 32'h10408000;
      29547: inst = 32'hc404244;
      29548: inst = 32'h8220000;
      29549: inst = 32'h10408000;
      29550: inst = 32'hc404245;
      29551: inst = 32'h8220000;
      29552: inst = 32'h10408000;
      29553: inst = 32'hc404246;
      29554: inst = 32'h8220000;
      29555: inst = 32'h10408000;
      29556: inst = 32'hc404247;
      29557: inst = 32'h8220000;
      29558: inst = 32'h10408000;
      29559: inst = 32'hc404248;
      29560: inst = 32'h8220000;
      29561: inst = 32'h10408000;
      29562: inst = 32'hc404249;
      29563: inst = 32'h8220000;
      29564: inst = 32'h10408000;
      29565: inst = 32'hc40424a;
      29566: inst = 32'h8220000;
      29567: inst = 32'h10408000;
      29568: inst = 32'hc40424b;
      29569: inst = 32'h8220000;
      29570: inst = 32'h10408000;
      29571: inst = 32'hc40424c;
      29572: inst = 32'h8220000;
      29573: inst = 32'h10408000;
      29574: inst = 32'hc40424d;
      29575: inst = 32'h8220000;
      29576: inst = 32'h10408000;
      29577: inst = 32'hc40424e;
      29578: inst = 32'h8220000;
      29579: inst = 32'h10408000;
      29580: inst = 32'hc40424f;
      29581: inst = 32'h8220000;
      29582: inst = 32'h10408000;
      29583: inst = 32'hc404250;
      29584: inst = 32'h8220000;
      29585: inst = 32'h10408000;
      29586: inst = 32'hc404251;
      29587: inst = 32'h8220000;
      29588: inst = 32'h10408000;
      29589: inst = 32'hc404252;
      29590: inst = 32'h8220000;
      29591: inst = 32'h10408000;
      29592: inst = 32'hc404253;
      29593: inst = 32'h8220000;
      29594: inst = 32'h10408000;
      29595: inst = 32'hc404254;
      29596: inst = 32'h8220000;
      29597: inst = 32'h10408000;
      29598: inst = 32'hc404255;
      29599: inst = 32'h8220000;
      29600: inst = 32'h10408000;
      29601: inst = 32'hc404256;
      29602: inst = 32'h8220000;
      29603: inst = 32'h10408000;
      29604: inst = 32'hc404257;
      29605: inst = 32'h8220000;
      29606: inst = 32'h10408000;
      29607: inst = 32'hc404258;
      29608: inst = 32'h8220000;
      29609: inst = 32'h10408000;
      29610: inst = 32'hc404259;
      29611: inst = 32'h8220000;
      29612: inst = 32'h10408000;
      29613: inst = 32'hc40425a;
      29614: inst = 32'h8220000;
      29615: inst = 32'h10408000;
      29616: inst = 32'hc40425b;
      29617: inst = 32'h8220000;
      29618: inst = 32'h10408000;
      29619: inst = 32'hc40425c;
      29620: inst = 32'h8220000;
      29621: inst = 32'h10408000;
      29622: inst = 32'hc40425d;
      29623: inst = 32'h8220000;
      29624: inst = 32'h10408000;
      29625: inst = 32'hc40425e;
      29626: inst = 32'h8220000;
      29627: inst = 32'h10408000;
      29628: inst = 32'hc40425f;
      29629: inst = 32'h8220000;
      29630: inst = 32'h10408000;
      29631: inst = 32'hc404260;
      29632: inst = 32'h8220000;
      29633: inst = 32'h10408000;
      29634: inst = 32'hc404261;
      29635: inst = 32'h8220000;
      29636: inst = 32'h10408000;
      29637: inst = 32'hc404262;
      29638: inst = 32'h8220000;
      29639: inst = 32'h10408000;
      29640: inst = 32'hc404263;
      29641: inst = 32'h8220000;
      29642: inst = 32'h10408000;
      29643: inst = 32'hc404264;
      29644: inst = 32'h8220000;
      29645: inst = 32'h10408000;
      29646: inst = 32'hc404265;
      29647: inst = 32'h8220000;
      29648: inst = 32'h10408000;
      29649: inst = 32'hc404266;
      29650: inst = 32'h8220000;
      29651: inst = 32'h10408000;
      29652: inst = 32'hc404267;
      29653: inst = 32'h8220000;
      29654: inst = 32'h10408000;
      29655: inst = 32'hc404268;
      29656: inst = 32'h8220000;
      29657: inst = 32'h10408000;
      29658: inst = 32'hc404269;
      29659: inst = 32'h8220000;
      29660: inst = 32'h10408000;
      29661: inst = 32'hc40426a;
      29662: inst = 32'h8220000;
      29663: inst = 32'h10408000;
      29664: inst = 32'hc40426b;
      29665: inst = 32'h8220000;
      29666: inst = 32'h10408000;
      29667: inst = 32'hc40426f;
      29668: inst = 32'h8220000;
      29669: inst = 32'h10408000;
      29670: inst = 32'hc404283;
      29671: inst = 32'h8220000;
      29672: inst = 32'h10408000;
      29673: inst = 32'hc40428d;
      29674: inst = 32'h8220000;
      29675: inst = 32'h10408000;
      29676: inst = 32'hc40428e;
      29677: inst = 32'h8220000;
      29678: inst = 32'h10408000;
      29679: inst = 32'hc404291;
      29680: inst = 32'h8220000;
      29681: inst = 32'h10408000;
      29682: inst = 32'hc404292;
      29683: inst = 32'h8220000;
      29684: inst = 32'h10408000;
      29685: inst = 32'hc404293;
      29686: inst = 32'h8220000;
      29687: inst = 32'h10408000;
      29688: inst = 32'hc404294;
      29689: inst = 32'h8220000;
      29690: inst = 32'h10408000;
      29691: inst = 32'hc404295;
      29692: inst = 32'h8220000;
      29693: inst = 32'h10408000;
      29694: inst = 32'hc404296;
      29695: inst = 32'h8220000;
      29696: inst = 32'h10408000;
      29697: inst = 32'hc404297;
      29698: inst = 32'h8220000;
      29699: inst = 32'h10408000;
      29700: inst = 32'hc404298;
      29701: inst = 32'h8220000;
      29702: inst = 32'h10408000;
      29703: inst = 32'hc404299;
      29704: inst = 32'h8220000;
      29705: inst = 32'h10408000;
      29706: inst = 32'hc40429a;
      29707: inst = 32'h8220000;
      29708: inst = 32'h10408000;
      29709: inst = 32'hc40429d;
      29710: inst = 32'h8220000;
      29711: inst = 32'h10408000;
      29712: inst = 32'hc40429e;
      29713: inst = 32'h8220000;
      29714: inst = 32'h10408000;
      29715: inst = 32'hc40429f;
      29716: inst = 32'h8220000;
      29717: inst = 32'h10408000;
      29718: inst = 32'hc4042a0;
      29719: inst = 32'h8220000;
      29720: inst = 32'h10408000;
      29721: inst = 32'hc4042a1;
      29722: inst = 32'h8220000;
      29723: inst = 32'h10408000;
      29724: inst = 32'hc4042a2;
      29725: inst = 32'h8220000;
      29726: inst = 32'h10408000;
      29727: inst = 32'hc4042a3;
      29728: inst = 32'h8220000;
      29729: inst = 32'h10408000;
      29730: inst = 32'hc4042a4;
      29731: inst = 32'h8220000;
      29732: inst = 32'h10408000;
      29733: inst = 32'hc4042a5;
      29734: inst = 32'h8220000;
      29735: inst = 32'h10408000;
      29736: inst = 32'hc4042a6;
      29737: inst = 32'h8220000;
      29738: inst = 32'h10408000;
      29739: inst = 32'hc4042a7;
      29740: inst = 32'h8220000;
      29741: inst = 32'h10408000;
      29742: inst = 32'hc4042a8;
      29743: inst = 32'h8220000;
      29744: inst = 32'h10408000;
      29745: inst = 32'hc4042a9;
      29746: inst = 32'h8220000;
      29747: inst = 32'h10408000;
      29748: inst = 32'hc4042aa;
      29749: inst = 32'h8220000;
      29750: inst = 32'h10408000;
      29751: inst = 32'hc4042ab;
      29752: inst = 32'h8220000;
      29753: inst = 32'h10408000;
      29754: inst = 32'hc4042ac;
      29755: inst = 32'h8220000;
      29756: inst = 32'h10408000;
      29757: inst = 32'hc4042ad;
      29758: inst = 32'h8220000;
      29759: inst = 32'h10408000;
      29760: inst = 32'hc4042ae;
      29761: inst = 32'h8220000;
      29762: inst = 32'h10408000;
      29763: inst = 32'hc4042af;
      29764: inst = 32'h8220000;
      29765: inst = 32'h10408000;
      29766: inst = 32'hc4042b0;
      29767: inst = 32'h8220000;
      29768: inst = 32'h10408000;
      29769: inst = 32'hc4042b1;
      29770: inst = 32'h8220000;
      29771: inst = 32'h10408000;
      29772: inst = 32'hc4042b2;
      29773: inst = 32'h8220000;
      29774: inst = 32'h10408000;
      29775: inst = 32'hc4042b3;
      29776: inst = 32'h8220000;
      29777: inst = 32'h10408000;
      29778: inst = 32'hc4042b4;
      29779: inst = 32'h8220000;
      29780: inst = 32'h10408000;
      29781: inst = 32'hc4042b5;
      29782: inst = 32'h8220000;
      29783: inst = 32'h10408000;
      29784: inst = 32'hc4042b6;
      29785: inst = 32'h8220000;
      29786: inst = 32'h10408000;
      29787: inst = 32'hc4042b7;
      29788: inst = 32'h8220000;
      29789: inst = 32'h10408000;
      29790: inst = 32'hc4042b8;
      29791: inst = 32'h8220000;
      29792: inst = 32'h10408000;
      29793: inst = 32'hc4042b9;
      29794: inst = 32'h8220000;
      29795: inst = 32'h10408000;
      29796: inst = 32'hc4042ba;
      29797: inst = 32'h8220000;
      29798: inst = 32'h10408000;
      29799: inst = 32'hc4042bb;
      29800: inst = 32'h8220000;
      29801: inst = 32'h10408000;
      29802: inst = 32'hc4042bc;
      29803: inst = 32'h8220000;
      29804: inst = 32'h10408000;
      29805: inst = 32'hc4042bd;
      29806: inst = 32'h8220000;
      29807: inst = 32'h10408000;
      29808: inst = 32'hc4042be;
      29809: inst = 32'h8220000;
      29810: inst = 32'h10408000;
      29811: inst = 32'hc4042bf;
      29812: inst = 32'h8220000;
      29813: inst = 32'h10408000;
      29814: inst = 32'hc4042c0;
      29815: inst = 32'h8220000;
      29816: inst = 32'h10408000;
      29817: inst = 32'hc4042c1;
      29818: inst = 32'h8220000;
      29819: inst = 32'h10408000;
      29820: inst = 32'hc4042c2;
      29821: inst = 32'h8220000;
      29822: inst = 32'h10408000;
      29823: inst = 32'hc4042c3;
      29824: inst = 32'h8220000;
      29825: inst = 32'h10408000;
      29826: inst = 32'hc4042c4;
      29827: inst = 32'h8220000;
      29828: inst = 32'h10408000;
      29829: inst = 32'hc4042c5;
      29830: inst = 32'h8220000;
      29831: inst = 32'h10408000;
      29832: inst = 32'hc4042c6;
      29833: inst = 32'h8220000;
      29834: inst = 32'h10408000;
      29835: inst = 32'hc4042c7;
      29836: inst = 32'h8220000;
      29837: inst = 32'h10408000;
      29838: inst = 32'hc4042c8;
      29839: inst = 32'h8220000;
      29840: inst = 32'h10408000;
      29841: inst = 32'hc4042c9;
      29842: inst = 32'h8220000;
      29843: inst = 32'h10408000;
      29844: inst = 32'hc4042ca;
      29845: inst = 32'h8220000;
      29846: inst = 32'h10408000;
      29847: inst = 32'hc4042cb;
      29848: inst = 32'h8220000;
      29849: inst = 32'h10408000;
      29850: inst = 32'hc4042cf;
      29851: inst = 32'h8220000;
      29852: inst = 32'h10408000;
      29853: inst = 32'hc4042d3;
      29854: inst = 32'h8220000;
      29855: inst = 32'h10408000;
      29856: inst = 32'hc4042da;
      29857: inst = 32'h8220000;
      29858: inst = 32'h10408000;
      29859: inst = 32'hc4042db;
      29860: inst = 32'h8220000;
      29861: inst = 32'h10408000;
      29862: inst = 32'hc4042e3;
      29863: inst = 32'h8220000;
      29864: inst = 32'h10408000;
      29865: inst = 32'hc4042ed;
      29866: inst = 32'h8220000;
      29867: inst = 32'h10408000;
      29868: inst = 32'hc4042ee;
      29869: inst = 32'h8220000;
      29870: inst = 32'h10408000;
      29871: inst = 32'hc4042ef;
      29872: inst = 32'h8220000;
      29873: inst = 32'h10408000;
      29874: inst = 32'hc4042f0;
      29875: inst = 32'h8220000;
      29876: inst = 32'h10408000;
      29877: inst = 32'hc4042f1;
      29878: inst = 32'h8220000;
      29879: inst = 32'h10408000;
      29880: inst = 32'hc4042f2;
      29881: inst = 32'h8220000;
      29882: inst = 32'h10408000;
      29883: inst = 32'hc4042f3;
      29884: inst = 32'h8220000;
      29885: inst = 32'h10408000;
      29886: inst = 32'hc4042f4;
      29887: inst = 32'h8220000;
      29888: inst = 32'h10408000;
      29889: inst = 32'hc4042f5;
      29890: inst = 32'h8220000;
      29891: inst = 32'h10408000;
      29892: inst = 32'hc4042f6;
      29893: inst = 32'h8220000;
      29894: inst = 32'h10408000;
      29895: inst = 32'hc4042f7;
      29896: inst = 32'h8220000;
      29897: inst = 32'h10408000;
      29898: inst = 32'hc4042f8;
      29899: inst = 32'h8220000;
      29900: inst = 32'h10408000;
      29901: inst = 32'hc4042f9;
      29902: inst = 32'h8220000;
      29903: inst = 32'h10408000;
      29904: inst = 32'hc4042fa;
      29905: inst = 32'h8220000;
      29906: inst = 32'h10408000;
      29907: inst = 32'hc4042fb;
      29908: inst = 32'h8220000;
      29909: inst = 32'h10408000;
      29910: inst = 32'hc4042fc;
      29911: inst = 32'h8220000;
      29912: inst = 32'h10408000;
      29913: inst = 32'hc4042fd;
      29914: inst = 32'h8220000;
      29915: inst = 32'h10408000;
      29916: inst = 32'hc4042fe;
      29917: inst = 32'h8220000;
      29918: inst = 32'h10408000;
      29919: inst = 32'hc4042ff;
      29920: inst = 32'h8220000;
      29921: inst = 32'h10408000;
      29922: inst = 32'hc404300;
      29923: inst = 32'h8220000;
      29924: inst = 32'h10408000;
      29925: inst = 32'hc404301;
      29926: inst = 32'h8220000;
      29927: inst = 32'h10408000;
      29928: inst = 32'hc404302;
      29929: inst = 32'h8220000;
      29930: inst = 32'h10408000;
      29931: inst = 32'hc404303;
      29932: inst = 32'h8220000;
      29933: inst = 32'h10408000;
      29934: inst = 32'hc404304;
      29935: inst = 32'h8220000;
      29936: inst = 32'h10408000;
      29937: inst = 32'hc404305;
      29938: inst = 32'h8220000;
      29939: inst = 32'h10408000;
      29940: inst = 32'hc404306;
      29941: inst = 32'h8220000;
      29942: inst = 32'h10408000;
      29943: inst = 32'hc404307;
      29944: inst = 32'h8220000;
      29945: inst = 32'h10408000;
      29946: inst = 32'hc404308;
      29947: inst = 32'h8220000;
      29948: inst = 32'h10408000;
      29949: inst = 32'hc404309;
      29950: inst = 32'h8220000;
      29951: inst = 32'h10408000;
      29952: inst = 32'hc40430a;
      29953: inst = 32'h8220000;
      29954: inst = 32'h10408000;
      29955: inst = 32'hc40430b;
      29956: inst = 32'h8220000;
      29957: inst = 32'h10408000;
      29958: inst = 32'hc40430c;
      29959: inst = 32'h8220000;
      29960: inst = 32'h10408000;
      29961: inst = 32'hc40430d;
      29962: inst = 32'h8220000;
      29963: inst = 32'h10408000;
      29964: inst = 32'hc40430e;
      29965: inst = 32'h8220000;
      29966: inst = 32'h10408000;
      29967: inst = 32'hc40430f;
      29968: inst = 32'h8220000;
      29969: inst = 32'h10408000;
      29970: inst = 32'hc404310;
      29971: inst = 32'h8220000;
      29972: inst = 32'h10408000;
      29973: inst = 32'hc404311;
      29974: inst = 32'h8220000;
      29975: inst = 32'h10408000;
      29976: inst = 32'hc404312;
      29977: inst = 32'h8220000;
      29978: inst = 32'h10408000;
      29979: inst = 32'hc404313;
      29980: inst = 32'h8220000;
      29981: inst = 32'h10408000;
      29982: inst = 32'hc404314;
      29983: inst = 32'h8220000;
      29984: inst = 32'h10408000;
      29985: inst = 32'hc404315;
      29986: inst = 32'h8220000;
      29987: inst = 32'h10408000;
      29988: inst = 32'hc404316;
      29989: inst = 32'h8220000;
      29990: inst = 32'h10408000;
      29991: inst = 32'hc404317;
      29992: inst = 32'h8220000;
      29993: inst = 32'h10408000;
      29994: inst = 32'hc404318;
      29995: inst = 32'h8220000;
      29996: inst = 32'h10408000;
      29997: inst = 32'hc404319;
      29998: inst = 32'h8220000;
      29999: inst = 32'h10408000;
      30000: inst = 32'hc40431a;
      30001: inst = 32'h8220000;
      30002: inst = 32'h10408000;
      30003: inst = 32'hc40431b;
      30004: inst = 32'h8220000;
      30005: inst = 32'h10408000;
      30006: inst = 32'hc40431c;
      30007: inst = 32'h8220000;
      30008: inst = 32'h10408000;
      30009: inst = 32'hc40431d;
      30010: inst = 32'h8220000;
      30011: inst = 32'h10408000;
      30012: inst = 32'hc40431e;
      30013: inst = 32'h8220000;
      30014: inst = 32'h10408000;
      30015: inst = 32'hc40431f;
      30016: inst = 32'h8220000;
      30017: inst = 32'h10408000;
      30018: inst = 32'hc404320;
      30019: inst = 32'h8220000;
      30020: inst = 32'h10408000;
      30021: inst = 32'hc404321;
      30022: inst = 32'h8220000;
      30023: inst = 32'h10408000;
      30024: inst = 32'hc404322;
      30025: inst = 32'h8220000;
      30026: inst = 32'h10408000;
      30027: inst = 32'hc404323;
      30028: inst = 32'h8220000;
      30029: inst = 32'h10408000;
      30030: inst = 32'hc404324;
      30031: inst = 32'h8220000;
      30032: inst = 32'h10408000;
      30033: inst = 32'hc404325;
      30034: inst = 32'h8220000;
      30035: inst = 32'h10408000;
      30036: inst = 32'hc404326;
      30037: inst = 32'h8220000;
      30038: inst = 32'h10408000;
      30039: inst = 32'hc404327;
      30040: inst = 32'h8220000;
      30041: inst = 32'h10408000;
      30042: inst = 32'hc404328;
      30043: inst = 32'h8220000;
      30044: inst = 32'h10408000;
      30045: inst = 32'hc404329;
      30046: inst = 32'h8220000;
      30047: inst = 32'h10408000;
      30048: inst = 32'hc40432a;
      30049: inst = 32'h8220000;
      30050: inst = 32'h10408000;
      30051: inst = 32'hc40432b;
      30052: inst = 32'h8220000;
      30053: inst = 32'h10408000;
      30054: inst = 32'hc40432f;
      30055: inst = 32'h8220000;
      30056: inst = 32'h10408000;
      30057: inst = 32'hc404330;
      30058: inst = 32'h8220000;
      30059: inst = 32'h10408000;
      30060: inst = 32'hc404333;
      30061: inst = 32'h8220000;
      30062: inst = 32'h10408000;
      30063: inst = 32'hc404334;
      30064: inst = 32'h8220000;
      30065: inst = 32'h10408000;
      30066: inst = 32'hc404343;
      30067: inst = 32'h8220000;
      30068: inst = 32'h10408000;
      30069: inst = 32'hc40434d;
      30070: inst = 32'h8220000;
      30071: inst = 32'h10408000;
      30072: inst = 32'hc40434e;
      30073: inst = 32'h8220000;
      30074: inst = 32'h10408000;
      30075: inst = 32'hc40434f;
      30076: inst = 32'h8220000;
      30077: inst = 32'h10408000;
      30078: inst = 32'hc404350;
      30079: inst = 32'h8220000;
      30080: inst = 32'h10408000;
      30081: inst = 32'hc404351;
      30082: inst = 32'h8220000;
      30083: inst = 32'h10408000;
      30084: inst = 32'hc404352;
      30085: inst = 32'h8220000;
      30086: inst = 32'h10408000;
      30087: inst = 32'hc404353;
      30088: inst = 32'h8220000;
      30089: inst = 32'h10408000;
      30090: inst = 32'hc404354;
      30091: inst = 32'h8220000;
      30092: inst = 32'h10408000;
      30093: inst = 32'hc404355;
      30094: inst = 32'h8220000;
      30095: inst = 32'h10408000;
      30096: inst = 32'hc404356;
      30097: inst = 32'h8220000;
      30098: inst = 32'h10408000;
      30099: inst = 32'hc404357;
      30100: inst = 32'h8220000;
      30101: inst = 32'h10408000;
      30102: inst = 32'hc404358;
      30103: inst = 32'h8220000;
      30104: inst = 32'h10408000;
      30105: inst = 32'hc404359;
      30106: inst = 32'h8220000;
      30107: inst = 32'h10408000;
      30108: inst = 32'hc40435a;
      30109: inst = 32'h8220000;
      30110: inst = 32'h10408000;
      30111: inst = 32'hc40435b;
      30112: inst = 32'h8220000;
      30113: inst = 32'h10408000;
      30114: inst = 32'hc40435c;
      30115: inst = 32'h8220000;
      30116: inst = 32'h10408000;
      30117: inst = 32'hc40435d;
      30118: inst = 32'h8220000;
      30119: inst = 32'h10408000;
      30120: inst = 32'hc40435e;
      30121: inst = 32'h8220000;
      30122: inst = 32'h10408000;
      30123: inst = 32'hc40435f;
      30124: inst = 32'h8220000;
      30125: inst = 32'h10408000;
      30126: inst = 32'hc404360;
      30127: inst = 32'h8220000;
      30128: inst = 32'h10408000;
      30129: inst = 32'hc404361;
      30130: inst = 32'h8220000;
      30131: inst = 32'h10408000;
      30132: inst = 32'hc404362;
      30133: inst = 32'h8220000;
      30134: inst = 32'h10408000;
      30135: inst = 32'hc404363;
      30136: inst = 32'h8220000;
      30137: inst = 32'h10408000;
      30138: inst = 32'hc404364;
      30139: inst = 32'h8220000;
      30140: inst = 32'h10408000;
      30141: inst = 32'hc404365;
      30142: inst = 32'h8220000;
      30143: inst = 32'h10408000;
      30144: inst = 32'hc404366;
      30145: inst = 32'h8220000;
      30146: inst = 32'h10408000;
      30147: inst = 32'hc404367;
      30148: inst = 32'h8220000;
      30149: inst = 32'h10408000;
      30150: inst = 32'hc404368;
      30151: inst = 32'h8220000;
      30152: inst = 32'h10408000;
      30153: inst = 32'hc404369;
      30154: inst = 32'h8220000;
      30155: inst = 32'h10408000;
      30156: inst = 32'hc40436a;
      30157: inst = 32'h8220000;
      30158: inst = 32'h10408000;
      30159: inst = 32'hc40436b;
      30160: inst = 32'h8220000;
      30161: inst = 32'h10408000;
      30162: inst = 32'hc40436c;
      30163: inst = 32'h8220000;
      30164: inst = 32'h10408000;
      30165: inst = 32'hc40436d;
      30166: inst = 32'h8220000;
      30167: inst = 32'h10408000;
      30168: inst = 32'hc40436e;
      30169: inst = 32'h8220000;
      30170: inst = 32'h10408000;
      30171: inst = 32'hc40436f;
      30172: inst = 32'h8220000;
      30173: inst = 32'h10408000;
      30174: inst = 32'hc404370;
      30175: inst = 32'h8220000;
      30176: inst = 32'h10408000;
      30177: inst = 32'hc404371;
      30178: inst = 32'h8220000;
      30179: inst = 32'h10408000;
      30180: inst = 32'hc404372;
      30181: inst = 32'h8220000;
      30182: inst = 32'h10408000;
      30183: inst = 32'hc404373;
      30184: inst = 32'h8220000;
      30185: inst = 32'h10408000;
      30186: inst = 32'hc404374;
      30187: inst = 32'h8220000;
      30188: inst = 32'h10408000;
      30189: inst = 32'hc404375;
      30190: inst = 32'h8220000;
      30191: inst = 32'h10408000;
      30192: inst = 32'hc404376;
      30193: inst = 32'h8220000;
      30194: inst = 32'h10408000;
      30195: inst = 32'hc404377;
      30196: inst = 32'h8220000;
      30197: inst = 32'h10408000;
      30198: inst = 32'hc404378;
      30199: inst = 32'h8220000;
      30200: inst = 32'h10408000;
      30201: inst = 32'hc404379;
      30202: inst = 32'h8220000;
      30203: inst = 32'h10408000;
      30204: inst = 32'hc40437a;
      30205: inst = 32'h8220000;
      30206: inst = 32'h10408000;
      30207: inst = 32'hc40437b;
      30208: inst = 32'h8220000;
      30209: inst = 32'h10408000;
      30210: inst = 32'hc40437c;
      30211: inst = 32'h8220000;
      30212: inst = 32'h10408000;
      30213: inst = 32'hc40437d;
      30214: inst = 32'h8220000;
      30215: inst = 32'h10408000;
      30216: inst = 32'hc40437e;
      30217: inst = 32'h8220000;
      30218: inst = 32'h10408000;
      30219: inst = 32'hc40437f;
      30220: inst = 32'h8220000;
      30221: inst = 32'h10408000;
      30222: inst = 32'hc404380;
      30223: inst = 32'h8220000;
      30224: inst = 32'h10408000;
      30225: inst = 32'hc404381;
      30226: inst = 32'h8220000;
      30227: inst = 32'h10408000;
      30228: inst = 32'hc404382;
      30229: inst = 32'h8220000;
      30230: inst = 32'h10408000;
      30231: inst = 32'hc404383;
      30232: inst = 32'h8220000;
      30233: inst = 32'h10408000;
      30234: inst = 32'hc404384;
      30235: inst = 32'h8220000;
      30236: inst = 32'h10408000;
      30237: inst = 32'hc404385;
      30238: inst = 32'h8220000;
      30239: inst = 32'h10408000;
      30240: inst = 32'hc404386;
      30241: inst = 32'h8220000;
      30242: inst = 32'h10408000;
      30243: inst = 32'hc404387;
      30244: inst = 32'h8220000;
      30245: inst = 32'h10408000;
      30246: inst = 32'hc404388;
      30247: inst = 32'h8220000;
      30248: inst = 32'h10408000;
      30249: inst = 32'hc404389;
      30250: inst = 32'h8220000;
      30251: inst = 32'h10408000;
      30252: inst = 32'hc40438a;
      30253: inst = 32'h8220000;
      30254: inst = 32'h10408000;
      30255: inst = 32'hc40438b;
      30256: inst = 32'h8220000;
      30257: inst = 32'h10408000;
      30258: inst = 32'hc40438f;
      30259: inst = 32'h8220000;
      30260: inst = 32'h10408000;
      30261: inst = 32'hc404390;
      30262: inst = 32'h8220000;
      30263: inst = 32'h10408000;
      30264: inst = 32'hc4043a3;
      30265: inst = 32'h8220000;
      30266: inst = 32'h10408000;
      30267: inst = 32'hc4043ad;
      30268: inst = 32'h8220000;
      30269: inst = 32'h10408000;
      30270: inst = 32'hc4043ae;
      30271: inst = 32'h8220000;
      30272: inst = 32'h10408000;
      30273: inst = 32'hc4043af;
      30274: inst = 32'h8220000;
      30275: inst = 32'h10408000;
      30276: inst = 32'hc4043b0;
      30277: inst = 32'h8220000;
      30278: inst = 32'h10408000;
      30279: inst = 32'hc4043b1;
      30280: inst = 32'h8220000;
      30281: inst = 32'h10408000;
      30282: inst = 32'hc4043b2;
      30283: inst = 32'h8220000;
      30284: inst = 32'h10408000;
      30285: inst = 32'hc4043b3;
      30286: inst = 32'h8220000;
      30287: inst = 32'h10408000;
      30288: inst = 32'hc4043b4;
      30289: inst = 32'h8220000;
      30290: inst = 32'h10408000;
      30291: inst = 32'hc4043b5;
      30292: inst = 32'h8220000;
      30293: inst = 32'h10408000;
      30294: inst = 32'hc4043b6;
      30295: inst = 32'h8220000;
      30296: inst = 32'h10408000;
      30297: inst = 32'hc4043b7;
      30298: inst = 32'h8220000;
      30299: inst = 32'h10408000;
      30300: inst = 32'hc4043b8;
      30301: inst = 32'h8220000;
      30302: inst = 32'h10408000;
      30303: inst = 32'hc4043b9;
      30304: inst = 32'h8220000;
      30305: inst = 32'h10408000;
      30306: inst = 32'hc4043ba;
      30307: inst = 32'h8220000;
      30308: inst = 32'h10408000;
      30309: inst = 32'hc4043bb;
      30310: inst = 32'h8220000;
      30311: inst = 32'h10408000;
      30312: inst = 32'hc4043bc;
      30313: inst = 32'h8220000;
      30314: inst = 32'h10408000;
      30315: inst = 32'hc4043bd;
      30316: inst = 32'h8220000;
      30317: inst = 32'h10408000;
      30318: inst = 32'hc4043be;
      30319: inst = 32'h8220000;
      30320: inst = 32'h10408000;
      30321: inst = 32'hc4043bf;
      30322: inst = 32'h8220000;
      30323: inst = 32'h10408000;
      30324: inst = 32'hc4043c0;
      30325: inst = 32'h8220000;
      30326: inst = 32'h10408000;
      30327: inst = 32'hc4043c1;
      30328: inst = 32'h8220000;
      30329: inst = 32'h10408000;
      30330: inst = 32'hc4043c2;
      30331: inst = 32'h8220000;
      30332: inst = 32'h10408000;
      30333: inst = 32'hc4043c3;
      30334: inst = 32'h8220000;
      30335: inst = 32'h10408000;
      30336: inst = 32'hc4043c4;
      30337: inst = 32'h8220000;
      30338: inst = 32'h10408000;
      30339: inst = 32'hc4043c5;
      30340: inst = 32'h8220000;
      30341: inst = 32'h10408000;
      30342: inst = 32'hc4043c6;
      30343: inst = 32'h8220000;
      30344: inst = 32'h10408000;
      30345: inst = 32'hc4043c7;
      30346: inst = 32'h8220000;
      30347: inst = 32'h10408000;
      30348: inst = 32'hc4043c8;
      30349: inst = 32'h8220000;
      30350: inst = 32'h10408000;
      30351: inst = 32'hc4043c9;
      30352: inst = 32'h8220000;
      30353: inst = 32'h10408000;
      30354: inst = 32'hc4043ca;
      30355: inst = 32'h8220000;
      30356: inst = 32'h10408000;
      30357: inst = 32'hc4043cb;
      30358: inst = 32'h8220000;
      30359: inst = 32'h10408000;
      30360: inst = 32'hc4043cc;
      30361: inst = 32'h8220000;
      30362: inst = 32'h10408000;
      30363: inst = 32'hc4043cd;
      30364: inst = 32'h8220000;
      30365: inst = 32'h10408000;
      30366: inst = 32'hc4043ce;
      30367: inst = 32'h8220000;
      30368: inst = 32'h10408000;
      30369: inst = 32'hc4043cf;
      30370: inst = 32'h8220000;
      30371: inst = 32'h10408000;
      30372: inst = 32'hc4043d0;
      30373: inst = 32'h8220000;
      30374: inst = 32'h10408000;
      30375: inst = 32'hc4043d1;
      30376: inst = 32'h8220000;
      30377: inst = 32'h10408000;
      30378: inst = 32'hc4043d2;
      30379: inst = 32'h8220000;
      30380: inst = 32'h10408000;
      30381: inst = 32'hc4043d3;
      30382: inst = 32'h8220000;
      30383: inst = 32'h10408000;
      30384: inst = 32'hc4043d4;
      30385: inst = 32'h8220000;
      30386: inst = 32'h10408000;
      30387: inst = 32'hc4043d5;
      30388: inst = 32'h8220000;
      30389: inst = 32'h10408000;
      30390: inst = 32'hc4043d6;
      30391: inst = 32'h8220000;
      30392: inst = 32'h10408000;
      30393: inst = 32'hc4043d7;
      30394: inst = 32'h8220000;
      30395: inst = 32'h10408000;
      30396: inst = 32'hc4043d8;
      30397: inst = 32'h8220000;
      30398: inst = 32'h10408000;
      30399: inst = 32'hc4043d9;
      30400: inst = 32'h8220000;
      30401: inst = 32'h10408000;
      30402: inst = 32'hc4043da;
      30403: inst = 32'h8220000;
      30404: inst = 32'h10408000;
      30405: inst = 32'hc4043db;
      30406: inst = 32'h8220000;
      30407: inst = 32'h10408000;
      30408: inst = 32'hc4043dc;
      30409: inst = 32'h8220000;
      30410: inst = 32'h10408000;
      30411: inst = 32'hc4043dd;
      30412: inst = 32'h8220000;
      30413: inst = 32'h10408000;
      30414: inst = 32'hc4043de;
      30415: inst = 32'h8220000;
      30416: inst = 32'h10408000;
      30417: inst = 32'hc4043df;
      30418: inst = 32'h8220000;
      30419: inst = 32'h10408000;
      30420: inst = 32'hc4043e0;
      30421: inst = 32'h8220000;
      30422: inst = 32'h10408000;
      30423: inst = 32'hc4043e1;
      30424: inst = 32'h8220000;
      30425: inst = 32'h10408000;
      30426: inst = 32'hc4043e2;
      30427: inst = 32'h8220000;
      30428: inst = 32'h10408000;
      30429: inst = 32'hc4043e3;
      30430: inst = 32'h8220000;
      30431: inst = 32'h10408000;
      30432: inst = 32'hc4043e4;
      30433: inst = 32'h8220000;
      30434: inst = 32'h10408000;
      30435: inst = 32'hc4043e5;
      30436: inst = 32'h8220000;
      30437: inst = 32'h10408000;
      30438: inst = 32'hc4043e6;
      30439: inst = 32'h8220000;
      30440: inst = 32'h10408000;
      30441: inst = 32'hc4043e7;
      30442: inst = 32'h8220000;
      30443: inst = 32'h10408000;
      30444: inst = 32'hc4043e8;
      30445: inst = 32'h8220000;
      30446: inst = 32'h10408000;
      30447: inst = 32'hc4043e9;
      30448: inst = 32'h8220000;
      30449: inst = 32'h10408000;
      30450: inst = 32'hc4043ea;
      30451: inst = 32'h8220000;
      30452: inst = 32'h10408000;
      30453: inst = 32'hc4043eb;
      30454: inst = 32'h8220000;
      30455: inst = 32'h10408000;
      30456: inst = 32'hc4043ef;
      30457: inst = 32'h8220000;
      30458: inst = 32'h10408000;
      30459: inst = 32'hc4043f9;
      30460: inst = 32'h8220000;
      30461: inst = 32'h10408000;
      30462: inst = 32'hc404403;
      30463: inst = 32'h8220000;
      30464: inst = 32'h10408000;
      30465: inst = 32'hc404404;
      30466: inst = 32'h8220000;
      30467: inst = 32'h10408000;
      30468: inst = 32'hc404405;
      30469: inst = 32'h8220000;
      30470: inst = 32'h10408000;
      30471: inst = 32'hc404406;
      30472: inst = 32'h8220000;
      30473: inst = 32'h10408000;
      30474: inst = 32'hc404407;
      30475: inst = 32'h8220000;
      30476: inst = 32'h10408000;
      30477: inst = 32'hc404408;
      30478: inst = 32'h8220000;
      30479: inst = 32'h10408000;
      30480: inst = 32'hc404409;
      30481: inst = 32'h8220000;
      30482: inst = 32'h10408000;
      30483: inst = 32'hc40440a;
      30484: inst = 32'h8220000;
      30485: inst = 32'h10408000;
      30486: inst = 32'hc40440b;
      30487: inst = 32'h8220000;
      30488: inst = 32'h10408000;
      30489: inst = 32'hc40440c;
      30490: inst = 32'h8220000;
      30491: inst = 32'h10408000;
      30492: inst = 32'hc40440d;
      30493: inst = 32'h8220000;
      30494: inst = 32'h10408000;
      30495: inst = 32'hc40440e;
      30496: inst = 32'h8220000;
      30497: inst = 32'h10408000;
      30498: inst = 32'hc40440f;
      30499: inst = 32'h8220000;
      30500: inst = 32'h10408000;
      30501: inst = 32'hc404410;
      30502: inst = 32'h8220000;
      30503: inst = 32'h10408000;
      30504: inst = 32'hc404411;
      30505: inst = 32'h8220000;
      30506: inst = 32'h10408000;
      30507: inst = 32'hc404412;
      30508: inst = 32'h8220000;
      30509: inst = 32'h10408000;
      30510: inst = 32'hc404413;
      30511: inst = 32'h8220000;
      30512: inst = 32'h10408000;
      30513: inst = 32'hc404414;
      30514: inst = 32'h8220000;
      30515: inst = 32'h10408000;
      30516: inst = 32'hc404415;
      30517: inst = 32'h8220000;
      30518: inst = 32'h10408000;
      30519: inst = 32'hc404416;
      30520: inst = 32'h8220000;
      30521: inst = 32'h10408000;
      30522: inst = 32'hc404417;
      30523: inst = 32'h8220000;
      30524: inst = 32'h10408000;
      30525: inst = 32'hc404418;
      30526: inst = 32'h8220000;
      30527: inst = 32'h10408000;
      30528: inst = 32'hc404419;
      30529: inst = 32'h8220000;
      30530: inst = 32'h10408000;
      30531: inst = 32'hc40441a;
      30532: inst = 32'h8220000;
      30533: inst = 32'h10408000;
      30534: inst = 32'hc40441b;
      30535: inst = 32'h8220000;
      30536: inst = 32'h10408000;
      30537: inst = 32'hc40441c;
      30538: inst = 32'h8220000;
      30539: inst = 32'h10408000;
      30540: inst = 32'hc40441d;
      30541: inst = 32'h8220000;
      30542: inst = 32'h10408000;
      30543: inst = 32'hc40441e;
      30544: inst = 32'h8220000;
      30545: inst = 32'h10408000;
      30546: inst = 32'hc40441f;
      30547: inst = 32'h8220000;
      30548: inst = 32'h10408000;
      30549: inst = 32'hc404420;
      30550: inst = 32'h8220000;
      30551: inst = 32'h10408000;
      30552: inst = 32'hc404421;
      30553: inst = 32'h8220000;
      30554: inst = 32'h10408000;
      30555: inst = 32'hc404422;
      30556: inst = 32'h8220000;
      30557: inst = 32'h10408000;
      30558: inst = 32'hc404423;
      30559: inst = 32'h8220000;
      30560: inst = 32'h10408000;
      30561: inst = 32'hc404424;
      30562: inst = 32'h8220000;
      30563: inst = 32'h10408000;
      30564: inst = 32'hc404425;
      30565: inst = 32'h8220000;
      30566: inst = 32'h10408000;
      30567: inst = 32'hc404426;
      30568: inst = 32'h8220000;
      30569: inst = 32'h10408000;
      30570: inst = 32'hc404427;
      30571: inst = 32'h8220000;
      30572: inst = 32'h10408000;
      30573: inst = 32'hc404428;
      30574: inst = 32'h8220000;
      30575: inst = 32'h10408000;
      30576: inst = 32'hc404429;
      30577: inst = 32'h8220000;
      30578: inst = 32'h10408000;
      30579: inst = 32'hc40442a;
      30580: inst = 32'h8220000;
      30581: inst = 32'h10408000;
      30582: inst = 32'hc40442b;
      30583: inst = 32'h8220000;
      30584: inst = 32'h10408000;
      30585: inst = 32'hc40442c;
      30586: inst = 32'h8220000;
      30587: inst = 32'h10408000;
      30588: inst = 32'hc40442d;
      30589: inst = 32'h8220000;
      30590: inst = 32'h10408000;
      30591: inst = 32'hc40442e;
      30592: inst = 32'h8220000;
      30593: inst = 32'h10408000;
      30594: inst = 32'hc40442f;
      30595: inst = 32'h8220000;
      30596: inst = 32'h10408000;
      30597: inst = 32'hc404430;
      30598: inst = 32'h8220000;
      30599: inst = 32'h10408000;
      30600: inst = 32'hc404431;
      30601: inst = 32'h8220000;
      30602: inst = 32'h10408000;
      30603: inst = 32'hc404432;
      30604: inst = 32'h8220000;
      30605: inst = 32'h10408000;
      30606: inst = 32'hc404433;
      30607: inst = 32'h8220000;
      30608: inst = 32'h10408000;
      30609: inst = 32'hc404434;
      30610: inst = 32'h8220000;
      30611: inst = 32'h10408000;
      30612: inst = 32'hc404435;
      30613: inst = 32'h8220000;
      30614: inst = 32'h10408000;
      30615: inst = 32'hc404436;
      30616: inst = 32'h8220000;
      30617: inst = 32'h10408000;
      30618: inst = 32'hc404437;
      30619: inst = 32'h8220000;
      30620: inst = 32'h10408000;
      30621: inst = 32'hc404438;
      30622: inst = 32'h8220000;
      30623: inst = 32'h10408000;
      30624: inst = 32'hc404439;
      30625: inst = 32'h8220000;
      30626: inst = 32'h10408000;
      30627: inst = 32'hc40443a;
      30628: inst = 32'h8220000;
      30629: inst = 32'h10408000;
      30630: inst = 32'hc40443b;
      30631: inst = 32'h8220000;
      30632: inst = 32'h10408000;
      30633: inst = 32'hc40443c;
      30634: inst = 32'h8220000;
      30635: inst = 32'h10408000;
      30636: inst = 32'hc40443d;
      30637: inst = 32'h8220000;
      30638: inst = 32'h10408000;
      30639: inst = 32'hc40443e;
      30640: inst = 32'h8220000;
      30641: inst = 32'h10408000;
      30642: inst = 32'hc40443f;
      30643: inst = 32'h8220000;
      30644: inst = 32'h10408000;
      30645: inst = 32'hc404440;
      30646: inst = 32'h8220000;
      30647: inst = 32'h10408000;
      30648: inst = 32'hc404441;
      30649: inst = 32'h8220000;
      30650: inst = 32'h10408000;
      30651: inst = 32'hc404442;
      30652: inst = 32'h8220000;
      30653: inst = 32'h10408000;
      30654: inst = 32'hc404443;
      30655: inst = 32'h8220000;
      30656: inst = 32'h10408000;
      30657: inst = 32'hc404444;
      30658: inst = 32'h8220000;
      30659: inst = 32'h10408000;
      30660: inst = 32'hc404445;
      30661: inst = 32'h8220000;
      30662: inst = 32'h10408000;
      30663: inst = 32'hc404446;
      30664: inst = 32'h8220000;
      30665: inst = 32'h10408000;
      30666: inst = 32'hc404447;
      30667: inst = 32'h8220000;
      30668: inst = 32'h10408000;
      30669: inst = 32'hc404448;
      30670: inst = 32'h8220000;
      30671: inst = 32'h10408000;
      30672: inst = 32'hc404449;
      30673: inst = 32'h8220000;
      30674: inst = 32'h10408000;
      30675: inst = 32'hc40444a;
      30676: inst = 32'h8220000;
      30677: inst = 32'h10408000;
      30678: inst = 32'hc40444b;
      30679: inst = 32'h8220000;
      30680: inst = 32'h10408000;
      30681: inst = 32'hc40444f;
      30682: inst = 32'h8220000;
      30683: inst = 32'h10408000;
      30684: inst = 32'hc404455;
      30685: inst = 32'h8220000;
      30686: inst = 32'h10408000;
      30687: inst = 32'hc404463;
      30688: inst = 32'h8220000;
      30689: inst = 32'h10408000;
      30690: inst = 32'hc404464;
      30691: inst = 32'h8220000;
      30692: inst = 32'h10408000;
      30693: inst = 32'hc404465;
      30694: inst = 32'h8220000;
      30695: inst = 32'h10408000;
      30696: inst = 32'hc404466;
      30697: inst = 32'h8220000;
      30698: inst = 32'h10408000;
      30699: inst = 32'hc404467;
      30700: inst = 32'h8220000;
      30701: inst = 32'h10408000;
      30702: inst = 32'hc404468;
      30703: inst = 32'h8220000;
      30704: inst = 32'h10408000;
      30705: inst = 32'hc404469;
      30706: inst = 32'h8220000;
      30707: inst = 32'h10408000;
      30708: inst = 32'hc40446a;
      30709: inst = 32'h8220000;
      30710: inst = 32'h10408000;
      30711: inst = 32'hc40446b;
      30712: inst = 32'h8220000;
      30713: inst = 32'h10408000;
      30714: inst = 32'hc40446c;
      30715: inst = 32'h8220000;
      30716: inst = 32'h10408000;
      30717: inst = 32'hc40446d;
      30718: inst = 32'h8220000;
      30719: inst = 32'h10408000;
      30720: inst = 32'hc40446e;
      30721: inst = 32'h8220000;
      30722: inst = 32'h10408000;
      30723: inst = 32'hc40446f;
      30724: inst = 32'h8220000;
      30725: inst = 32'h10408000;
      30726: inst = 32'hc404470;
      30727: inst = 32'h8220000;
      30728: inst = 32'h10408000;
      30729: inst = 32'hc404471;
      30730: inst = 32'h8220000;
      30731: inst = 32'h10408000;
      30732: inst = 32'hc404472;
      30733: inst = 32'h8220000;
      30734: inst = 32'h10408000;
      30735: inst = 32'hc404473;
      30736: inst = 32'h8220000;
      30737: inst = 32'h10408000;
      30738: inst = 32'hc404474;
      30739: inst = 32'h8220000;
      30740: inst = 32'h10408000;
      30741: inst = 32'hc404475;
      30742: inst = 32'h8220000;
      30743: inst = 32'h10408000;
      30744: inst = 32'hc404476;
      30745: inst = 32'h8220000;
      30746: inst = 32'h10408000;
      30747: inst = 32'hc404477;
      30748: inst = 32'h8220000;
      30749: inst = 32'h10408000;
      30750: inst = 32'hc404478;
      30751: inst = 32'h8220000;
      30752: inst = 32'h10408000;
      30753: inst = 32'hc404479;
      30754: inst = 32'h8220000;
      30755: inst = 32'h10408000;
      30756: inst = 32'hc40447a;
      30757: inst = 32'h8220000;
      30758: inst = 32'h10408000;
      30759: inst = 32'hc40447b;
      30760: inst = 32'h8220000;
      30761: inst = 32'h10408000;
      30762: inst = 32'hc40447c;
      30763: inst = 32'h8220000;
      30764: inst = 32'h10408000;
      30765: inst = 32'hc40447d;
      30766: inst = 32'h8220000;
      30767: inst = 32'h10408000;
      30768: inst = 32'hc40447e;
      30769: inst = 32'h8220000;
      30770: inst = 32'h10408000;
      30771: inst = 32'hc40447f;
      30772: inst = 32'h8220000;
      30773: inst = 32'h10408000;
      30774: inst = 32'hc404480;
      30775: inst = 32'h8220000;
      30776: inst = 32'h10408000;
      30777: inst = 32'hc404481;
      30778: inst = 32'h8220000;
      30779: inst = 32'h10408000;
      30780: inst = 32'hc404482;
      30781: inst = 32'h8220000;
      30782: inst = 32'h10408000;
      30783: inst = 32'hc404483;
      30784: inst = 32'h8220000;
      30785: inst = 32'h10408000;
      30786: inst = 32'hc404484;
      30787: inst = 32'h8220000;
      30788: inst = 32'h10408000;
      30789: inst = 32'hc404485;
      30790: inst = 32'h8220000;
      30791: inst = 32'h10408000;
      30792: inst = 32'hc404486;
      30793: inst = 32'h8220000;
      30794: inst = 32'h10408000;
      30795: inst = 32'hc404487;
      30796: inst = 32'h8220000;
      30797: inst = 32'h10408000;
      30798: inst = 32'hc404488;
      30799: inst = 32'h8220000;
      30800: inst = 32'h10408000;
      30801: inst = 32'hc404489;
      30802: inst = 32'h8220000;
      30803: inst = 32'h10408000;
      30804: inst = 32'hc40448a;
      30805: inst = 32'h8220000;
      30806: inst = 32'h10408000;
      30807: inst = 32'hc40448b;
      30808: inst = 32'h8220000;
      30809: inst = 32'h10408000;
      30810: inst = 32'hc40448c;
      30811: inst = 32'h8220000;
      30812: inst = 32'h10408000;
      30813: inst = 32'hc40448d;
      30814: inst = 32'h8220000;
      30815: inst = 32'h10408000;
      30816: inst = 32'hc40448e;
      30817: inst = 32'h8220000;
      30818: inst = 32'h10408000;
      30819: inst = 32'hc40448f;
      30820: inst = 32'h8220000;
      30821: inst = 32'h10408000;
      30822: inst = 32'hc404490;
      30823: inst = 32'h8220000;
      30824: inst = 32'h10408000;
      30825: inst = 32'hc404491;
      30826: inst = 32'h8220000;
      30827: inst = 32'h10408000;
      30828: inst = 32'hc404492;
      30829: inst = 32'h8220000;
      30830: inst = 32'h10408000;
      30831: inst = 32'hc404493;
      30832: inst = 32'h8220000;
      30833: inst = 32'h10408000;
      30834: inst = 32'hc404494;
      30835: inst = 32'h8220000;
      30836: inst = 32'h10408000;
      30837: inst = 32'hc404495;
      30838: inst = 32'h8220000;
      30839: inst = 32'h10408000;
      30840: inst = 32'hc404496;
      30841: inst = 32'h8220000;
      30842: inst = 32'h10408000;
      30843: inst = 32'hc404497;
      30844: inst = 32'h8220000;
      30845: inst = 32'h10408000;
      30846: inst = 32'hc404498;
      30847: inst = 32'h8220000;
      30848: inst = 32'h10408000;
      30849: inst = 32'hc404499;
      30850: inst = 32'h8220000;
      30851: inst = 32'h10408000;
      30852: inst = 32'hc40449a;
      30853: inst = 32'h8220000;
      30854: inst = 32'h10408000;
      30855: inst = 32'hc40449b;
      30856: inst = 32'h8220000;
      30857: inst = 32'h10408000;
      30858: inst = 32'hc40449c;
      30859: inst = 32'h8220000;
      30860: inst = 32'h10408000;
      30861: inst = 32'hc40449d;
      30862: inst = 32'h8220000;
      30863: inst = 32'h10408000;
      30864: inst = 32'hc40449e;
      30865: inst = 32'h8220000;
      30866: inst = 32'h10408000;
      30867: inst = 32'hc40449f;
      30868: inst = 32'h8220000;
      30869: inst = 32'h10408000;
      30870: inst = 32'hc4044a0;
      30871: inst = 32'h8220000;
      30872: inst = 32'h10408000;
      30873: inst = 32'hc4044a1;
      30874: inst = 32'h8220000;
      30875: inst = 32'h10408000;
      30876: inst = 32'hc4044a2;
      30877: inst = 32'h8220000;
      30878: inst = 32'h10408000;
      30879: inst = 32'hc4044a3;
      30880: inst = 32'h8220000;
      30881: inst = 32'h10408000;
      30882: inst = 32'hc4044a4;
      30883: inst = 32'h8220000;
      30884: inst = 32'h10408000;
      30885: inst = 32'hc4044a5;
      30886: inst = 32'h8220000;
      30887: inst = 32'h10408000;
      30888: inst = 32'hc4044a6;
      30889: inst = 32'h8220000;
      30890: inst = 32'h10408000;
      30891: inst = 32'hc4044a7;
      30892: inst = 32'h8220000;
      30893: inst = 32'h10408000;
      30894: inst = 32'hc4044a8;
      30895: inst = 32'h8220000;
      30896: inst = 32'h10408000;
      30897: inst = 32'hc4044a9;
      30898: inst = 32'h8220000;
      30899: inst = 32'h10408000;
      30900: inst = 32'hc4044aa;
      30901: inst = 32'h8220000;
      30902: inst = 32'h10408000;
      30903: inst = 32'hc4044ab;
      30904: inst = 32'h8220000;
      30905: inst = 32'h10408000;
      30906: inst = 32'hc4044af;
      30907: inst = 32'h8220000;
      30908: inst = 32'h10408000;
      30909: inst = 32'hc4044b0;
      30910: inst = 32'h8220000;
      30911: inst = 32'h10408000;
      30912: inst = 32'hc4044b1;
      30913: inst = 32'h8220000;
      30914: inst = 32'h10408000;
      30915: inst = 32'hc4044b2;
      30916: inst = 32'h8220000;
      30917: inst = 32'h10408000;
      30918: inst = 32'hc4044b7;
      30919: inst = 32'h8220000;
      30920: inst = 32'h10408000;
      30921: inst = 32'hc4044c3;
      30922: inst = 32'h8220000;
      30923: inst = 32'h10408000;
      30924: inst = 32'hc4044c4;
      30925: inst = 32'h8220000;
      30926: inst = 32'h10408000;
      30927: inst = 32'hc4044c5;
      30928: inst = 32'h8220000;
      30929: inst = 32'h10408000;
      30930: inst = 32'hc4044c6;
      30931: inst = 32'h8220000;
      30932: inst = 32'h10408000;
      30933: inst = 32'hc4044c7;
      30934: inst = 32'h8220000;
      30935: inst = 32'h10408000;
      30936: inst = 32'hc4044c8;
      30937: inst = 32'h8220000;
      30938: inst = 32'h10408000;
      30939: inst = 32'hc4044c9;
      30940: inst = 32'h8220000;
      30941: inst = 32'h10408000;
      30942: inst = 32'hc4044ca;
      30943: inst = 32'h8220000;
      30944: inst = 32'h10408000;
      30945: inst = 32'hc4044cb;
      30946: inst = 32'h8220000;
      30947: inst = 32'h10408000;
      30948: inst = 32'hc4044cc;
      30949: inst = 32'h8220000;
      30950: inst = 32'h10408000;
      30951: inst = 32'hc4044cd;
      30952: inst = 32'h8220000;
      30953: inst = 32'h10408000;
      30954: inst = 32'hc4044ce;
      30955: inst = 32'h8220000;
      30956: inst = 32'h10408000;
      30957: inst = 32'hc4044cf;
      30958: inst = 32'h8220000;
      30959: inst = 32'h10408000;
      30960: inst = 32'hc4044d0;
      30961: inst = 32'h8220000;
      30962: inst = 32'h10408000;
      30963: inst = 32'hc4044d1;
      30964: inst = 32'h8220000;
      30965: inst = 32'h10408000;
      30966: inst = 32'hc4044d2;
      30967: inst = 32'h8220000;
      30968: inst = 32'h10408000;
      30969: inst = 32'hc4044d3;
      30970: inst = 32'h8220000;
      30971: inst = 32'h10408000;
      30972: inst = 32'hc4044d4;
      30973: inst = 32'h8220000;
      30974: inst = 32'h10408000;
      30975: inst = 32'hc4044d5;
      30976: inst = 32'h8220000;
      30977: inst = 32'h10408000;
      30978: inst = 32'hc4044d6;
      30979: inst = 32'h8220000;
      30980: inst = 32'h10408000;
      30981: inst = 32'hc4044d7;
      30982: inst = 32'h8220000;
      30983: inst = 32'h10408000;
      30984: inst = 32'hc4044d8;
      30985: inst = 32'h8220000;
      30986: inst = 32'h10408000;
      30987: inst = 32'hc4044d9;
      30988: inst = 32'h8220000;
      30989: inst = 32'h10408000;
      30990: inst = 32'hc4044da;
      30991: inst = 32'h8220000;
      30992: inst = 32'h10408000;
      30993: inst = 32'hc4044db;
      30994: inst = 32'h8220000;
      30995: inst = 32'h10408000;
      30996: inst = 32'hc4044dc;
      30997: inst = 32'h8220000;
      30998: inst = 32'h10408000;
      30999: inst = 32'hc4044dd;
      31000: inst = 32'h8220000;
      31001: inst = 32'h10408000;
      31002: inst = 32'hc4044de;
      31003: inst = 32'h8220000;
      31004: inst = 32'h10408000;
      31005: inst = 32'hc4044df;
      31006: inst = 32'h8220000;
      31007: inst = 32'h10408000;
      31008: inst = 32'hc4044e0;
      31009: inst = 32'h8220000;
      31010: inst = 32'h10408000;
      31011: inst = 32'hc4044e1;
      31012: inst = 32'h8220000;
      31013: inst = 32'h10408000;
      31014: inst = 32'hc4044e2;
      31015: inst = 32'h8220000;
      31016: inst = 32'h10408000;
      31017: inst = 32'hc4044e3;
      31018: inst = 32'h8220000;
      31019: inst = 32'h10408000;
      31020: inst = 32'hc4044e4;
      31021: inst = 32'h8220000;
      31022: inst = 32'h10408000;
      31023: inst = 32'hc4044e5;
      31024: inst = 32'h8220000;
      31025: inst = 32'h10408000;
      31026: inst = 32'hc4044e6;
      31027: inst = 32'h8220000;
      31028: inst = 32'h10408000;
      31029: inst = 32'hc4044e7;
      31030: inst = 32'h8220000;
      31031: inst = 32'h10408000;
      31032: inst = 32'hc4044e8;
      31033: inst = 32'h8220000;
      31034: inst = 32'h10408000;
      31035: inst = 32'hc4044e9;
      31036: inst = 32'h8220000;
      31037: inst = 32'h10408000;
      31038: inst = 32'hc4044ea;
      31039: inst = 32'h8220000;
      31040: inst = 32'h10408000;
      31041: inst = 32'hc4044eb;
      31042: inst = 32'h8220000;
      31043: inst = 32'h10408000;
      31044: inst = 32'hc4044ec;
      31045: inst = 32'h8220000;
      31046: inst = 32'h10408000;
      31047: inst = 32'hc4044ed;
      31048: inst = 32'h8220000;
      31049: inst = 32'h10408000;
      31050: inst = 32'hc4044ee;
      31051: inst = 32'h8220000;
      31052: inst = 32'h10408000;
      31053: inst = 32'hc4044ef;
      31054: inst = 32'h8220000;
      31055: inst = 32'h10408000;
      31056: inst = 32'hc4044f0;
      31057: inst = 32'h8220000;
      31058: inst = 32'h10408000;
      31059: inst = 32'hc4044f1;
      31060: inst = 32'h8220000;
      31061: inst = 32'h10408000;
      31062: inst = 32'hc4044f2;
      31063: inst = 32'h8220000;
      31064: inst = 32'h10408000;
      31065: inst = 32'hc4044f3;
      31066: inst = 32'h8220000;
      31067: inst = 32'h10408000;
      31068: inst = 32'hc4044f4;
      31069: inst = 32'h8220000;
      31070: inst = 32'h10408000;
      31071: inst = 32'hc4044f5;
      31072: inst = 32'h8220000;
      31073: inst = 32'h10408000;
      31074: inst = 32'hc4044f6;
      31075: inst = 32'h8220000;
      31076: inst = 32'h10408000;
      31077: inst = 32'hc4044f7;
      31078: inst = 32'h8220000;
      31079: inst = 32'h10408000;
      31080: inst = 32'hc4044f8;
      31081: inst = 32'h8220000;
      31082: inst = 32'h10408000;
      31083: inst = 32'hc4044f9;
      31084: inst = 32'h8220000;
      31085: inst = 32'h10408000;
      31086: inst = 32'hc4044fa;
      31087: inst = 32'h8220000;
      31088: inst = 32'h10408000;
      31089: inst = 32'hc4044fb;
      31090: inst = 32'h8220000;
      31091: inst = 32'h10408000;
      31092: inst = 32'hc4044fc;
      31093: inst = 32'h8220000;
      31094: inst = 32'h10408000;
      31095: inst = 32'hc4044fd;
      31096: inst = 32'h8220000;
      31097: inst = 32'h10408000;
      31098: inst = 32'hc4044fe;
      31099: inst = 32'h8220000;
      31100: inst = 32'h10408000;
      31101: inst = 32'hc4044ff;
      31102: inst = 32'h8220000;
      31103: inst = 32'h10408000;
      31104: inst = 32'hc404500;
      31105: inst = 32'h8220000;
      31106: inst = 32'h10408000;
      31107: inst = 32'hc404501;
      31108: inst = 32'h8220000;
      31109: inst = 32'h10408000;
      31110: inst = 32'hc404502;
      31111: inst = 32'h8220000;
      31112: inst = 32'h10408000;
      31113: inst = 32'hc404503;
      31114: inst = 32'h8220000;
      31115: inst = 32'h10408000;
      31116: inst = 32'hc404504;
      31117: inst = 32'h8220000;
      31118: inst = 32'h10408000;
      31119: inst = 32'hc404505;
      31120: inst = 32'h8220000;
      31121: inst = 32'h10408000;
      31122: inst = 32'hc404506;
      31123: inst = 32'h8220000;
      31124: inst = 32'h10408000;
      31125: inst = 32'hc404507;
      31126: inst = 32'h8220000;
      31127: inst = 32'h10408000;
      31128: inst = 32'hc404508;
      31129: inst = 32'h8220000;
      31130: inst = 32'h10408000;
      31131: inst = 32'hc404509;
      31132: inst = 32'h8220000;
      31133: inst = 32'h10408000;
      31134: inst = 32'hc40450a;
      31135: inst = 32'h8220000;
      31136: inst = 32'h10408000;
      31137: inst = 32'hc40450b;
      31138: inst = 32'h8220000;
      31139: inst = 32'h10408000;
      31140: inst = 32'hc40450f;
      31141: inst = 32'h8220000;
      31142: inst = 32'h10408000;
      31143: inst = 32'hc404512;
      31144: inst = 32'h8220000;
      31145: inst = 32'h10408000;
      31146: inst = 32'hc404513;
      31147: inst = 32'h8220000;
      31148: inst = 32'h10408000;
      31149: inst = 32'hc404523;
      31150: inst = 32'h8220000;
      31151: inst = 32'h10408000;
      31152: inst = 32'hc404524;
      31153: inst = 32'h8220000;
      31154: inst = 32'h10408000;
      31155: inst = 32'hc404525;
      31156: inst = 32'h8220000;
      31157: inst = 32'h10408000;
      31158: inst = 32'hc404526;
      31159: inst = 32'h8220000;
      31160: inst = 32'h10408000;
      31161: inst = 32'hc404527;
      31162: inst = 32'h8220000;
      31163: inst = 32'h10408000;
      31164: inst = 32'hc404528;
      31165: inst = 32'h8220000;
      31166: inst = 32'h10408000;
      31167: inst = 32'hc404529;
      31168: inst = 32'h8220000;
      31169: inst = 32'h10408000;
      31170: inst = 32'hc40452a;
      31171: inst = 32'h8220000;
      31172: inst = 32'h10408000;
      31173: inst = 32'hc40452b;
      31174: inst = 32'h8220000;
      31175: inst = 32'h10408000;
      31176: inst = 32'hc40452c;
      31177: inst = 32'h8220000;
      31178: inst = 32'h10408000;
      31179: inst = 32'hc40452d;
      31180: inst = 32'h8220000;
      31181: inst = 32'h10408000;
      31182: inst = 32'hc40452e;
      31183: inst = 32'h8220000;
      31184: inst = 32'h10408000;
      31185: inst = 32'hc40452f;
      31186: inst = 32'h8220000;
      31187: inst = 32'h10408000;
      31188: inst = 32'hc404530;
      31189: inst = 32'h8220000;
      31190: inst = 32'h10408000;
      31191: inst = 32'hc404531;
      31192: inst = 32'h8220000;
      31193: inst = 32'h10408000;
      31194: inst = 32'hc404532;
      31195: inst = 32'h8220000;
      31196: inst = 32'h10408000;
      31197: inst = 32'hc404533;
      31198: inst = 32'h8220000;
      31199: inst = 32'h10408000;
      31200: inst = 32'hc404534;
      31201: inst = 32'h8220000;
      31202: inst = 32'h10408000;
      31203: inst = 32'hc404535;
      31204: inst = 32'h8220000;
      31205: inst = 32'h10408000;
      31206: inst = 32'hc404536;
      31207: inst = 32'h8220000;
      31208: inst = 32'h10408000;
      31209: inst = 32'hc404537;
      31210: inst = 32'h8220000;
      31211: inst = 32'h10408000;
      31212: inst = 32'hc404538;
      31213: inst = 32'h8220000;
      31214: inst = 32'h10408000;
      31215: inst = 32'hc404539;
      31216: inst = 32'h8220000;
      31217: inst = 32'h10408000;
      31218: inst = 32'hc40453a;
      31219: inst = 32'h8220000;
      31220: inst = 32'h10408000;
      31221: inst = 32'hc40453b;
      31222: inst = 32'h8220000;
      31223: inst = 32'h10408000;
      31224: inst = 32'hc40453c;
      31225: inst = 32'h8220000;
      31226: inst = 32'h10408000;
      31227: inst = 32'hc40453d;
      31228: inst = 32'h8220000;
      31229: inst = 32'h10408000;
      31230: inst = 32'hc40453e;
      31231: inst = 32'h8220000;
      31232: inst = 32'h10408000;
      31233: inst = 32'hc40453f;
      31234: inst = 32'h8220000;
      31235: inst = 32'h10408000;
      31236: inst = 32'hc404540;
      31237: inst = 32'h8220000;
      31238: inst = 32'h10408000;
      31239: inst = 32'hc404541;
      31240: inst = 32'h8220000;
      31241: inst = 32'h10408000;
      31242: inst = 32'hc404542;
      31243: inst = 32'h8220000;
      31244: inst = 32'h10408000;
      31245: inst = 32'hc404543;
      31246: inst = 32'h8220000;
      31247: inst = 32'h10408000;
      31248: inst = 32'hc404544;
      31249: inst = 32'h8220000;
      31250: inst = 32'h10408000;
      31251: inst = 32'hc404545;
      31252: inst = 32'h8220000;
      31253: inst = 32'h10408000;
      31254: inst = 32'hc404546;
      31255: inst = 32'h8220000;
      31256: inst = 32'h10408000;
      31257: inst = 32'hc404547;
      31258: inst = 32'h8220000;
      31259: inst = 32'h10408000;
      31260: inst = 32'hc404548;
      31261: inst = 32'h8220000;
      31262: inst = 32'h10408000;
      31263: inst = 32'hc404549;
      31264: inst = 32'h8220000;
      31265: inst = 32'h10408000;
      31266: inst = 32'hc40454a;
      31267: inst = 32'h8220000;
      31268: inst = 32'h10408000;
      31269: inst = 32'hc40454b;
      31270: inst = 32'h8220000;
      31271: inst = 32'h10408000;
      31272: inst = 32'hc40454c;
      31273: inst = 32'h8220000;
      31274: inst = 32'h10408000;
      31275: inst = 32'hc40454d;
      31276: inst = 32'h8220000;
      31277: inst = 32'h10408000;
      31278: inst = 32'hc40454e;
      31279: inst = 32'h8220000;
      31280: inst = 32'h10408000;
      31281: inst = 32'hc40454f;
      31282: inst = 32'h8220000;
      31283: inst = 32'h10408000;
      31284: inst = 32'hc404550;
      31285: inst = 32'h8220000;
      31286: inst = 32'h10408000;
      31287: inst = 32'hc404551;
      31288: inst = 32'h8220000;
      31289: inst = 32'h10408000;
      31290: inst = 32'hc404552;
      31291: inst = 32'h8220000;
      31292: inst = 32'h10408000;
      31293: inst = 32'hc404553;
      31294: inst = 32'h8220000;
      31295: inst = 32'h10408000;
      31296: inst = 32'hc404554;
      31297: inst = 32'h8220000;
      31298: inst = 32'h10408000;
      31299: inst = 32'hc404555;
      31300: inst = 32'h8220000;
      31301: inst = 32'h10408000;
      31302: inst = 32'hc404556;
      31303: inst = 32'h8220000;
      31304: inst = 32'h10408000;
      31305: inst = 32'hc404557;
      31306: inst = 32'h8220000;
      31307: inst = 32'h10408000;
      31308: inst = 32'hc404558;
      31309: inst = 32'h8220000;
      31310: inst = 32'h10408000;
      31311: inst = 32'hc404559;
      31312: inst = 32'h8220000;
      31313: inst = 32'h10408000;
      31314: inst = 32'hc40455a;
      31315: inst = 32'h8220000;
      31316: inst = 32'h10408000;
      31317: inst = 32'hc40455b;
      31318: inst = 32'h8220000;
      31319: inst = 32'h10408000;
      31320: inst = 32'hc40455c;
      31321: inst = 32'h8220000;
      31322: inst = 32'h10408000;
      31323: inst = 32'hc40455d;
      31324: inst = 32'h8220000;
      31325: inst = 32'h10408000;
      31326: inst = 32'hc40455e;
      31327: inst = 32'h8220000;
      31328: inst = 32'h10408000;
      31329: inst = 32'hc40455f;
      31330: inst = 32'h8220000;
      31331: inst = 32'h10408000;
      31332: inst = 32'hc404560;
      31333: inst = 32'h8220000;
      31334: inst = 32'h10408000;
      31335: inst = 32'hc404561;
      31336: inst = 32'h8220000;
      31337: inst = 32'h10408000;
      31338: inst = 32'hc404562;
      31339: inst = 32'h8220000;
      31340: inst = 32'h10408000;
      31341: inst = 32'hc404563;
      31342: inst = 32'h8220000;
      31343: inst = 32'h10408000;
      31344: inst = 32'hc404564;
      31345: inst = 32'h8220000;
      31346: inst = 32'h10408000;
      31347: inst = 32'hc404565;
      31348: inst = 32'h8220000;
      31349: inst = 32'h10408000;
      31350: inst = 32'hc404566;
      31351: inst = 32'h8220000;
      31352: inst = 32'h10408000;
      31353: inst = 32'hc404567;
      31354: inst = 32'h8220000;
      31355: inst = 32'h10408000;
      31356: inst = 32'hc404568;
      31357: inst = 32'h8220000;
      31358: inst = 32'h10408000;
      31359: inst = 32'hc404569;
      31360: inst = 32'h8220000;
      31361: inst = 32'h10408000;
      31362: inst = 32'hc40456a;
      31363: inst = 32'h8220000;
      31364: inst = 32'h10408000;
      31365: inst = 32'hc40456b;
      31366: inst = 32'h8220000;
      31367: inst = 32'h10408000;
      31368: inst = 32'hc40456f;
      31369: inst = 32'h8220000;
      31370: inst = 32'h10408000;
      31371: inst = 32'hc40457a;
      31372: inst = 32'h8220000;
      31373: inst = 32'h10408000;
      31374: inst = 32'hc40457b;
      31375: inst = 32'h8220000;
      31376: inst = 32'h10408000;
      31377: inst = 32'hc40457c;
      31378: inst = 32'h8220000;
      31379: inst = 32'h10408000;
      31380: inst = 32'hc404583;
      31381: inst = 32'h8220000;
      31382: inst = 32'h10408000;
      31383: inst = 32'hc404584;
      31384: inst = 32'h8220000;
      31385: inst = 32'h10408000;
      31386: inst = 32'hc404585;
      31387: inst = 32'h8220000;
      31388: inst = 32'h10408000;
      31389: inst = 32'hc404586;
      31390: inst = 32'h8220000;
      31391: inst = 32'h10408000;
      31392: inst = 32'hc404587;
      31393: inst = 32'h8220000;
      31394: inst = 32'h10408000;
      31395: inst = 32'hc404588;
      31396: inst = 32'h8220000;
      31397: inst = 32'h10408000;
      31398: inst = 32'hc404589;
      31399: inst = 32'h8220000;
      31400: inst = 32'h10408000;
      31401: inst = 32'hc40458a;
      31402: inst = 32'h8220000;
      31403: inst = 32'h10408000;
      31404: inst = 32'hc40458b;
      31405: inst = 32'h8220000;
      31406: inst = 32'h10408000;
      31407: inst = 32'hc40458c;
      31408: inst = 32'h8220000;
      31409: inst = 32'h10408000;
      31410: inst = 32'hc40458d;
      31411: inst = 32'h8220000;
      31412: inst = 32'h10408000;
      31413: inst = 32'hc40458e;
      31414: inst = 32'h8220000;
      31415: inst = 32'h10408000;
      31416: inst = 32'hc40458f;
      31417: inst = 32'h8220000;
      31418: inst = 32'h10408000;
      31419: inst = 32'hc404590;
      31420: inst = 32'h8220000;
      31421: inst = 32'h10408000;
      31422: inst = 32'hc404591;
      31423: inst = 32'h8220000;
      31424: inst = 32'h10408000;
      31425: inst = 32'hc404592;
      31426: inst = 32'h8220000;
      31427: inst = 32'h10408000;
      31428: inst = 32'hc404593;
      31429: inst = 32'h8220000;
      31430: inst = 32'h10408000;
      31431: inst = 32'hc404594;
      31432: inst = 32'h8220000;
      31433: inst = 32'h10408000;
      31434: inst = 32'hc404595;
      31435: inst = 32'h8220000;
      31436: inst = 32'h10408000;
      31437: inst = 32'hc404596;
      31438: inst = 32'h8220000;
      31439: inst = 32'h10408000;
      31440: inst = 32'hc404597;
      31441: inst = 32'h8220000;
      31442: inst = 32'h10408000;
      31443: inst = 32'hc404598;
      31444: inst = 32'h8220000;
      31445: inst = 32'h10408000;
      31446: inst = 32'hc404599;
      31447: inst = 32'h8220000;
      31448: inst = 32'h10408000;
      31449: inst = 32'hc40459a;
      31450: inst = 32'h8220000;
      31451: inst = 32'h10408000;
      31452: inst = 32'hc40459b;
      31453: inst = 32'h8220000;
      31454: inst = 32'h10408000;
      31455: inst = 32'hc40459c;
      31456: inst = 32'h8220000;
      31457: inst = 32'h10408000;
      31458: inst = 32'hc40459d;
      31459: inst = 32'h8220000;
      31460: inst = 32'h10408000;
      31461: inst = 32'hc40459e;
      31462: inst = 32'h8220000;
      31463: inst = 32'h10408000;
      31464: inst = 32'hc40459f;
      31465: inst = 32'h8220000;
      31466: inst = 32'h10408000;
      31467: inst = 32'hc4045a0;
      31468: inst = 32'h8220000;
      31469: inst = 32'h10408000;
      31470: inst = 32'hc4045a1;
      31471: inst = 32'h8220000;
      31472: inst = 32'h10408000;
      31473: inst = 32'hc4045a2;
      31474: inst = 32'h8220000;
      31475: inst = 32'h10408000;
      31476: inst = 32'hc4045a3;
      31477: inst = 32'h8220000;
      31478: inst = 32'h10408000;
      31479: inst = 32'hc4045a4;
      31480: inst = 32'h8220000;
      31481: inst = 32'h10408000;
      31482: inst = 32'hc4045a5;
      31483: inst = 32'h8220000;
      31484: inst = 32'h10408000;
      31485: inst = 32'hc4045a6;
      31486: inst = 32'h8220000;
      31487: inst = 32'h10408000;
      31488: inst = 32'hc4045a7;
      31489: inst = 32'h8220000;
      31490: inst = 32'h10408000;
      31491: inst = 32'hc4045a8;
      31492: inst = 32'h8220000;
      31493: inst = 32'h10408000;
      31494: inst = 32'hc4045a9;
      31495: inst = 32'h8220000;
      31496: inst = 32'h10408000;
      31497: inst = 32'hc4045aa;
      31498: inst = 32'h8220000;
      31499: inst = 32'h10408000;
      31500: inst = 32'hc4045ab;
      31501: inst = 32'h8220000;
      31502: inst = 32'h10408000;
      31503: inst = 32'hc4045ac;
      31504: inst = 32'h8220000;
      31505: inst = 32'h10408000;
      31506: inst = 32'hc4045ad;
      31507: inst = 32'h8220000;
      31508: inst = 32'h10408000;
      31509: inst = 32'hc4045ae;
      31510: inst = 32'h8220000;
      31511: inst = 32'h10408000;
      31512: inst = 32'hc4045af;
      31513: inst = 32'h8220000;
      31514: inst = 32'h10408000;
      31515: inst = 32'hc4045b0;
      31516: inst = 32'h8220000;
      31517: inst = 32'h10408000;
      31518: inst = 32'hc4045b1;
      31519: inst = 32'h8220000;
      31520: inst = 32'h10408000;
      31521: inst = 32'hc4045b2;
      31522: inst = 32'h8220000;
      31523: inst = 32'h10408000;
      31524: inst = 32'hc4045b3;
      31525: inst = 32'h8220000;
      31526: inst = 32'h10408000;
      31527: inst = 32'hc4045b4;
      31528: inst = 32'h8220000;
      31529: inst = 32'h10408000;
      31530: inst = 32'hc4045b5;
      31531: inst = 32'h8220000;
      31532: inst = 32'h10408000;
      31533: inst = 32'hc4045b6;
      31534: inst = 32'h8220000;
      31535: inst = 32'h10408000;
      31536: inst = 32'hc4045b7;
      31537: inst = 32'h8220000;
      31538: inst = 32'h10408000;
      31539: inst = 32'hc4045b8;
      31540: inst = 32'h8220000;
      31541: inst = 32'h10408000;
      31542: inst = 32'hc4045b9;
      31543: inst = 32'h8220000;
      31544: inst = 32'h10408000;
      31545: inst = 32'hc4045ba;
      31546: inst = 32'h8220000;
      31547: inst = 32'h10408000;
      31548: inst = 32'hc4045bb;
      31549: inst = 32'h8220000;
      31550: inst = 32'h10408000;
      31551: inst = 32'hc4045bc;
      31552: inst = 32'h8220000;
      31553: inst = 32'h10408000;
      31554: inst = 32'hc4045bd;
      31555: inst = 32'h8220000;
      31556: inst = 32'h10408000;
      31557: inst = 32'hc4045be;
      31558: inst = 32'h8220000;
      31559: inst = 32'h10408000;
      31560: inst = 32'hc4045bf;
      31561: inst = 32'h8220000;
      31562: inst = 32'h10408000;
      31563: inst = 32'hc4045c0;
      31564: inst = 32'h8220000;
      31565: inst = 32'h10408000;
      31566: inst = 32'hc4045c1;
      31567: inst = 32'h8220000;
      31568: inst = 32'h10408000;
      31569: inst = 32'hc4045c2;
      31570: inst = 32'h8220000;
      31571: inst = 32'h10408000;
      31572: inst = 32'hc4045c3;
      31573: inst = 32'h8220000;
      31574: inst = 32'h10408000;
      31575: inst = 32'hc4045c4;
      31576: inst = 32'h8220000;
      31577: inst = 32'h10408000;
      31578: inst = 32'hc4045c5;
      31579: inst = 32'h8220000;
      31580: inst = 32'h10408000;
      31581: inst = 32'hc4045c6;
      31582: inst = 32'h8220000;
      31583: inst = 32'h10408000;
      31584: inst = 32'hc4045c7;
      31585: inst = 32'h8220000;
      31586: inst = 32'h10408000;
      31587: inst = 32'hc4045c8;
      31588: inst = 32'h8220000;
      31589: inst = 32'h10408000;
      31590: inst = 32'hc4045c9;
      31591: inst = 32'h8220000;
      31592: inst = 32'h10408000;
      31593: inst = 32'hc4045ca;
      31594: inst = 32'h8220000;
      31595: inst = 32'h10408000;
      31596: inst = 32'hc4045cb;
      31597: inst = 32'h8220000;
      31598: inst = 32'h10408000;
      31599: inst = 32'hc4045cf;
      31600: inst = 32'h8220000;
      31601: inst = 32'h10408000;
      31602: inst = 32'hc4045d0;
      31603: inst = 32'h8220000;
      31604: inst = 32'h10408000;
      31605: inst = 32'hc4045d4;
      31606: inst = 32'h8220000;
      31607: inst = 32'h10408000;
      31608: inst = 32'hc4045d5;
      31609: inst = 32'h8220000;
      31610: inst = 32'h10408000;
      31611: inst = 32'hc4045d6;
      31612: inst = 32'h8220000;
      31613: inst = 32'h10408000;
      31614: inst = 32'hc4045d7;
      31615: inst = 32'h8220000;
      31616: inst = 32'h10408000;
      31617: inst = 32'hc4045da;
      31618: inst = 32'h8220000;
      31619: inst = 32'h10408000;
      31620: inst = 32'hc4045db;
      31621: inst = 32'h8220000;
      31622: inst = 32'h10408000;
      31623: inst = 32'hc4045e3;
      31624: inst = 32'h8220000;
      31625: inst = 32'h10408000;
      31626: inst = 32'hc4045e4;
      31627: inst = 32'h8220000;
      31628: inst = 32'h10408000;
      31629: inst = 32'hc4045e5;
      31630: inst = 32'h8220000;
      31631: inst = 32'h10408000;
      31632: inst = 32'hc4045e6;
      31633: inst = 32'h8220000;
      31634: inst = 32'h10408000;
      31635: inst = 32'hc4045e7;
      31636: inst = 32'h8220000;
      31637: inst = 32'h10408000;
      31638: inst = 32'hc4045e8;
      31639: inst = 32'h8220000;
      31640: inst = 32'h10408000;
      31641: inst = 32'hc4045e9;
      31642: inst = 32'h8220000;
      31643: inst = 32'h10408000;
      31644: inst = 32'hc4045ea;
      31645: inst = 32'h8220000;
      31646: inst = 32'h10408000;
      31647: inst = 32'hc4045eb;
      31648: inst = 32'h8220000;
      31649: inst = 32'h10408000;
      31650: inst = 32'hc4045ec;
      31651: inst = 32'h8220000;
      31652: inst = 32'h10408000;
      31653: inst = 32'hc4045ed;
      31654: inst = 32'h8220000;
      31655: inst = 32'h10408000;
      31656: inst = 32'hc4045ee;
      31657: inst = 32'h8220000;
      31658: inst = 32'h10408000;
      31659: inst = 32'hc4045ef;
      31660: inst = 32'h8220000;
      31661: inst = 32'h10408000;
      31662: inst = 32'hc4045f0;
      31663: inst = 32'h8220000;
      31664: inst = 32'h10408000;
      31665: inst = 32'hc4045f1;
      31666: inst = 32'h8220000;
      31667: inst = 32'h10408000;
      31668: inst = 32'hc4045f2;
      31669: inst = 32'h8220000;
      31670: inst = 32'h10408000;
      31671: inst = 32'hc4045f3;
      31672: inst = 32'h8220000;
      31673: inst = 32'h10408000;
      31674: inst = 32'hc4045f4;
      31675: inst = 32'h8220000;
      31676: inst = 32'h10408000;
      31677: inst = 32'hc4045f5;
      31678: inst = 32'h8220000;
      31679: inst = 32'h10408000;
      31680: inst = 32'hc4045f6;
      31681: inst = 32'h8220000;
      31682: inst = 32'h10408000;
      31683: inst = 32'hc4045f7;
      31684: inst = 32'h8220000;
      31685: inst = 32'h10408000;
      31686: inst = 32'hc4045f8;
      31687: inst = 32'h8220000;
      31688: inst = 32'h10408000;
      31689: inst = 32'hc4045f9;
      31690: inst = 32'h8220000;
      31691: inst = 32'h10408000;
      31692: inst = 32'hc4045fa;
      31693: inst = 32'h8220000;
      31694: inst = 32'h10408000;
      31695: inst = 32'hc4045fb;
      31696: inst = 32'h8220000;
      31697: inst = 32'h10408000;
      31698: inst = 32'hc4045fc;
      31699: inst = 32'h8220000;
      31700: inst = 32'h10408000;
      31701: inst = 32'hc4045fd;
      31702: inst = 32'h8220000;
      31703: inst = 32'h10408000;
      31704: inst = 32'hc4045fe;
      31705: inst = 32'h8220000;
      31706: inst = 32'h10408000;
      31707: inst = 32'hc4045ff;
      31708: inst = 32'h8220000;
      31709: inst = 32'h10408000;
      31710: inst = 32'hc404600;
      31711: inst = 32'h8220000;
      31712: inst = 32'h10408000;
      31713: inst = 32'hc404601;
      31714: inst = 32'h8220000;
      31715: inst = 32'h10408000;
      31716: inst = 32'hc404602;
      31717: inst = 32'h8220000;
      31718: inst = 32'h10408000;
      31719: inst = 32'hc404603;
      31720: inst = 32'h8220000;
      31721: inst = 32'h10408000;
      31722: inst = 32'hc404604;
      31723: inst = 32'h8220000;
      31724: inst = 32'h10408000;
      31725: inst = 32'hc404605;
      31726: inst = 32'h8220000;
      31727: inst = 32'h10408000;
      31728: inst = 32'hc404606;
      31729: inst = 32'h8220000;
      31730: inst = 32'h10408000;
      31731: inst = 32'hc404607;
      31732: inst = 32'h8220000;
      31733: inst = 32'h10408000;
      31734: inst = 32'hc404608;
      31735: inst = 32'h8220000;
      31736: inst = 32'h10408000;
      31737: inst = 32'hc404609;
      31738: inst = 32'h8220000;
      31739: inst = 32'h10408000;
      31740: inst = 32'hc40460a;
      31741: inst = 32'h8220000;
      31742: inst = 32'h10408000;
      31743: inst = 32'hc40460b;
      31744: inst = 32'h8220000;
      31745: inst = 32'h10408000;
      31746: inst = 32'hc40460c;
      31747: inst = 32'h8220000;
      31748: inst = 32'h10408000;
      31749: inst = 32'hc40460d;
      31750: inst = 32'h8220000;
      31751: inst = 32'h10408000;
      31752: inst = 32'hc40460e;
      31753: inst = 32'h8220000;
      31754: inst = 32'h10408000;
      31755: inst = 32'hc40460f;
      31756: inst = 32'h8220000;
      31757: inst = 32'h10408000;
      31758: inst = 32'hc404610;
      31759: inst = 32'h8220000;
      31760: inst = 32'h10408000;
      31761: inst = 32'hc404611;
      31762: inst = 32'h8220000;
      31763: inst = 32'h10408000;
      31764: inst = 32'hc404612;
      31765: inst = 32'h8220000;
      31766: inst = 32'h10408000;
      31767: inst = 32'hc404613;
      31768: inst = 32'h8220000;
      31769: inst = 32'h10408000;
      31770: inst = 32'hc404614;
      31771: inst = 32'h8220000;
      31772: inst = 32'h10408000;
      31773: inst = 32'hc404615;
      31774: inst = 32'h8220000;
      31775: inst = 32'h10408000;
      31776: inst = 32'hc404616;
      31777: inst = 32'h8220000;
      31778: inst = 32'h10408000;
      31779: inst = 32'hc404617;
      31780: inst = 32'h8220000;
      31781: inst = 32'h10408000;
      31782: inst = 32'hc404618;
      31783: inst = 32'h8220000;
      31784: inst = 32'h10408000;
      31785: inst = 32'hc404619;
      31786: inst = 32'h8220000;
      31787: inst = 32'h10408000;
      31788: inst = 32'hc40461a;
      31789: inst = 32'h8220000;
      31790: inst = 32'h10408000;
      31791: inst = 32'hc40461b;
      31792: inst = 32'h8220000;
      31793: inst = 32'h10408000;
      31794: inst = 32'hc40461c;
      31795: inst = 32'h8220000;
      31796: inst = 32'h10408000;
      31797: inst = 32'hc40461d;
      31798: inst = 32'h8220000;
      31799: inst = 32'h10408000;
      31800: inst = 32'hc40461e;
      31801: inst = 32'h8220000;
      31802: inst = 32'h10408000;
      31803: inst = 32'hc40461f;
      31804: inst = 32'h8220000;
      31805: inst = 32'h10408000;
      31806: inst = 32'hc404620;
      31807: inst = 32'h8220000;
      31808: inst = 32'h10408000;
      31809: inst = 32'hc404621;
      31810: inst = 32'h8220000;
      31811: inst = 32'h10408000;
      31812: inst = 32'hc404622;
      31813: inst = 32'h8220000;
      31814: inst = 32'h10408000;
      31815: inst = 32'hc404623;
      31816: inst = 32'h8220000;
      31817: inst = 32'h10408000;
      31818: inst = 32'hc404624;
      31819: inst = 32'h8220000;
      31820: inst = 32'h10408000;
      31821: inst = 32'hc404625;
      31822: inst = 32'h8220000;
      31823: inst = 32'h10408000;
      31824: inst = 32'hc404626;
      31825: inst = 32'h8220000;
      31826: inst = 32'h10408000;
      31827: inst = 32'hc404627;
      31828: inst = 32'h8220000;
      31829: inst = 32'h10408000;
      31830: inst = 32'hc404628;
      31831: inst = 32'h8220000;
      31832: inst = 32'h10408000;
      31833: inst = 32'hc404629;
      31834: inst = 32'h8220000;
      31835: inst = 32'h10408000;
      31836: inst = 32'hc40462a;
      31837: inst = 32'h8220000;
      31838: inst = 32'h10408000;
      31839: inst = 32'hc40462b;
      31840: inst = 32'h8220000;
      31841: inst = 32'h10408000;
      31842: inst = 32'hc40462f;
      31843: inst = 32'h8220000;
      31844: inst = 32'h10408000;
      31845: inst = 32'hc404630;
      31846: inst = 32'h8220000;
      31847: inst = 32'h10408000;
      31848: inst = 32'hc404631;
      31849: inst = 32'h8220000;
      31850: inst = 32'h10408000;
      31851: inst = 32'hc404632;
      31852: inst = 32'h8220000;
      31853: inst = 32'h10408000;
      31854: inst = 32'hc404633;
      31855: inst = 32'h8220000;
      31856: inst = 32'h10408000;
      31857: inst = 32'hc404634;
      31858: inst = 32'h8220000;
      31859: inst = 32'h10408000;
      31860: inst = 32'hc404635;
      31861: inst = 32'h8220000;
      31862: inst = 32'h10408000;
      31863: inst = 32'hc404636;
      31864: inst = 32'h8220000;
      31865: inst = 32'h10408000;
      31866: inst = 32'hc404637;
      31867: inst = 32'h8220000;
      31868: inst = 32'h10408000;
      31869: inst = 32'hc404638;
      31870: inst = 32'h8220000;
      31871: inst = 32'h10408000;
      31872: inst = 32'hc404639;
      31873: inst = 32'h8220000;
      31874: inst = 32'h10408000;
      31875: inst = 32'hc40463a;
      31876: inst = 32'h8220000;
      31877: inst = 32'h10408000;
      31878: inst = 32'hc40463b;
      31879: inst = 32'h8220000;
      31880: inst = 32'h10408000;
      31881: inst = 32'hc40463c;
      31882: inst = 32'h8220000;
      31883: inst = 32'h10408000;
      31884: inst = 32'hc404643;
      31885: inst = 32'h8220000;
      31886: inst = 32'h10408000;
      31887: inst = 32'hc404644;
      31888: inst = 32'h8220000;
      31889: inst = 32'h10408000;
      31890: inst = 32'hc404645;
      31891: inst = 32'h8220000;
      31892: inst = 32'h10408000;
      31893: inst = 32'hc404646;
      31894: inst = 32'h8220000;
      31895: inst = 32'h10408000;
      31896: inst = 32'hc404647;
      31897: inst = 32'h8220000;
      31898: inst = 32'h10408000;
      31899: inst = 32'hc404648;
      31900: inst = 32'h8220000;
      31901: inst = 32'h10408000;
      31902: inst = 32'hc404649;
      31903: inst = 32'h8220000;
      31904: inst = 32'h10408000;
      31905: inst = 32'hc40464a;
      31906: inst = 32'h8220000;
      31907: inst = 32'h10408000;
      31908: inst = 32'hc40464b;
      31909: inst = 32'h8220000;
      31910: inst = 32'h10408000;
      31911: inst = 32'hc40464c;
      31912: inst = 32'h8220000;
      31913: inst = 32'h10408000;
      31914: inst = 32'hc40464d;
      31915: inst = 32'h8220000;
      31916: inst = 32'h10408000;
      31917: inst = 32'hc40467a;
      31918: inst = 32'h8220000;
      31919: inst = 32'h10408000;
      31920: inst = 32'hc40467b;
      31921: inst = 32'h8220000;
      31922: inst = 32'h10408000;
      31923: inst = 32'hc40467c;
      31924: inst = 32'h8220000;
      31925: inst = 32'h10408000;
      31926: inst = 32'hc40467d;
      31927: inst = 32'h8220000;
      31928: inst = 32'h10408000;
      31929: inst = 32'hc40467e;
      31930: inst = 32'h8220000;
      31931: inst = 32'h10408000;
      31932: inst = 32'hc40467f;
      31933: inst = 32'h8220000;
      31934: inst = 32'h10408000;
      31935: inst = 32'hc404680;
      31936: inst = 32'h8220000;
      31937: inst = 32'h10408000;
      31938: inst = 32'hc404681;
      31939: inst = 32'h8220000;
      31940: inst = 32'h10408000;
      31941: inst = 32'hc404682;
      31942: inst = 32'h8220000;
      31943: inst = 32'h10408000;
      31944: inst = 32'hc404683;
      31945: inst = 32'h8220000;
      31946: inst = 32'h10408000;
      31947: inst = 32'hc404684;
      31948: inst = 32'h8220000;
      31949: inst = 32'h10408000;
      31950: inst = 32'hc404685;
      31951: inst = 32'h8220000;
      31952: inst = 32'h10408000;
      31953: inst = 32'hc404686;
      31954: inst = 32'h8220000;
      31955: inst = 32'h10408000;
      31956: inst = 32'hc404687;
      31957: inst = 32'h8220000;
      31958: inst = 32'h10408000;
      31959: inst = 32'hc404688;
      31960: inst = 32'h8220000;
      31961: inst = 32'h10408000;
      31962: inst = 32'hc404689;
      31963: inst = 32'h8220000;
      31964: inst = 32'h10408000;
      31965: inst = 32'hc40468a;
      31966: inst = 32'h8220000;
      31967: inst = 32'h10408000;
      31968: inst = 32'hc40468b;
      31969: inst = 32'h8220000;
      31970: inst = 32'h10408000;
      31971: inst = 32'hc40468f;
      31972: inst = 32'h8220000;
      31973: inst = 32'h10408000;
      31974: inst = 32'hc404690;
      31975: inst = 32'h8220000;
      31976: inst = 32'h10408000;
      31977: inst = 32'hc404691;
      31978: inst = 32'h8220000;
      31979: inst = 32'h10408000;
      31980: inst = 32'hc404692;
      31981: inst = 32'h8220000;
      31982: inst = 32'h10408000;
      31983: inst = 32'hc404693;
      31984: inst = 32'h8220000;
      31985: inst = 32'h10408000;
      31986: inst = 32'hc404694;
      31987: inst = 32'h8220000;
      31988: inst = 32'h10408000;
      31989: inst = 32'hc404695;
      31990: inst = 32'h8220000;
      31991: inst = 32'h10408000;
      31992: inst = 32'hc404696;
      31993: inst = 32'h8220000;
      31994: inst = 32'h10408000;
      31995: inst = 32'hc404697;
      31996: inst = 32'h8220000;
      31997: inst = 32'h10408000;
      31998: inst = 32'hc404698;
      31999: inst = 32'h8220000;
      32000: inst = 32'h10408000;
      32001: inst = 32'hc404699;
      32002: inst = 32'h8220000;
      32003: inst = 32'h10408000;
      32004: inst = 32'hc40469a;
      32005: inst = 32'h8220000;
      32006: inst = 32'h10408000;
      32007: inst = 32'hc40469b;
      32008: inst = 32'h8220000;
      32009: inst = 32'h10408000;
      32010: inst = 32'hc40469c;
      32011: inst = 32'h8220000;
      32012: inst = 32'h10408000;
      32013: inst = 32'hc4046a3;
      32014: inst = 32'h8220000;
      32015: inst = 32'h10408000;
      32016: inst = 32'hc4046a4;
      32017: inst = 32'h8220000;
      32018: inst = 32'h10408000;
      32019: inst = 32'hc4046a5;
      32020: inst = 32'h8220000;
      32021: inst = 32'h10408000;
      32022: inst = 32'hc4046a6;
      32023: inst = 32'h8220000;
      32024: inst = 32'h10408000;
      32025: inst = 32'hc4046a7;
      32026: inst = 32'h8220000;
      32027: inst = 32'h10408000;
      32028: inst = 32'hc4046a8;
      32029: inst = 32'h8220000;
      32030: inst = 32'h10408000;
      32031: inst = 32'hc4046a9;
      32032: inst = 32'h8220000;
      32033: inst = 32'h10408000;
      32034: inst = 32'hc4046aa;
      32035: inst = 32'h8220000;
      32036: inst = 32'h10408000;
      32037: inst = 32'hc4046ab;
      32038: inst = 32'h8220000;
      32039: inst = 32'h10408000;
      32040: inst = 32'hc4046ac;
      32041: inst = 32'h8220000;
      32042: inst = 32'h10408000;
      32043: inst = 32'hc4046ad;
      32044: inst = 32'h8220000;
      32045: inst = 32'h10408000;
      32046: inst = 32'hc4046da;
      32047: inst = 32'h8220000;
      32048: inst = 32'h10408000;
      32049: inst = 32'hc4046db;
      32050: inst = 32'h8220000;
      32051: inst = 32'h10408000;
      32052: inst = 32'hc4046dc;
      32053: inst = 32'h8220000;
      32054: inst = 32'h10408000;
      32055: inst = 32'hc4046dd;
      32056: inst = 32'h8220000;
      32057: inst = 32'h10408000;
      32058: inst = 32'hc4046de;
      32059: inst = 32'h8220000;
      32060: inst = 32'h10408000;
      32061: inst = 32'hc4046df;
      32062: inst = 32'h8220000;
      32063: inst = 32'h10408000;
      32064: inst = 32'hc4046e0;
      32065: inst = 32'h8220000;
      32066: inst = 32'h10408000;
      32067: inst = 32'hc4046e1;
      32068: inst = 32'h8220000;
      32069: inst = 32'h10408000;
      32070: inst = 32'hc4046e2;
      32071: inst = 32'h8220000;
      32072: inst = 32'h10408000;
      32073: inst = 32'hc4046e3;
      32074: inst = 32'h8220000;
      32075: inst = 32'h10408000;
      32076: inst = 32'hc4046e4;
      32077: inst = 32'h8220000;
      32078: inst = 32'h10408000;
      32079: inst = 32'hc4046e5;
      32080: inst = 32'h8220000;
      32081: inst = 32'h10408000;
      32082: inst = 32'hc4046e6;
      32083: inst = 32'h8220000;
      32084: inst = 32'h10408000;
      32085: inst = 32'hc4046e7;
      32086: inst = 32'h8220000;
      32087: inst = 32'h10408000;
      32088: inst = 32'hc4046e8;
      32089: inst = 32'h8220000;
      32090: inst = 32'h10408000;
      32091: inst = 32'hc4046e9;
      32092: inst = 32'h8220000;
      32093: inst = 32'h10408000;
      32094: inst = 32'hc4046ea;
      32095: inst = 32'h8220000;
      32096: inst = 32'h10408000;
      32097: inst = 32'hc4046eb;
      32098: inst = 32'h8220000;
      32099: inst = 32'h10408000;
      32100: inst = 32'hc4046ef;
      32101: inst = 32'h8220000;
      32102: inst = 32'h10408000;
      32103: inst = 32'hc4046f0;
      32104: inst = 32'h8220000;
      32105: inst = 32'h10408000;
      32106: inst = 32'hc4046f1;
      32107: inst = 32'h8220000;
      32108: inst = 32'h10408000;
      32109: inst = 32'hc4046f2;
      32110: inst = 32'h8220000;
      32111: inst = 32'h10408000;
      32112: inst = 32'hc4046f3;
      32113: inst = 32'h8220000;
      32114: inst = 32'h10408000;
      32115: inst = 32'hc4046f4;
      32116: inst = 32'h8220000;
      32117: inst = 32'h10408000;
      32118: inst = 32'hc4046f5;
      32119: inst = 32'h8220000;
      32120: inst = 32'h10408000;
      32121: inst = 32'hc4046f6;
      32122: inst = 32'h8220000;
      32123: inst = 32'h10408000;
      32124: inst = 32'hc4046f7;
      32125: inst = 32'h8220000;
      32126: inst = 32'h10408000;
      32127: inst = 32'hc4046f8;
      32128: inst = 32'h8220000;
      32129: inst = 32'h10408000;
      32130: inst = 32'hc4046f9;
      32131: inst = 32'h8220000;
      32132: inst = 32'h10408000;
      32133: inst = 32'hc4046fa;
      32134: inst = 32'h8220000;
      32135: inst = 32'h10408000;
      32136: inst = 32'hc4046fb;
      32137: inst = 32'h8220000;
      32138: inst = 32'h10408000;
      32139: inst = 32'hc4046fc;
      32140: inst = 32'h8220000;
      32141: inst = 32'h10408000;
      32142: inst = 32'hc404703;
      32143: inst = 32'h8220000;
      32144: inst = 32'h10408000;
      32145: inst = 32'hc404704;
      32146: inst = 32'h8220000;
      32147: inst = 32'h10408000;
      32148: inst = 32'hc404705;
      32149: inst = 32'h8220000;
      32150: inst = 32'h10408000;
      32151: inst = 32'hc404706;
      32152: inst = 32'h8220000;
      32153: inst = 32'h10408000;
      32154: inst = 32'hc404707;
      32155: inst = 32'h8220000;
      32156: inst = 32'h10408000;
      32157: inst = 32'hc404708;
      32158: inst = 32'h8220000;
      32159: inst = 32'h10408000;
      32160: inst = 32'hc404709;
      32161: inst = 32'h8220000;
      32162: inst = 32'h10408000;
      32163: inst = 32'hc40470a;
      32164: inst = 32'h8220000;
      32165: inst = 32'h10408000;
      32166: inst = 32'hc40470b;
      32167: inst = 32'h8220000;
      32168: inst = 32'h10408000;
      32169: inst = 32'hc40470c;
      32170: inst = 32'h8220000;
      32171: inst = 32'h10408000;
      32172: inst = 32'hc40470d;
      32173: inst = 32'h8220000;
      32174: inst = 32'h10408000;
      32175: inst = 32'hc40473a;
      32176: inst = 32'h8220000;
      32177: inst = 32'h10408000;
      32178: inst = 32'hc40473b;
      32179: inst = 32'h8220000;
      32180: inst = 32'h10408000;
      32181: inst = 32'hc40473c;
      32182: inst = 32'h8220000;
      32183: inst = 32'h10408000;
      32184: inst = 32'hc40473d;
      32185: inst = 32'h8220000;
      32186: inst = 32'h10408000;
      32187: inst = 32'hc40473e;
      32188: inst = 32'h8220000;
      32189: inst = 32'h10408000;
      32190: inst = 32'hc40473f;
      32191: inst = 32'h8220000;
      32192: inst = 32'h10408000;
      32193: inst = 32'hc404740;
      32194: inst = 32'h8220000;
      32195: inst = 32'h10408000;
      32196: inst = 32'hc404741;
      32197: inst = 32'h8220000;
      32198: inst = 32'h10408000;
      32199: inst = 32'hc404742;
      32200: inst = 32'h8220000;
      32201: inst = 32'h10408000;
      32202: inst = 32'hc404743;
      32203: inst = 32'h8220000;
      32204: inst = 32'h10408000;
      32205: inst = 32'hc404744;
      32206: inst = 32'h8220000;
      32207: inst = 32'h10408000;
      32208: inst = 32'hc404745;
      32209: inst = 32'h8220000;
      32210: inst = 32'h10408000;
      32211: inst = 32'hc404746;
      32212: inst = 32'h8220000;
      32213: inst = 32'h10408000;
      32214: inst = 32'hc404747;
      32215: inst = 32'h8220000;
      32216: inst = 32'h10408000;
      32217: inst = 32'hc404748;
      32218: inst = 32'h8220000;
      32219: inst = 32'h10408000;
      32220: inst = 32'hc404749;
      32221: inst = 32'h8220000;
      32222: inst = 32'h10408000;
      32223: inst = 32'hc40474a;
      32224: inst = 32'h8220000;
      32225: inst = 32'h10408000;
      32226: inst = 32'hc40474b;
      32227: inst = 32'h8220000;
      32228: inst = 32'h10408000;
      32229: inst = 32'hc40474f;
      32230: inst = 32'h8220000;
      32231: inst = 32'h10408000;
      32232: inst = 32'hc404750;
      32233: inst = 32'h8220000;
      32234: inst = 32'h10408000;
      32235: inst = 32'hc404751;
      32236: inst = 32'h8220000;
      32237: inst = 32'h10408000;
      32238: inst = 32'hc404752;
      32239: inst = 32'h8220000;
      32240: inst = 32'h10408000;
      32241: inst = 32'hc404753;
      32242: inst = 32'h8220000;
      32243: inst = 32'h10408000;
      32244: inst = 32'hc404754;
      32245: inst = 32'h8220000;
      32246: inst = 32'h10408000;
      32247: inst = 32'hc404755;
      32248: inst = 32'h8220000;
      32249: inst = 32'h10408000;
      32250: inst = 32'hc404756;
      32251: inst = 32'h8220000;
      32252: inst = 32'h10408000;
      32253: inst = 32'hc404757;
      32254: inst = 32'h8220000;
      32255: inst = 32'h10408000;
      32256: inst = 32'hc404758;
      32257: inst = 32'h8220000;
      32258: inst = 32'h10408000;
      32259: inst = 32'hc404759;
      32260: inst = 32'h8220000;
      32261: inst = 32'h10408000;
      32262: inst = 32'hc40475a;
      32263: inst = 32'h8220000;
      32264: inst = 32'h10408000;
      32265: inst = 32'hc40475b;
      32266: inst = 32'h8220000;
      32267: inst = 32'h10408000;
      32268: inst = 32'hc40475c;
      32269: inst = 32'h8220000;
      32270: inst = 32'h10408000;
      32271: inst = 32'hc404763;
      32272: inst = 32'h8220000;
      32273: inst = 32'h10408000;
      32274: inst = 32'hc404764;
      32275: inst = 32'h8220000;
      32276: inst = 32'h10408000;
      32277: inst = 32'hc404765;
      32278: inst = 32'h8220000;
      32279: inst = 32'h10408000;
      32280: inst = 32'hc404766;
      32281: inst = 32'h8220000;
      32282: inst = 32'h10408000;
      32283: inst = 32'hc404767;
      32284: inst = 32'h8220000;
      32285: inst = 32'h10408000;
      32286: inst = 32'hc404768;
      32287: inst = 32'h8220000;
      32288: inst = 32'h10408000;
      32289: inst = 32'hc404769;
      32290: inst = 32'h8220000;
      32291: inst = 32'h10408000;
      32292: inst = 32'hc40476a;
      32293: inst = 32'h8220000;
      32294: inst = 32'h10408000;
      32295: inst = 32'hc40476b;
      32296: inst = 32'h8220000;
      32297: inst = 32'h10408000;
      32298: inst = 32'hc40476c;
      32299: inst = 32'h8220000;
      32300: inst = 32'h10408000;
      32301: inst = 32'hc40476d;
      32302: inst = 32'h8220000;
      32303: inst = 32'h10408000;
      32304: inst = 32'hc404771;
      32305: inst = 32'h8220000;
      32306: inst = 32'h10408000;
      32307: inst = 32'hc404772;
      32308: inst = 32'h8220000;
      32309: inst = 32'h10408000;
      32310: inst = 32'hc404773;
      32311: inst = 32'h8220000;
      32312: inst = 32'h10408000;
      32313: inst = 32'hc404774;
      32314: inst = 32'h8220000;
      32315: inst = 32'h10408000;
      32316: inst = 32'hc404775;
      32317: inst = 32'h8220000;
      32318: inst = 32'h10408000;
      32319: inst = 32'hc404776;
      32320: inst = 32'h8220000;
      32321: inst = 32'h10408000;
      32322: inst = 32'hc404777;
      32323: inst = 32'h8220000;
      32324: inst = 32'h10408000;
      32325: inst = 32'hc404778;
      32326: inst = 32'h8220000;
      32327: inst = 32'h10408000;
      32328: inst = 32'hc404779;
      32329: inst = 32'h8220000;
      32330: inst = 32'h10408000;
      32331: inst = 32'hc40477a;
      32332: inst = 32'h8220000;
      32333: inst = 32'h10408000;
      32334: inst = 32'hc40477b;
      32335: inst = 32'h8220000;
      32336: inst = 32'h10408000;
      32337: inst = 32'hc40477c;
      32338: inst = 32'h8220000;
      32339: inst = 32'h10408000;
      32340: inst = 32'hc40477d;
      32341: inst = 32'h8220000;
      32342: inst = 32'h10408000;
      32343: inst = 32'hc40477e;
      32344: inst = 32'h8220000;
      32345: inst = 32'h10408000;
      32346: inst = 32'hc40477f;
      32347: inst = 32'h8220000;
      32348: inst = 32'h10408000;
      32349: inst = 32'hc404780;
      32350: inst = 32'h8220000;
      32351: inst = 32'h10408000;
      32352: inst = 32'hc404781;
      32353: inst = 32'h8220000;
      32354: inst = 32'h10408000;
      32355: inst = 32'hc404782;
      32356: inst = 32'h8220000;
      32357: inst = 32'h10408000;
      32358: inst = 32'hc404783;
      32359: inst = 32'h8220000;
      32360: inst = 32'h10408000;
      32361: inst = 32'hc404784;
      32362: inst = 32'h8220000;
      32363: inst = 32'h10408000;
      32364: inst = 32'hc404785;
      32365: inst = 32'h8220000;
      32366: inst = 32'h10408000;
      32367: inst = 32'hc404786;
      32368: inst = 32'h8220000;
      32369: inst = 32'h10408000;
      32370: inst = 32'hc404787;
      32371: inst = 32'h8220000;
      32372: inst = 32'h10408000;
      32373: inst = 32'hc404788;
      32374: inst = 32'h8220000;
      32375: inst = 32'h10408000;
      32376: inst = 32'hc404789;
      32377: inst = 32'h8220000;
      32378: inst = 32'h10408000;
      32379: inst = 32'hc40478a;
      32380: inst = 32'h8220000;
      32381: inst = 32'h10408000;
      32382: inst = 32'hc404795;
      32383: inst = 32'h8220000;
      32384: inst = 32'h10408000;
      32385: inst = 32'hc404796;
      32386: inst = 32'h8220000;
      32387: inst = 32'h10408000;
      32388: inst = 32'hc404797;
      32389: inst = 32'h8220000;
      32390: inst = 32'h10408000;
      32391: inst = 32'hc404799;
      32392: inst = 32'h8220000;
      32393: inst = 32'h10408000;
      32394: inst = 32'hc40479a;
      32395: inst = 32'h8220000;
      32396: inst = 32'h10408000;
      32397: inst = 32'hc40479b;
      32398: inst = 32'h8220000;
      32399: inst = 32'h10408000;
      32400: inst = 32'hc40479c;
      32401: inst = 32'h8220000;
      32402: inst = 32'h10408000;
      32403: inst = 32'hc40479d;
      32404: inst = 32'h8220000;
      32405: inst = 32'h10408000;
      32406: inst = 32'hc40479e;
      32407: inst = 32'h8220000;
      32408: inst = 32'h10408000;
      32409: inst = 32'hc40479f;
      32410: inst = 32'h8220000;
      32411: inst = 32'h10408000;
      32412: inst = 32'hc4047a0;
      32413: inst = 32'h8220000;
      32414: inst = 32'h10408000;
      32415: inst = 32'hc4047a1;
      32416: inst = 32'h8220000;
      32417: inst = 32'h10408000;
      32418: inst = 32'hc4047a2;
      32419: inst = 32'h8220000;
      32420: inst = 32'h10408000;
      32421: inst = 32'hc4047a3;
      32422: inst = 32'h8220000;
      32423: inst = 32'h10408000;
      32424: inst = 32'hc4047a4;
      32425: inst = 32'h8220000;
      32426: inst = 32'h10408000;
      32427: inst = 32'hc4047a5;
      32428: inst = 32'h8220000;
      32429: inst = 32'h10408000;
      32430: inst = 32'hc4047a6;
      32431: inst = 32'h8220000;
      32432: inst = 32'h10408000;
      32433: inst = 32'hc4047a7;
      32434: inst = 32'h8220000;
      32435: inst = 32'h10408000;
      32436: inst = 32'hc4047a8;
      32437: inst = 32'h8220000;
      32438: inst = 32'h10408000;
      32439: inst = 32'hc4047a9;
      32440: inst = 32'h8220000;
      32441: inst = 32'h10408000;
      32442: inst = 32'hc4047aa;
      32443: inst = 32'h8220000;
      32444: inst = 32'h10408000;
      32445: inst = 32'hc4047ab;
      32446: inst = 32'h8220000;
      32447: inst = 32'h10408000;
      32448: inst = 32'hc4047af;
      32449: inst = 32'h8220000;
      32450: inst = 32'h10408000;
      32451: inst = 32'hc4047b0;
      32452: inst = 32'h8220000;
      32453: inst = 32'h10408000;
      32454: inst = 32'hc4047b1;
      32455: inst = 32'h8220000;
      32456: inst = 32'h10408000;
      32457: inst = 32'hc4047b2;
      32458: inst = 32'h8220000;
      32459: inst = 32'h10408000;
      32460: inst = 32'hc4047b3;
      32461: inst = 32'h8220000;
      32462: inst = 32'h10408000;
      32463: inst = 32'hc4047b4;
      32464: inst = 32'h8220000;
      32465: inst = 32'h10408000;
      32466: inst = 32'hc4047b5;
      32467: inst = 32'h8220000;
      32468: inst = 32'h10408000;
      32469: inst = 32'hc4047b6;
      32470: inst = 32'h8220000;
      32471: inst = 32'h10408000;
      32472: inst = 32'hc4047b7;
      32473: inst = 32'h8220000;
      32474: inst = 32'h10408000;
      32475: inst = 32'hc4047b8;
      32476: inst = 32'h8220000;
      32477: inst = 32'h10408000;
      32478: inst = 32'hc4047b9;
      32479: inst = 32'h8220000;
      32480: inst = 32'h10408000;
      32481: inst = 32'hc4047ba;
      32482: inst = 32'h8220000;
      32483: inst = 32'h10408000;
      32484: inst = 32'hc4047bb;
      32485: inst = 32'h8220000;
      32486: inst = 32'h10408000;
      32487: inst = 32'hc4047bc;
      32488: inst = 32'h8220000;
      32489: inst = 32'h10408000;
      32490: inst = 32'hc4047c3;
      32491: inst = 32'h8220000;
      32492: inst = 32'h10408000;
      32493: inst = 32'hc4047c4;
      32494: inst = 32'h8220000;
      32495: inst = 32'h10408000;
      32496: inst = 32'hc4047c5;
      32497: inst = 32'h8220000;
      32498: inst = 32'h10408000;
      32499: inst = 32'hc4047c6;
      32500: inst = 32'h8220000;
      32501: inst = 32'h10408000;
      32502: inst = 32'hc4047c7;
      32503: inst = 32'h8220000;
      32504: inst = 32'h10408000;
      32505: inst = 32'hc4047c8;
      32506: inst = 32'h8220000;
      32507: inst = 32'h10408000;
      32508: inst = 32'hc4047c9;
      32509: inst = 32'h8220000;
      32510: inst = 32'h10408000;
      32511: inst = 32'hc4047ca;
      32512: inst = 32'h8220000;
      32513: inst = 32'h10408000;
      32514: inst = 32'hc4047cb;
      32515: inst = 32'h8220000;
      32516: inst = 32'h10408000;
      32517: inst = 32'hc4047cc;
      32518: inst = 32'h8220000;
      32519: inst = 32'h10408000;
      32520: inst = 32'hc4047cd;
      32521: inst = 32'h8220000;
      32522: inst = 32'h10408000;
      32523: inst = 32'hc4047d1;
      32524: inst = 32'h8220000;
      32525: inst = 32'h10408000;
      32526: inst = 32'hc4047d2;
      32527: inst = 32'h8220000;
      32528: inst = 32'h10408000;
      32529: inst = 32'hc4047d3;
      32530: inst = 32'h8220000;
      32531: inst = 32'h10408000;
      32532: inst = 32'hc4047d4;
      32533: inst = 32'h8220000;
      32534: inst = 32'h10408000;
      32535: inst = 32'hc4047d5;
      32536: inst = 32'h8220000;
      32537: inst = 32'h10408000;
      32538: inst = 32'hc4047d6;
      32539: inst = 32'h8220000;
      32540: inst = 32'h10408000;
      32541: inst = 32'hc4047d7;
      32542: inst = 32'h8220000;
      32543: inst = 32'h10408000;
      32544: inst = 32'hc4047d8;
      32545: inst = 32'h8220000;
      32546: inst = 32'h10408000;
      32547: inst = 32'hc4047d9;
      32548: inst = 32'h8220000;
      32549: inst = 32'h10408000;
      32550: inst = 32'hc4047da;
      32551: inst = 32'h8220000;
      32552: inst = 32'h10408000;
      32553: inst = 32'hc4047db;
      32554: inst = 32'h8220000;
      32555: inst = 32'h10408000;
      32556: inst = 32'hc4047dc;
      32557: inst = 32'h8220000;
      32558: inst = 32'h10408000;
      32559: inst = 32'hc4047dd;
      32560: inst = 32'h8220000;
      32561: inst = 32'h10408000;
      32562: inst = 32'hc4047de;
      32563: inst = 32'h8220000;
      32564: inst = 32'h10408000;
      32565: inst = 32'hc4047df;
      32566: inst = 32'h8220000;
      32567: inst = 32'h10408000;
      32568: inst = 32'hc4047e0;
      32569: inst = 32'h8220000;
      32570: inst = 32'h10408000;
      32571: inst = 32'hc4047e1;
      32572: inst = 32'h8220000;
      32573: inst = 32'h10408000;
      32574: inst = 32'hc4047e2;
      32575: inst = 32'h8220000;
      32576: inst = 32'h10408000;
      32577: inst = 32'hc4047e3;
      32578: inst = 32'h8220000;
      32579: inst = 32'h10408000;
      32580: inst = 32'hc4047e4;
      32581: inst = 32'h8220000;
      32582: inst = 32'h10408000;
      32583: inst = 32'hc4047e5;
      32584: inst = 32'h8220000;
      32585: inst = 32'h10408000;
      32586: inst = 32'hc4047e6;
      32587: inst = 32'h8220000;
      32588: inst = 32'h10408000;
      32589: inst = 32'hc4047e7;
      32590: inst = 32'h8220000;
      32591: inst = 32'h10408000;
      32592: inst = 32'hc4047e8;
      32593: inst = 32'h8220000;
      32594: inst = 32'h10408000;
      32595: inst = 32'hc4047e9;
      32596: inst = 32'h8220000;
      32597: inst = 32'h10408000;
      32598: inst = 32'hc4047ea;
      32599: inst = 32'h8220000;
      32600: inst = 32'h10408000;
      32601: inst = 32'hc4047ee;
      32602: inst = 32'h8220000;
      32603: inst = 32'h10408000;
      32604: inst = 32'hc4047ef;
      32605: inst = 32'h8220000;
      32606: inst = 32'h10408000;
      32607: inst = 32'hc4047f6;
      32608: inst = 32'h8220000;
      32609: inst = 32'h10408000;
      32610: inst = 32'hc4047f7;
      32611: inst = 32'h8220000;
      32612: inst = 32'h10408000;
      32613: inst = 32'hc4047fa;
      32614: inst = 32'h8220000;
      32615: inst = 32'h10408000;
      32616: inst = 32'hc4047fb;
      32617: inst = 32'h8220000;
      32618: inst = 32'h10408000;
      32619: inst = 32'hc4047fc;
      32620: inst = 32'h8220000;
      32621: inst = 32'h10408000;
      32622: inst = 32'hc4047fd;
      32623: inst = 32'h8220000;
      32624: inst = 32'h10408000;
      32625: inst = 32'hc4047fe;
      32626: inst = 32'h8220000;
      32627: inst = 32'h10408000;
      32628: inst = 32'hc4047ff;
      32629: inst = 32'h8220000;
      32630: inst = 32'h10408000;
      32631: inst = 32'hc404800;
      32632: inst = 32'h8220000;
      32633: inst = 32'h10408000;
      32634: inst = 32'hc404801;
      32635: inst = 32'h8220000;
      32636: inst = 32'h10408000;
      32637: inst = 32'hc404802;
      32638: inst = 32'h8220000;
      32639: inst = 32'h10408000;
      32640: inst = 32'hc404803;
      32641: inst = 32'h8220000;
      32642: inst = 32'h10408000;
      32643: inst = 32'hc404804;
      32644: inst = 32'h8220000;
      32645: inst = 32'h10408000;
      32646: inst = 32'hc404805;
      32647: inst = 32'h8220000;
      32648: inst = 32'h10408000;
      32649: inst = 32'hc404806;
      32650: inst = 32'h8220000;
      32651: inst = 32'h10408000;
      32652: inst = 32'hc404807;
      32653: inst = 32'h8220000;
      32654: inst = 32'h10408000;
      32655: inst = 32'hc404808;
      32656: inst = 32'h8220000;
      32657: inst = 32'h10408000;
      32658: inst = 32'hc404809;
      32659: inst = 32'h8220000;
      32660: inst = 32'h10408000;
      32661: inst = 32'hc40480a;
      32662: inst = 32'h8220000;
      32663: inst = 32'h10408000;
      32664: inst = 32'hc40480b;
      32665: inst = 32'h8220000;
      32666: inst = 32'h10408000;
      32667: inst = 32'hc40480f;
      32668: inst = 32'h8220000;
      32669: inst = 32'h10408000;
      32670: inst = 32'hc404810;
      32671: inst = 32'h8220000;
      32672: inst = 32'h10408000;
      32673: inst = 32'hc404811;
      32674: inst = 32'h8220000;
      32675: inst = 32'h10408000;
      32676: inst = 32'hc404812;
      32677: inst = 32'h8220000;
      32678: inst = 32'h10408000;
      32679: inst = 32'hc404813;
      32680: inst = 32'h8220000;
      32681: inst = 32'h10408000;
      32682: inst = 32'hc404814;
      32683: inst = 32'h8220000;
      32684: inst = 32'h10408000;
      32685: inst = 32'hc404815;
      32686: inst = 32'h8220000;
      32687: inst = 32'h10408000;
      32688: inst = 32'hc404816;
      32689: inst = 32'h8220000;
      32690: inst = 32'h10408000;
      32691: inst = 32'hc404817;
      32692: inst = 32'h8220000;
      32693: inst = 32'h10408000;
      32694: inst = 32'hc404818;
      32695: inst = 32'h8220000;
      32696: inst = 32'h10408000;
      32697: inst = 32'hc404819;
      32698: inst = 32'h8220000;
      32699: inst = 32'h10408000;
      32700: inst = 32'hc40481a;
      32701: inst = 32'h8220000;
      32702: inst = 32'h10408000;
      32703: inst = 32'hc40481b;
      32704: inst = 32'h8220000;
      32705: inst = 32'h10408000;
      32706: inst = 32'hc40481c;
      32707: inst = 32'h8220000;
      32708: inst = 32'h10408000;
      32709: inst = 32'hc404823;
      32710: inst = 32'h8220000;
      32711: inst = 32'h10408000;
      32712: inst = 32'hc404824;
      32713: inst = 32'h8220000;
      32714: inst = 32'h10408000;
      32715: inst = 32'hc404825;
      32716: inst = 32'h8220000;
      32717: inst = 32'h10408000;
      32718: inst = 32'hc404826;
      32719: inst = 32'h8220000;
      32720: inst = 32'h10408000;
      32721: inst = 32'hc404827;
      32722: inst = 32'h8220000;
      32723: inst = 32'h10408000;
      32724: inst = 32'hc404828;
      32725: inst = 32'h8220000;
      32726: inst = 32'h10408000;
      32727: inst = 32'hc404829;
      32728: inst = 32'h8220000;
      32729: inst = 32'h10408000;
      32730: inst = 32'hc40482a;
      32731: inst = 32'h8220000;
      32732: inst = 32'h10408000;
      32733: inst = 32'hc40482b;
      32734: inst = 32'h8220000;
      32735: inst = 32'h10408000;
      32736: inst = 32'hc40482c;
      32737: inst = 32'h8220000;
      32738: inst = 32'h10408000;
      32739: inst = 32'hc40482d;
      32740: inst = 32'h8220000;
      32741: inst = 32'h10408000;
      32742: inst = 32'hc404831;
      32743: inst = 32'h8220000;
      32744: inst = 32'h10408000;
      32745: inst = 32'hc404832;
      32746: inst = 32'h8220000;
      32747: inst = 32'h10408000;
      32748: inst = 32'hc404833;
      32749: inst = 32'h8220000;
      32750: inst = 32'h10408000;
      32751: inst = 32'hc404834;
      32752: inst = 32'h8220000;
      32753: inst = 32'h10408000;
      32754: inst = 32'hc404835;
      32755: inst = 32'h8220000;
      32756: inst = 32'h10408000;
      32757: inst = 32'hc404836;
      32758: inst = 32'h8220000;
      32759: inst = 32'h10408000;
      32760: inst = 32'hc404837;
      32761: inst = 32'h8220000;
      32762: inst = 32'h10408000;
      32763: inst = 32'hc404838;
      32764: inst = 32'h8220000;
      32765: inst = 32'h10408000;
      32766: inst = 32'hc404839;
      32767: inst = 32'h8220000;
      32768: inst = 32'h10408000;
      32769: inst = 32'hc40483a;
      32770: inst = 32'h8220000;
      32771: inst = 32'h10408000;
      32772: inst = 32'hc40483b;
      32773: inst = 32'h8220000;
      32774: inst = 32'h10408000;
      32775: inst = 32'hc40483c;
      32776: inst = 32'h8220000;
      32777: inst = 32'h10408000;
      32778: inst = 32'hc40483d;
      32779: inst = 32'h8220000;
      32780: inst = 32'h10408000;
      32781: inst = 32'hc40483e;
      32782: inst = 32'h8220000;
      32783: inst = 32'h10408000;
      32784: inst = 32'hc40483f;
      32785: inst = 32'h8220000;
      32786: inst = 32'h10408000;
      32787: inst = 32'hc404840;
      32788: inst = 32'h8220000;
      32789: inst = 32'h10408000;
      32790: inst = 32'hc404841;
      32791: inst = 32'h8220000;
      32792: inst = 32'h10408000;
      32793: inst = 32'hc404842;
      32794: inst = 32'h8220000;
      32795: inst = 32'h10408000;
      32796: inst = 32'hc404843;
      32797: inst = 32'h8220000;
      32798: inst = 32'h10408000;
      32799: inst = 32'hc404844;
      32800: inst = 32'h8220000;
      32801: inst = 32'h10408000;
      32802: inst = 32'hc404845;
      32803: inst = 32'h8220000;
      32804: inst = 32'h10408000;
      32805: inst = 32'hc404846;
      32806: inst = 32'h8220000;
      32807: inst = 32'h10408000;
      32808: inst = 32'hc404847;
      32809: inst = 32'h8220000;
      32810: inst = 32'h10408000;
      32811: inst = 32'hc404848;
      32812: inst = 32'h8220000;
      32813: inst = 32'h10408000;
      32814: inst = 32'hc404849;
      32815: inst = 32'h8220000;
      32816: inst = 32'h10408000;
      32817: inst = 32'hc40484a;
      32818: inst = 32'h8220000;
      32819: inst = 32'h10408000;
      32820: inst = 32'hc40484b;
      32821: inst = 32'h8220000;
      32822: inst = 32'h10408000;
      32823: inst = 32'hc40484c;
      32824: inst = 32'h8220000;
      32825: inst = 32'h10408000;
      32826: inst = 32'hc40484d;
      32827: inst = 32'h8220000;
      32828: inst = 32'h10408000;
      32829: inst = 32'hc40484e;
      32830: inst = 32'h8220000;
      32831: inst = 32'h10408000;
      32832: inst = 32'hc40484f;
      32833: inst = 32'h8220000;
      32834: inst = 32'h10408000;
      32835: inst = 32'hc404850;
      32836: inst = 32'h8220000;
      32837: inst = 32'h10408000;
      32838: inst = 32'hc404851;
      32839: inst = 32'h8220000;
      32840: inst = 32'h10408000;
      32841: inst = 32'hc404852;
      32842: inst = 32'h8220000;
      32843: inst = 32'h10408000;
      32844: inst = 32'hc404853;
      32845: inst = 32'h8220000;
      32846: inst = 32'h10408000;
      32847: inst = 32'hc40485a;
      32848: inst = 32'h8220000;
      32849: inst = 32'h10408000;
      32850: inst = 32'hc40485b;
      32851: inst = 32'h8220000;
      32852: inst = 32'h10408000;
      32853: inst = 32'hc40485c;
      32854: inst = 32'h8220000;
      32855: inst = 32'h10408000;
      32856: inst = 32'hc40485d;
      32857: inst = 32'h8220000;
      32858: inst = 32'h10408000;
      32859: inst = 32'hc40485e;
      32860: inst = 32'h8220000;
      32861: inst = 32'h10408000;
      32862: inst = 32'hc40485f;
      32863: inst = 32'h8220000;
      32864: inst = 32'h10408000;
      32865: inst = 32'hc404860;
      32866: inst = 32'h8220000;
      32867: inst = 32'h10408000;
      32868: inst = 32'hc404861;
      32869: inst = 32'h8220000;
      32870: inst = 32'h10408000;
      32871: inst = 32'hc404862;
      32872: inst = 32'h8220000;
      32873: inst = 32'h10408000;
      32874: inst = 32'hc404863;
      32875: inst = 32'h8220000;
      32876: inst = 32'h10408000;
      32877: inst = 32'hc404864;
      32878: inst = 32'h8220000;
      32879: inst = 32'h10408000;
      32880: inst = 32'hc404865;
      32881: inst = 32'h8220000;
      32882: inst = 32'h10408000;
      32883: inst = 32'hc404866;
      32884: inst = 32'h8220000;
      32885: inst = 32'h10408000;
      32886: inst = 32'hc404867;
      32887: inst = 32'h8220000;
      32888: inst = 32'h10408000;
      32889: inst = 32'hc404868;
      32890: inst = 32'h8220000;
      32891: inst = 32'h10408000;
      32892: inst = 32'hc404869;
      32893: inst = 32'h8220000;
      32894: inst = 32'h10408000;
      32895: inst = 32'hc40486a;
      32896: inst = 32'h8220000;
      32897: inst = 32'h10408000;
      32898: inst = 32'hc40486b;
      32899: inst = 32'h8220000;
      32900: inst = 32'h10408000;
      32901: inst = 32'hc40486f;
      32902: inst = 32'h8220000;
      32903: inst = 32'h10408000;
      32904: inst = 32'hc404870;
      32905: inst = 32'h8220000;
      32906: inst = 32'h10408000;
      32907: inst = 32'hc404871;
      32908: inst = 32'h8220000;
      32909: inst = 32'h10408000;
      32910: inst = 32'hc404872;
      32911: inst = 32'h8220000;
      32912: inst = 32'h10408000;
      32913: inst = 32'hc404873;
      32914: inst = 32'h8220000;
      32915: inst = 32'h10408000;
      32916: inst = 32'hc404874;
      32917: inst = 32'h8220000;
      32918: inst = 32'h10408000;
      32919: inst = 32'hc404875;
      32920: inst = 32'h8220000;
      32921: inst = 32'h10408000;
      32922: inst = 32'hc404876;
      32923: inst = 32'h8220000;
      32924: inst = 32'h10408000;
      32925: inst = 32'hc404877;
      32926: inst = 32'h8220000;
      32927: inst = 32'h10408000;
      32928: inst = 32'hc404878;
      32929: inst = 32'h8220000;
      32930: inst = 32'h10408000;
      32931: inst = 32'hc404879;
      32932: inst = 32'h8220000;
      32933: inst = 32'h10408000;
      32934: inst = 32'hc40487a;
      32935: inst = 32'h8220000;
      32936: inst = 32'h10408000;
      32937: inst = 32'hc40487b;
      32938: inst = 32'h8220000;
      32939: inst = 32'h10408000;
      32940: inst = 32'hc40487c;
      32941: inst = 32'h8220000;
      32942: inst = 32'h10408000;
      32943: inst = 32'hc404883;
      32944: inst = 32'h8220000;
      32945: inst = 32'h10408000;
      32946: inst = 32'hc404884;
      32947: inst = 32'h8220000;
      32948: inst = 32'h10408000;
      32949: inst = 32'hc404885;
      32950: inst = 32'h8220000;
      32951: inst = 32'h10408000;
      32952: inst = 32'hc404886;
      32953: inst = 32'h8220000;
      32954: inst = 32'h10408000;
      32955: inst = 32'hc404887;
      32956: inst = 32'h8220000;
      32957: inst = 32'h10408000;
      32958: inst = 32'hc404888;
      32959: inst = 32'h8220000;
      32960: inst = 32'h10408000;
      32961: inst = 32'hc404889;
      32962: inst = 32'h8220000;
      32963: inst = 32'h10408000;
      32964: inst = 32'hc40488a;
      32965: inst = 32'h8220000;
      32966: inst = 32'h10408000;
      32967: inst = 32'hc40488b;
      32968: inst = 32'h8220000;
      32969: inst = 32'h10408000;
      32970: inst = 32'hc40488c;
      32971: inst = 32'h8220000;
      32972: inst = 32'h10408000;
      32973: inst = 32'hc40488d;
      32974: inst = 32'h8220000;
      32975: inst = 32'h10408000;
      32976: inst = 32'hc404891;
      32977: inst = 32'h8220000;
      32978: inst = 32'h10408000;
      32979: inst = 32'hc404892;
      32980: inst = 32'h8220000;
      32981: inst = 32'h10408000;
      32982: inst = 32'hc404893;
      32983: inst = 32'h8220000;
      32984: inst = 32'h10408000;
      32985: inst = 32'hc404894;
      32986: inst = 32'h8220000;
      32987: inst = 32'h10408000;
      32988: inst = 32'hc404895;
      32989: inst = 32'h8220000;
      32990: inst = 32'h10408000;
      32991: inst = 32'hc404896;
      32992: inst = 32'h8220000;
      32993: inst = 32'h10408000;
      32994: inst = 32'hc404897;
      32995: inst = 32'h8220000;
      32996: inst = 32'h10408000;
      32997: inst = 32'hc404898;
      32998: inst = 32'h8220000;
      32999: inst = 32'h10408000;
      33000: inst = 32'hc404899;
      33001: inst = 32'h8220000;
      33002: inst = 32'h10408000;
      33003: inst = 32'hc40489a;
      33004: inst = 32'h8220000;
      33005: inst = 32'h10408000;
      33006: inst = 32'hc40489b;
      33007: inst = 32'h8220000;
      33008: inst = 32'h10408000;
      33009: inst = 32'hc40489c;
      33010: inst = 32'h8220000;
      33011: inst = 32'h10408000;
      33012: inst = 32'hc40489d;
      33013: inst = 32'h8220000;
      33014: inst = 32'h10408000;
      33015: inst = 32'hc40489e;
      33016: inst = 32'h8220000;
      33017: inst = 32'h10408000;
      33018: inst = 32'hc40489f;
      33019: inst = 32'h8220000;
      33020: inst = 32'h10408000;
      33021: inst = 32'hc4048a0;
      33022: inst = 32'h8220000;
      33023: inst = 32'h10408000;
      33024: inst = 32'hc4048a1;
      33025: inst = 32'h8220000;
      33026: inst = 32'h10408000;
      33027: inst = 32'hc4048a2;
      33028: inst = 32'h8220000;
      33029: inst = 32'h10408000;
      33030: inst = 32'hc4048a3;
      33031: inst = 32'h8220000;
      33032: inst = 32'h10408000;
      33033: inst = 32'hc4048a4;
      33034: inst = 32'h8220000;
      33035: inst = 32'h10408000;
      33036: inst = 32'hc4048a5;
      33037: inst = 32'h8220000;
      33038: inst = 32'h10408000;
      33039: inst = 32'hc4048a6;
      33040: inst = 32'h8220000;
      33041: inst = 32'h10408000;
      33042: inst = 32'hc4048a7;
      33043: inst = 32'h8220000;
      33044: inst = 32'h10408000;
      33045: inst = 32'hc4048a8;
      33046: inst = 32'h8220000;
      33047: inst = 32'h10408000;
      33048: inst = 32'hc4048a9;
      33049: inst = 32'h8220000;
      33050: inst = 32'h10408000;
      33051: inst = 32'hc4048aa;
      33052: inst = 32'h8220000;
      33053: inst = 32'h10408000;
      33054: inst = 32'hc4048ab;
      33055: inst = 32'h8220000;
      33056: inst = 32'h10408000;
      33057: inst = 32'hc4048ac;
      33058: inst = 32'h8220000;
      33059: inst = 32'h10408000;
      33060: inst = 32'hc4048ad;
      33061: inst = 32'h8220000;
      33062: inst = 32'h10408000;
      33063: inst = 32'hc4048ae;
      33064: inst = 32'h8220000;
      33065: inst = 32'h10408000;
      33066: inst = 32'hc4048af;
      33067: inst = 32'h8220000;
      33068: inst = 32'h10408000;
      33069: inst = 32'hc4048b0;
      33070: inst = 32'h8220000;
      33071: inst = 32'h10408000;
      33072: inst = 32'hc4048b1;
      33073: inst = 32'h8220000;
      33074: inst = 32'h10408000;
      33075: inst = 32'hc4048b2;
      33076: inst = 32'h8220000;
      33077: inst = 32'h10408000;
      33078: inst = 32'hc4048b3;
      33079: inst = 32'h8220000;
      33080: inst = 32'h10408000;
      33081: inst = 32'hc4048ba;
      33082: inst = 32'h8220000;
      33083: inst = 32'h10408000;
      33084: inst = 32'hc4048bb;
      33085: inst = 32'h8220000;
      33086: inst = 32'h10408000;
      33087: inst = 32'hc4048bc;
      33088: inst = 32'h8220000;
      33089: inst = 32'h10408000;
      33090: inst = 32'hc4048bd;
      33091: inst = 32'h8220000;
      33092: inst = 32'h10408000;
      33093: inst = 32'hc4048be;
      33094: inst = 32'h8220000;
      33095: inst = 32'h10408000;
      33096: inst = 32'hc4048bf;
      33097: inst = 32'h8220000;
      33098: inst = 32'h10408000;
      33099: inst = 32'hc4048c0;
      33100: inst = 32'h8220000;
      33101: inst = 32'h10408000;
      33102: inst = 32'hc4048c1;
      33103: inst = 32'h8220000;
      33104: inst = 32'h10408000;
      33105: inst = 32'hc4048c2;
      33106: inst = 32'h8220000;
      33107: inst = 32'h10408000;
      33108: inst = 32'hc4048c3;
      33109: inst = 32'h8220000;
      33110: inst = 32'h10408000;
      33111: inst = 32'hc4048c4;
      33112: inst = 32'h8220000;
      33113: inst = 32'h10408000;
      33114: inst = 32'hc4048c5;
      33115: inst = 32'h8220000;
      33116: inst = 32'h10408000;
      33117: inst = 32'hc4048c6;
      33118: inst = 32'h8220000;
      33119: inst = 32'h10408000;
      33120: inst = 32'hc4048c7;
      33121: inst = 32'h8220000;
      33122: inst = 32'h10408000;
      33123: inst = 32'hc4048c8;
      33124: inst = 32'h8220000;
      33125: inst = 32'h10408000;
      33126: inst = 32'hc4048c9;
      33127: inst = 32'h8220000;
      33128: inst = 32'h10408000;
      33129: inst = 32'hc4048ca;
      33130: inst = 32'h8220000;
      33131: inst = 32'h10408000;
      33132: inst = 32'hc4048cb;
      33133: inst = 32'h8220000;
      33134: inst = 32'h10408000;
      33135: inst = 32'hc4048cf;
      33136: inst = 32'h8220000;
      33137: inst = 32'h10408000;
      33138: inst = 32'hc4048d0;
      33139: inst = 32'h8220000;
      33140: inst = 32'h10408000;
      33141: inst = 32'hc4048d1;
      33142: inst = 32'h8220000;
      33143: inst = 32'h10408000;
      33144: inst = 32'hc4048d2;
      33145: inst = 32'h8220000;
      33146: inst = 32'h10408000;
      33147: inst = 32'hc4048d3;
      33148: inst = 32'h8220000;
      33149: inst = 32'h10408000;
      33150: inst = 32'hc4048d4;
      33151: inst = 32'h8220000;
      33152: inst = 32'h10408000;
      33153: inst = 32'hc4048d5;
      33154: inst = 32'h8220000;
      33155: inst = 32'h10408000;
      33156: inst = 32'hc4048d6;
      33157: inst = 32'h8220000;
      33158: inst = 32'h10408000;
      33159: inst = 32'hc4048d7;
      33160: inst = 32'h8220000;
      33161: inst = 32'h10408000;
      33162: inst = 32'hc4048d8;
      33163: inst = 32'h8220000;
      33164: inst = 32'h10408000;
      33165: inst = 32'hc4048d9;
      33166: inst = 32'h8220000;
      33167: inst = 32'h10408000;
      33168: inst = 32'hc4048da;
      33169: inst = 32'h8220000;
      33170: inst = 32'h10408000;
      33171: inst = 32'hc4048db;
      33172: inst = 32'h8220000;
      33173: inst = 32'h10408000;
      33174: inst = 32'hc4048dc;
      33175: inst = 32'h8220000;
      33176: inst = 32'h10408000;
      33177: inst = 32'hc4048e3;
      33178: inst = 32'h8220000;
      33179: inst = 32'h10408000;
      33180: inst = 32'hc4048e4;
      33181: inst = 32'h8220000;
      33182: inst = 32'h10408000;
      33183: inst = 32'hc4048e5;
      33184: inst = 32'h8220000;
      33185: inst = 32'h10408000;
      33186: inst = 32'hc4048e6;
      33187: inst = 32'h8220000;
      33188: inst = 32'h10408000;
      33189: inst = 32'hc4048e7;
      33190: inst = 32'h8220000;
      33191: inst = 32'h10408000;
      33192: inst = 32'hc4048e8;
      33193: inst = 32'h8220000;
      33194: inst = 32'h10408000;
      33195: inst = 32'hc4048e9;
      33196: inst = 32'h8220000;
      33197: inst = 32'h10408000;
      33198: inst = 32'hc4048ea;
      33199: inst = 32'h8220000;
      33200: inst = 32'h10408000;
      33201: inst = 32'hc4048eb;
      33202: inst = 32'h8220000;
      33203: inst = 32'h10408000;
      33204: inst = 32'hc4048ec;
      33205: inst = 32'h8220000;
      33206: inst = 32'h10408000;
      33207: inst = 32'hc4048ed;
      33208: inst = 32'h8220000;
      33209: inst = 32'h10408000;
      33210: inst = 32'hc4048f1;
      33211: inst = 32'h8220000;
      33212: inst = 32'h10408000;
      33213: inst = 32'hc4048f2;
      33214: inst = 32'h8220000;
      33215: inst = 32'h10408000;
      33216: inst = 32'hc4048f3;
      33217: inst = 32'h8220000;
      33218: inst = 32'h10408000;
      33219: inst = 32'hc4048f4;
      33220: inst = 32'h8220000;
      33221: inst = 32'h10408000;
      33222: inst = 32'hc4048f5;
      33223: inst = 32'h8220000;
      33224: inst = 32'h10408000;
      33225: inst = 32'hc4048f6;
      33226: inst = 32'h8220000;
      33227: inst = 32'h10408000;
      33228: inst = 32'hc4048f7;
      33229: inst = 32'h8220000;
      33230: inst = 32'h10408000;
      33231: inst = 32'hc4048f8;
      33232: inst = 32'h8220000;
      33233: inst = 32'h10408000;
      33234: inst = 32'hc4048f9;
      33235: inst = 32'h8220000;
      33236: inst = 32'h10408000;
      33237: inst = 32'hc4048fa;
      33238: inst = 32'h8220000;
      33239: inst = 32'h10408000;
      33240: inst = 32'hc4048fb;
      33241: inst = 32'h8220000;
      33242: inst = 32'h10408000;
      33243: inst = 32'hc4048fc;
      33244: inst = 32'h8220000;
      33245: inst = 32'h10408000;
      33246: inst = 32'hc4048fd;
      33247: inst = 32'h8220000;
      33248: inst = 32'h10408000;
      33249: inst = 32'hc4048fe;
      33250: inst = 32'h8220000;
      33251: inst = 32'h10408000;
      33252: inst = 32'hc4048ff;
      33253: inst = 32'h8220000;
      33254: inst = 32'h10408000;
      33255: inst = 32'hc404900;
      33256: inst = 32'h8220000;
      33257: inst = 32'h10408000;
      33258: inst = 32'hc404901;
      33259: inst = 32'h8220000;
      33260: inst = 32'h10408000;
      33261: inst = 32'hc404902;
      33262: inst = 32'h8220000;
      33263: inst = 32'h10408000;
      33264: inst = 32'hc404903;
      33265: inst = 32'h8220000;
      33266: inst = 32'h10408000;
      33267: inst = 32'hc404904;
      33268: inst = 32'h8220000;
      33269: inst = 32'h10408000;
      33270: inst = 32'hc404905;
      33271: inst = 32'h8220000;
      33272: inst = 32'h10408000;
      33273: inst = 32'hc404906;
      33274: inst = 32'h8220000;
      33275: inst = 32'h10408000;
      33276: inst = 32'hc404907;
      33277: inst = 32'h8220000;
      33278: inst = 32'h10408000;
      33279: inst = 32'hc404908;
      33280: inst = 32'h8220000;
      33281: inst = 32'h10408000;
      33282: inst = 32'hc404909;
      33283: inst = 32'h8220000;
      33284: inst = 32'h10408000;
      33285: inst = 32'hc40490a;
      33286: inst = 32'h8220000;
      33287: inst = 32'h10408000;
      33288: inst = 32'hc40490b;
      33289: inst = 32'h8220000;
      33290: inst = 32'h10408000;
      33291: inst = 32'hc40490c;
      33292: inst = 32'h8220000;
      33293: inst = 32'h10408000;
      33294: inst = 32'hc40490d;
      33295: inst = 32'h8220000;
      33296: inst = 32'h10408000;
      33297: inst = 32'hc40490e;
      33298: inst = 32'h8220000;
      33299: inst = 32'h10408000;
      33300: inst = 32'hc40490f;
      33301: inst = 32'h8220000;
      33302: inst = 32'h10408000;
      33303: inst = 32'hc404910;
      33304: inst = 32'h8220000;
      33305: inst = 32'h10408000;
      33306: inst = 32'hc404911;
      33307: inst = 32'h8220000;
      33308: inst = 32'h10408000;
      33309: inst = 32'hc404912;
      33310: inst = 32'h8220000;
      33311: inst = 32'h10408000;
      33312: inst = 32'hc404913;
      33313: inst = 32'h8220000;
      33314: inst = 32'h10408000;
      33315: inst = 32'hc404916;
      33316: inst = 32'h8220000;
      33317: inst = 32'h10408000;
      33318: inst = 32'hc40491a;
      33319: inst = 32'h8220000;
      33320: inst = 32'h10408000;
      33321: inst = 32'hc40491b;
      33322: inst = 32'h8220000;
      33323: inst = 32'h10408000;
      33324: inst = 32'hc40491c;
      33325: inst = 32'h8220000;
      33326: inst = 32'h10408000;
      33327: inst = 32'hc40491d;
      33328: inst = 32'h8220000;
      33329: inst = 32'h10408000;
      33330: inst = 32'hc40491e;
      33331: inst = 32'h8220000;
      33332: inst = 32'h10408000;
      33333: inst = 32'hc40491f;
      33334: inst = 32'h8220000;
      33335: inst = 32'h10408000;
      33336: inst = 32'hc404920;
      33337: inst = 32'h8220000;
      33338: inst = 32'h10408000;
      33339: inst = 32'hc404921;
      33340: inst = 32'h8220000;
      33341: inst = 32'h10408000;
      33342: inst = 32'hc404922;
      33343: inst = 32'h8220000;
      33344: inst = 32'h10408000;
      33345: inst = 32'hc404923;
      33346: inst = 32'h8220000;
      33347: inst = 32'h10408000;
      33348: inst = 32'hc404924;
      33349: inst = 32'h8220000;
      33350: inst = 32'h10408000;
      33351: inst = 32'hc404925;
      33352: inst = 32'h8220000;
      33353: inst = 32'h10408000;
      33354: inst = 32'hc404926;
      33355: inst = 32'h8220000;
      33356: inst = 32'h10408000;
      33357: inst = 32'hc404927;
      33358: inst = 32'h8220000;
      33359: inst = 32'h10408000;
      33360: inst = 32'hc404928;
      33361: inst = 32'h8220000;
      33362: inst = 32'h10408000;
      33363: inst = 32'hc404929;
      33364: inst = 32'h8220000;
      33365: inst = 32'h10408000;
      33366: inst = 32'hc40492a;
      33367: inst = 32'h8220000;
      33368: inst = 32'h10408000;
      33369: inst = 32'hc40492b;
      33370: inst = 32'h8220000;
      33371: inst = 32'h10408000;
      33372: inst = 32'hc40492f;
      33373: inst = 32'h8220000;
      33374: inst = 32'h10408000;
      33375: inst = 32'hc404930;
      33376: inst = 32'h8220000;
      33377: inst = 32'h10408000;
      33378: inst = 32'hc404931;
      33379: inst = 32'h8220000;
      33380: inst = 32'h10408000;
      33381: inst = 32'hc404932;
      33382: inst = 32'h8220000;
      33383: inst = 32'h10408000;
      33384: inst = 32'hc404933;
      33385: inst = 32'h8220000;
      33386: inst = 32'h10408000;
      33387: inst = 32'hc404934;
      33388: inst = 32'h8220000;
      33389: inst = 32'h10408000;
      33390: inst = 32'hc404935;
      33391: inst = 32'h8220000;
      33392: inst = 32'h10408000;
      33393: inst = 32'hc404936;
      33394: inst = 32'h8220000;
      33395: inst = 32'h10408000;
      33396: inst = 32'hc404937;
      33397: inst = 32'h8220000;
      33398: inst = 32'h10408000;
      33399: inst = 32'hc404938;
      33400: inst = 32'h8220000;
      33401: inst = 32'h10408000;
      33402: inst = 32'hc404939;
      33403: inst = 32'h8220000;
      33404: inst = 32'h10408000;
      33405: inst = 32'hc40493a;
      33406: inst = 32'h8220000;
      33407: inst = 32'h10408000;
      33408: inst = 32'hc40493b;
      33409: inst = 32'h8220000;
      33410: inst = 32'h10408000;
      33411: inst = 32'hc40493c;
      33412: inst = 32'h8220000;
      33413: inst = 32'h10408000;
      33414: inst = 32'hc404943;
      33415: inst = 32'h8220000;
      33416: inst = 32'h10408000;
      33417: inst = 32'hc404944;
      33418: inst = 32'h8220000;
      33419: inst = 32'h10408000;
      33420: inst = 32'hc404945;
      33421: inst = 32'h8220000;
      33422: inst = 32'h10408000;
      33423: inst = 32'hc404946;
      33424: inst = 32'h8220000;
      33425: inst = 32'h10408000;
      33426: inst = 32'hc404947;
      33427: inst = 32'h8220000;
      33428: inst = 32'h10408000;
      33429: inst = 32'hc404948;
      33430: inst = 32'h8220000;
      33431: inst = 32'h10408000;
      33432: inst = 32'hc404949;
      33433: inst = 32'h8220000;
      33434: inst = 32'h10408000;
      33435: inst = 32'hc40494a;
      33436: inst = 32'h8220000;
      33437: inst = 32'h10408000;
      33438: inst = 32'hc40494b;
      33439: inst = 32'h8220000;
      33440: inst = 32'h10408000;
      33441: inst = 32'hc40494c;
      33442: inst = 32'h8220000;
      33443: inst = 32'h10408000;
      33444: inst = 32'hc40494d;
      33445: inst = 32'h8220000;
      33446: inst = 32'h10408000;
      33447: inst = 32'hc404951;
      33448: inst = 32'h8220000;
      33449: inst = 32'h10408000;
      33450: inst = 32'hc404952;
      33451: inst = 32'h8220000;
      33452: inst = 32'h10408000;
      33453: inst = 32'hc404953;
      33454: inst = 32'h8220000;
      33455: inst = 32'h10408000;
      33456: inst = 32'hc404954;
      33457: inst = 32'h8220000;
      33458: inst = 32'h10408000;
      33459: inst = 32'hc404955;
      33460: inst = 32'h8220000;
      33461: inst = 32'h10408000;
      33462: inst = 32'hc404956;
      33463: inst = 32'h8220000;
      33464: inst = 32'h10408000;
      33465: inst = 32'hc404957;
      33466: inst = 32'h8220000;
      33467: inst = 32'h10408000;
      33468: inst = 32'hc404958;
      33469: inst = 32'h8220000;
      33470: inst = 32'h10408000;
      33471: inst = 32'hc404959;
      33472: inst = 32'h8220000;
      33473: inst = 32'h10408000;
      33474: inst = 32'hc40495a;
      33475: inst = 32'h8220000;
      33476: inst = 32'h10408000;
      33477: inst = 32'hc40495b;
      33478: inst = 32'h8220000;
      33479: inst = 32'h10408000;
      33480: inst = 32'hc40495c;
      33481: inst = 32'h8220000;
      33482: inst = 32'h10408000;
      33483: inst = 32'hc40495d;
      33484: inst = 32'h8220000;
      33485: inst = 32'h10408000;
      33486: inst = 32'hc40495e;
      33487: inst = 32'h8220000;
      33488: inst = 32'h10408000;
      33489: inst = 32'hc40495f;
      33490: inst = 32'h8220000;
      33491: inst = 32'h10408000;
      33492: inst = 32'hc404960;
      33493: inst = 32'h8220000;
      33494: inst = 32'h10408000;
      33495: inst = 32'hc404961;
      33496: inst = 32'h8220000;
      33497: inst = 32'h10408000;
      33498: inst = 32'hc404962;
      33499: inst = 32'h8220000;
      33500: inst = 32'h10408000;
      33501: inst = 32'hc404963;
      33502: inst = 32'h8220000;
      33503: inst = 32'h10408000;
      33504: inst = 32'hc404964;
      33505: inst = 32'h8220000;
      33506: inst = 32'h10408000;
      33507: inst = 32'hc404965;
      33508: inst = 32'h8220000;
      33509: inst = 32'h10408000;
      33510: inst = 32'hc404966;
      33511: inst = 32'h8220000;
      33512: inst = 32'h10408000;
      33513: inst = 32'hc404967;
      33514: inst = 32'h8220000;
      33515: inst = 32'h10408000;
      33516: inst = 32'hc404968;
      33517: inst = 32'h8220000;
      33518: inst = 32'h10408000;
      33519: inst = 32'hc404969;
      33520: inst = 32'h8220000;
      33521: inst = 32'h10408000;
      33522: inst = 32'hc40496a;
      33523: inst = 32'h8220000;
      33524: inst = 32'h10408000;
      33525: inst = 32'hc40496b;
      33526: inst = 32'h8220000;
      33527: inst = 32'h10408000;
      33528: inst = 32'hc40496c;
      33529: inst = 32'h8220000;
      33530: inst = 32'h10408000;
      33531: inst = 32'hc40496d;
      33532: inst = 32'h8220000;
      33533: inst = 32'h10408000;
      33534: inst = 32'hc40496e;
      33535: inst = 32'h8220000;
      33536: inst = 32'h10408000;
      33537: inst = 32'hc40496f;
      33538: inst = 32'h8220000;
      33539: inst = 32'h10408000;
      33540: inst = 32'hc404970;
      33541: inst = 32'h8220000;
      33542: inst = 32'h10408000;
      33543: inst = 32'hc404971;
      33544: inst = 32'h8220000;
      33545: inst = 32'h10408000;
      33546: inst = 32'hc404972;
      33547: inst = 32'h8220000;
      33548: inst = 32'h10408000;
      33549: inst = 32'hc404973;
      33550: inst = 32'h8220000;
      33551: inst = 32'h10408000;
      33552: inst = 32'hc404974;
      33553: inst = 32'h8220000;
      33554: inst = 32'h10408000;
      33555: inst = 32'hc404975;
      33556: inst = 32'h8220000;
      33557: inst = 32'h10408000;
      33558: inst = 32'hc404976;
      33559: inst = 32'h8220000;
      33560: inst = 32'h10408000;
      33561: inst = 32'hc404977;
      33562: inst = 32'h8220000;
      33563: inst = 32'h10408000;
      33564: inst = 32'hc404978;
      33565: inst = 32'h8220000;
      33566: inst = 32'h10408000;
      33567: inst = 32'hc404979;
      33568: inst = 32'h8220000;
      33569: inst = 32'h10408000;
      33570: inst = 32'hc40497a;
      33571: inst = 32'h8220000;
      33572: inst = 32'h10408000;
      33573: inst = 32'hc40497b;
      33574: inst = 32'h8220000;
      33575: inst = 32'h10408000;
      33576: inst = 32'hc40497c;
      33577: inst = 32'h8220000;
      33578: inst = 32'h10408000;
      33579: inst = 32'hc40497d;
      33580: inst = 32'h8220000;
      33581: inst = 32'h10408000;
      33582: inst = 32'hc40497e;
      33583: inst = 32'h8220000;
      33584: inst = 32'h10408000;
      33585: inst = 32'hc40497f;
      33586: inst = 32'h8220000;
      33587: inst = 32'h10408000;
      33588: inst = 32'hc404980;
      33589: inst = 32'h8220000;
      33590: inst = 32'h10408000;
      33591: inst = 32'hc404981;
      33592: inst = 32'h8220000;
      33593: inst = 32'h10408000;
      33594: inst = 32'hc404982;
      33595: inst = 32'h8220000;
      33596: inst = 32'h10408000;
      33597: inst = 32'hc404983;
      33598: inst = 32'h8220000;
      33599: inst = 32'h10408000;
      33600: inst = 32'hc404984;
      33601: inst = 32'h8220000;
      33602: inst = 32'h10408000;
      33603: inst = 32'hc404985;
      33604: inst = 32'h8220000;
      33605: inst = 32'h10408000;
      33606: inst = 32'hc40498f;
      33607: inst = 32'h8220000;
      33608: inst = 32'h10408000;
      33609: inst = 32'hc404990;
      33610: inst = 32'h8220000;
      33611: inst = 32'h10408000;
      33612: inst = 32'hc404991;
      33613: inst = 32'h8220000;
      33614: inst = 32'h10408000;
      33615: inst = 32'hc404992;
      33616: inst = 32'h8220000;
      33617: inst = 32'h10408000;
      33618: inst = 32'hc404993;
      33619: inst = 32'h8220000;
      33620: inst = 32'h10408000;
      33621: inst = 32'hc404994;
      33622: inst = 32'h8220000;
      33623: inst = 32'h10408000;
      33624: inst = 32'hc404995;
      33625: inst = 32'h8220000;
      33626: inst = 32'h10408000;
      33627: inst = 32'hc404996;
      33628: inst = 32'h8220000;
      33629: inst = 32'h10408000;
      33630: inst = 32'hc404997;
      33631: inst = 32'h8220000;
      33632: inst = 32'h10408000;
      33633: inst = 32'hc404998;
      33634: inst = 32'h8220000;
      33635: inst = 32'h10408000;
      33636: inst = 32'hc404999;
      33637: inst = 32'h8220000;
      33638: inst = 32'h10408000;
      33639: inst = 32'hc40499a;
      33640: inst = 32'h8220000;
      33641: inst = 32'h10408000;
      33642: inst = 32'hc40499b;
      33643: inst = 32'h8220000;
      33644: inst = 32'h10408000;
      33645: inst = 32'hc40499c;
      33646: inst = 32'h8220000;
      33647: inst = 32'h10408000;
      33648: inst = 32'hc4049a3;
      33649: inst = 32'h8220000;
      33650: inst = 32'h10408000;
      33651: inst = 32'hc4049a4;
      33652: inst = 32'h8220000;
      33653: inst = 32'h10408000;
      33654: inst = 32'hc4049a5;
      33655: inst = 32'h8220000;
      33656: inst = 32'h10408000;
      33657: inst = 32'hc4049a6;
      33658: inst = 32'h8220000;
      33659: inst = 32'h10408000;
      33660: inst = 32'hc4049a7;
      33661: inst = 32'h8220000;
      33662: inst = 32'h10408000;
      33663: inst = 32'hc4049a8;
      33664: inst = 32'h8220000;
      33665: inst = 32'h10408000;
      33666: inst = 32'hc4049a9;
      33667: inst = 32'h8220000;
      33668: inst = 32'h10408000;
      33669: inst = 32'hc4049aa;
      33670: inst = 32'h8220000;
      33671: inst = 32'h10408000;
      33672: inst = 32'hc4049ab;
      33673: inst = 32'h8220000;
      33674: inst = 32'h10408000;
      33675: inst = 32'hc4049ac;
      33676: inst = 32'h8220000;
      33677: inst = 32'h10408000;
      33678: inst = 32'hc4049ad;
      33679: inst = 32'h8220000;
      33680: inst = 32'h10408000;
      33681: inst = 32'hc4049b1;
      33682: inst = 32'h8220000;
      33683: inst = 32'h10408000;
      33684: inst = 32'hc4049b2;
      33685: inst = 32'h8220000;
      33686: inst = 32'h10408000;
      33687: inst = 32'hc4049b3;
      33688: inst = 32'h8220000;
      33689: inst = 32'h10408000;
      33690: inst = 32'hc4049b4;
      33691: inst = 32'h8220000;
      33692: inst = 32'h10408000;
      33693: inst = 32'hc4049b5;
      33694: inst = 32'h8220000;
      33695: inst = 32'h10408000;
      33696: inst = 32'hc4049b6;
      33697: inst = 32'h8220000;
      33698: inst = 32'h10408000;
      33699: inst = 32'hc4049b7;
      33700: inst = 32'h8220000;
      33701: inst = 32'h10408000;
      33702: inst = 32'hc4049b8;
      33703: inst = 32'h8220000;
      33704: inst = 32'h10408000;
      33705: inst = 32'hc4049b9;
      33706: inst = 32'h8220000;
      33707: inst = 32'h10408000;
      33708: inst = 32'hc4049ba;
      33709: inst = 32'h8220000;
      33710: inst = 32'h10408000;
      33711: inst = 32'hc4049bb;
      33712: inst = 32'h8220000;
      33713: inst = 32'h10408000;
      33714: inst = 32'hc4049bc;
      33715: inst = 32'h8220000;
      33716: inst = 32'h10408000;
      33717: inst = 32'hc4049bd;
      33718: inst = 32'h8220000;
      33719: inst = 32'h10408000;
      33720: inst = 32'hc4049be;
      33721: inst = 32'h8220000;
      33722: inst = 32'h10408000;
      33723: inst = 32'hc4049bf;
      33724: inst = 32'h8220000;
      33725: inst = 32'h10408000;
      33726: inst = 32'hc4049c0;
      33727: inst = 32'h8220000;
      33728: inst = 32'h10408000;
      33729: inst = 32'hc4049c1;
      33730: inst = 32'h8220000;
      33731: inst = 32'h10408000;
      33732: inst = 32'hc4049c2;
      33733: inst = 32'h8220000;
      33734: inst = 32'h10408000;
      33735: inst = 32'hc4049c3;
      33736: inst = 32'h8220000;
      33737: inst = 32'h10408000;
      33738: inst = 32'hc4049c4;
      33739: inst = 32'h8220000;
      33740: inst = 32'h10408000;
      33741: inst = 32'hc4049c5;
      33742: inst = 32'h8220000;
      33743: inst = 32'h10408000;
      33744: inst = 32'hc4049c6;
      33745: inst = 32'h8220000;
      33746: inst = 32'h10408000;
      33747: inst = 32'hc4049c7;
      33748: inst = 32'h8220000;
      33749: inst = 32'h10408000;
      33750: inst = 32'hc4049c8;
      33751: inst = 32'h8220000;
      33752: inst = 32'h10408000;
      33753: inst = 32'hc4049c9;
      33754: inst = 32'h8220000;
      33755: inst = 32'h10408000;
      33756: inst = 32'hc4049ca;
      33757: inst = 32'h8220000;
      33758: inst = 32'h10408000;
      33759: inst = 32'hc4049cb;
      33760: inst = 32'h8220000;
      33761: inst = 32'h10408000;
      33762: inst = 32'hc4049cc;
      33763: inst = 32'h8220000;
      33764: inst = 32'h10408000;
      33765: inst = 32'hc4049cd;
      33766: inst = 32'h8220000;
      33767: inst = 32'h10408000;
      33768: inst = 32'hc4049ce;
      33769: inst = 32'h8220000;
      33770: inst = 32'h10408000;
      33771: inst = 32'hc4049cf;
      33772: inst = 32'h8220000;
      33773: inst = 32'h10408000;
      33774: inst = 32'hc4049d0;
      33775: inst = 32'h8220000;
      33776: inst = 32'h10408000;
      33777: inst = 32'hc4049d1;
      33778: inst = 32'h8220000;
      33779: inst = 32'h10408000;
      33780: inst = 32'hc4049d2;
      33781: inst = 32'h8220000;
      33782: inst = 32'h10408000;
      33783: inst = 32'hc4049d3;
      33784: inst = 32'h8220000;
      33785: inst = 32'h10408000;
      33786: inst = 32'hc4049d4;
      33787: inst = 32'h8220000;
      33788: inst = 32'h10408000;
      33789: inst = 32'hc4049d5;
      33790: inst = 32'h8220000;
      33791: inst = 32'h10408000;
      33792: inst = 32'hc4049d6;
      33793: inst = 32'h8220000;
      33794: inst = 32'h10408000;
      33795: inst = 32'hc4049d7;
      33796: inst = 32'h8220000;
      33797: inst = 32'h10408000;
      33798: inst = 32'hc4049d8;
      33799: inst = 32'h8220000;
      33800: inst = 32'h10408000;
      33801: inst = 32'hc4049d9;
      33802: inst = 32'h8220000;
      33803: inst = 32'h10408000;
      33804: inst = 32'hc4049da;
      33805: inst = 32'h8220000;
      33806: inst = 32'h10408000;
      33807: inst = 32'hc4049db;
      33808: inst = 32'h8220000;
      33809: inst = 32'h10408000;
      33810: inst = 32'hc4049dc;
      33811: inst = 32'h8220000;
      33812: inst = 32'h10408000;
      33813: inst = 32'hc4049dd;
      33814: inst = 32'h8220000;
      33815: inst = 32'h10408000;
      33816: inst = 32'hc4049de;
      33817: inst = 32'h8220000;
      33818: inst = 32'h10408000;
      33819: inst = 32'hc4049df;
      33820: inst = 32'h8220000;
      33821: inst = 32'h10408000;
      33822: inst = 32'hc4049e0;
      33823: inst = 32'h8220000;
      33824: inst = 32'h10408000;
      33825: inst = 32'hc4049e1;
      33826: inst = 32'h8220000;
      33827: inst = 32'h10408000;
      33828: inst = 32'hc4049e2;
      33829: inst = 32'h8220000;
      33830: inst = 32'h10408000;
      33831: inst = 32'hc4049e3;
      33832: inst = 32'h8220000;
      33833: inst = 32'h10408000;
      33834: inst = 32'hc4049e4;
      33835: inst = 32'h8220000;
      33836: inst = 32'h10408000;
      33837: inst = 32'hc4049e5;
      33838: inst = 32'h8220000;
      33839: inst = 32'h10408000;
      33840: inst = 32'hc4049ef;
      33841: inst = 32'h8220000;
      33842: inst = 32'h10408000;
      33843: inst = 32'hc4049f0;
      33844: inst = 32'h8220000;
      33845: inst = 32'h10408000;
      33846: inst = 32'hc4049f1;
      33847: inst = 32'h8220000;
      33848: inst = 32'h10408000;
      33849: inst = 32'hc4049f2;
      33850: inst = 32'h8220000;
      33851: inst = 32'h10408000;
      33852: inst = 32'hc4049f3;
      33853: inst = 32'h8220000;
      33854: inst = 32'h10408000;
      33855: inst = 32'hc4049f4;
      33856: inst = 32'h8220000;
      33857: inst = 32'h10408000;
      33858: inst = 32'hc4049f5;
      33859: inst = 32'h8220000;
      33860: inst = 32'h10408000;
      33861: inst = 32'hc4049f6;
      33862: inst = 32'h8220000;
      33863: inst = 32'h10408000;
      33864: inst = 32'hc4049f7;
      33865: inst = 32'h8220000;
      33866: inst = 32'h10408000;
      33867: inst = 32'hc4049f8;
      33868: inst = 32'h8220000;
      33869: inst = 32'h10408000;
      33870: inst = 32'hc4049f9;
      33871: inst = 32'h8220000;
      33872: inst = 32'h10408000;
      33873: inst = 32'hc4049fa;
      33874: inst = 32'h8220000;
      33875: inst = 32'h10408000;
      33876: inst = 32'hc4049fb;
      33877: inst = 32'h8220000;
      33878: inst = 32'h10408000;
      33879: inst = 32'hc4049fc;
      33880: inst = 32'h8220000;
      33881: inst = 32'h10408000;
      33882: inst = 32'hc404a03;
      33883: inst = 32'h8220000;
      33884: inst = 32'h10408000;
      33885: inst = 32'hc404a04;
      33886: inst = 32'h8220000;
      33887: inst = 32'h10408000;
      33888: inst = 32'hc404a05;
      33889: inst = 32'h8220000;
      33890: inst = 32'h10408000;
      33891: inst = 32'hc404a06;
      33892: inst = 32'h8220000;
      33893: inst = 32'h10408000;
      33894: inst = 32'hc404a07;
      33895: inst = 32'h8220000;
      33896: inst = 32'h10408000;
      33897: inst = 32'hc404a08;
      33898: inst = 32'h8220000;
      33899: inst = 32'h10408000;
      33900: inst = 32'hc404a09;
      33901: inst = 32'h8220000;
      33902: inst = 32'h10408000;
      33903: inst = 32'hc404a0a;
      33904: inst = 32'h8220000;
      33905: inst = 32'h10408000;
      33906: inst = 32'hc404a0b;
      33907: inst = 32'h8220000;
      33908: inst = 32'h10408000;
      33909: inst = 32'hc404a0c;
      33910: inst = 32'h8220000;
      33911: inst = 32'h10408000;
      33912: inst = 32'hc404a0d;
      33913: inst = 32'h8220000;
      33914: inst = 32'h10408000;
      33915: inst = 32'hc404a11;
      33916: inst = 32'h8220000;
      33917: inst = 32'h10408000;
      33918: inst = 32'hc404a12;
      33919: inst = 32'h8220000;
      33920: inst = 32'h10408000;
      33921: inst = 32'hc404a13;
      33922: inst = 32'h8220000;
      33923: inst = 32'h10408000;
      33924: inst = 32'hc404a14;
      33925: inst = 32'h8220000;
      33926: inst = 32'h10408000;
      33927: inst = 32'hc404a15;
      33928: inst = 32'h8220000;
      33929: inst = 32'h10408000;
      33930: inst = 32'hc404a16;
      33931: inst = 32'h8220000;
      33932: inst = 32'h10408000;
      33933: inst = 32'hc404a17;
      33934: inst = 32'h8220000;
      33935: inst = 32'h10408000;
      33936: inst = 32'hc404a18;
      33937: inst = 32'h8220000;
      33938: inst = 32'h10408000;
      33939: inst = 32'hc404a19;
      33940: inst = 32'h8220000;
      33941: inst = 32'h10408000;
      33942: inst = 32'hc404a1a;
      33943: inst = 32'h8220000;
      33944: inst = 32'h10408000;
      33945: inst = 32'hc404a1b;
      33946: inst = 32'h8220000;
      33947: inst = 32'h10408000;
      33948: inst = 32'hc404a1c;
      33949: inst = 32'h8220000;
      33950: inst = 32'h10408000;
      33951: inst = 32'hc404a1d;
      33952: inst = 32'h8220000;
      33953: inst = 32'h10408000;
      33954: inst = 32'hc404a1e;
      33955: inst = 32'h8220000;
      33956: inst = 32'h10408000;
      33957: inst = 32'hc404a1f;
      33958: inst = 32'h8220000;
      33959: inst = 32'h10408000;
      33960: inst = 32'hc404a20;
      33961: inst = 32'h8220000;
      33962: inst = 32'h10408000;
      33963: inst = 32'hc404a21;
      33964: inst = 32'h8220000;
      33965: inst = 32'h10408000;
      33966: inst = 32'hc404a22;
      33967: inst = 32'h8220000;
      33968: inst = 32'h10408000;
      33969: inst = 32'hc404a23;
      33970: inst = 32'h8220000;
      33971: inst = 32'h10408000;
      33972: inst = 32'hc404a24;
      33973: inst = 32'h8220000;
      33974: inst = 32'h10408000;
      33975: inst = 32'hc404a25;
      33976: inst = 32'h8220000;
      33977: inst = 32'h10408000;
      33978: inst = 32'hc404a26;
      33979: inst = 32'h8220000;
      33980: inst = 32'h10408000;
      33981: inst = 32'hc404a27;
      33982: inst = 32'h8220000;
      33983: inst = 32'h10408000;
      33984: inst = 32'hc404a28;
      33985: inst = 32'h8220000;
      33986: inst = 32'h10408000;
      33987: inst = 32'hc404a29;
      33988: inst = 32'h8220000;
      33989: inst = 32'h10408000;
      33990: inst = 32'hc404a2a;
      33991: inst = 32'h8220000;
      33992: inst = 32'h10408000;
      33993: inst = 32'hc404a2b;
      33994: inst = 32'h8220000;
      33995: inst = 32'h10408000;
      33996: inst = 32'hc404a2c;
      33997: inst = 32'h8220000;
      33998: inst = 32'h10408000;
      33999: inst = 32'hc404a2d;
      34000: inst = 32'h8220000;
      34001: inst = 32'h10408000;
      34002: inst = 32'hc404a2e;
      34003: inst = 32'h8220000;
      34004: inst = 32'h10408000;
      34005: inst = 32'hc404a2f;
      34006: inst = 32'h8220000;
      34007: inst = 32'h10408000;
      34008: inst = 32'hc404a30;
      34009: inst = 32'h8220000;
      34010: inst = 32'h10408000;
      34011: inst = 32'hc404a31;
      34012: inst = 32'h8220000;
      34013: inst = 32'h10408000;
      34014: inst = 32'hc404a32;
      34015: inst = 32'h8220000;
      34016: inst = 32'h10408000;
      34017: inst = 32'hc404a33;
      34018: inst = 32'h8220000;
      34019: inst = 32'h10408000;
      34020: inst = 32'hc404a34;
      34021: inst = 32'h8220000;
      34022: inst = 32'h10408000;
      34023: inst = 32'hc404a35;
      34024: inst = 32'h8220000;
      34025: inst = 32'h10408000;
      34026: inst = 32'hc404a36;
      34027: inst = 32'h8220000;
      34028: inst = 32'h10408000;
      34029: inst = 32'hc404a37;
      34030: inst = 32'h8220000;
      34031: inst = 32'h10408000;
      34032: inst = 32'hc404a38;
      34033: inst = 32'h8220000;
      34034: inst = 32'h10408000;
      34035: inst = 32'hc404a39;
      34036: inst = 32'h8220000;
      34037: inst = 32'h10408000;
      34038: inst = 32'hc404a3a;
      34039: inst = 32'h8220000;
      34040: inst = 32'h10408000;
      34041: inst = 32'hc404a3b;
      34042: inst = 32'h8220000;
      34043: inst = 32'h10408000;
      34044: inst = 32'hc404a3c;
      34045: inst = 32'h8220000;
      34046: inst = 32'h10408000;
      34047: inst = 32'hc404a3d;
      34048: inst = 32'h8220000;
      34049: inst = 32'h10408000;
      34050: inst = 32'hc404a3e;
      34051: inst = 32'h8220000;
      34052: inst = 32'h10408000;
      34053: inst = 32'hc404a3f;
      34054: inst = 32'h8220000;
      34055: inst = 32'h10408000;
      34056: inst = 32'hc404a40;
      34057: inst = 32'h8220000;
      34058: inst = 32'h10408000;
      34059: inst = 32'hc404a41;
      34060: inst = 32'h8220000;
      34061: inst = 32'h10408000;
      34062: inst = 32'hc404a42;
      34063: inst = 32'h8220000;
      34064: inst = 32'h10408000;
      34065: inst = 32'hc404a43;
      34066: inst = 32'h8220000;
      34067: inst = 32'h10408000;
      34068: inst = 32'hc404a44;
      34069: inst = 32'h8220000;
      34070: inst = 32'h10408000;
      34071: inst = 32'hc404a45;
      34072: inst = 32'h8220000;
      34073: inst = 32'h10408000;
      34074: inst = 32'hc404a4f;
      34075: inst = 32'h8220000;
      34076: inst = 32'h10408000;
      34077: inst = 32'hc404a50;
      34078: inst = 32'h8220000;
      34079: inst = 32'h10408000;
      34080: inst = 32'hc404a51;
      34081: inst = 32'h8220000;
      34082: inst = 32'h10408000;
      34083: inst = 32'hc404a52;
      34084: inst = 32'h8220000;
      34085: inst = 32'h10408000;
      34086: inst = 32'hc404a53;
      34087: inst = 32'h8220000;
      34088: inst = 32'h10408000;
      34089: inst = 32'hc404a54;
      34090: inst = 32'h8220000;
      34091: inst = 32'h10408000;
      34092: inst = 32'hc404a55;
      34093: inst = 32'h8220000;
      34094: inst = 32'h10408000;
      34095: inst = 32'hc404a56;
      34096: inst = 32'h8220000;
      34097: inst = 32'h10408000;
      34098: inst = 32'hc404a57;
      34099: inst = 32'h8220000;
      34100: inst = 32'h10408000;
      34101: inst = 32'hc404a58;
      34102: inst = 32'h8220000;
      34103: inst = 32'h10408000;
      34104: inst = 32'hc404a59;
      34105: inst = 32'h8220000;
      34106: inst = 32'h10408000;
      34107: inst = 32'hc404a5a;
      34108: inst = 32'h8220000;
      34109: inst = 32'h10408000;
      34110: inst = 32'hc404a5b;
      34111: inst = 32'h8220000;
      34112: inst = 32'h10408000;
      34113: inst = 32'hc404a5c;
      34114: inst = 32'h8220000;
      34115: inst = 32'h10408000;
      34116: inst = 32'hc404a63;
      34117: inst = 32'h8220000;
      34118: inst = 32'h10408000;
      34119: inst = 32'hc404a64;
      34120: inst = 32'h8220000;
      34121: inst = 32'h10408000;
      34122: inst = 32'hc404a65;
      34123: inst = 32'h8220000;
      34124: inst = 32'h10408000;
      34125: inst = 32'hc404a66;
      34126: inst = 32'h8220000;
      34127: inst = 32'h10408000;
      34128: inst = 32'hc404a67;
      34129: inst = 32'h8220000;
      34130: inst = 32'h10408000;
      34131: inst = 32'hc404a68;
      34132: inst = 32'h8220000;
      34133: inst = 32'h10408000;
      34134: inst = 32'hc404a69;
      34135: inst = 32'h8220000;
      34136: inst = 32'h10408000;
      34137: inst = 32'hc404a6a;
      34138: inst = 32'h8220000;
      34139: inst = 32'h10408000;
      34140: inst = 32'hc404a6b;
      34141: inst = 32'h8220000;
      34142: inst = 32'h10408000;
      34143: inst = 32'hc404a6c;
      34144: inst = 32'h8220000;
      34145: inst = 32'h10408000;
      34146: inst = 32'hc404a6d;
      34147: inst = 32'h8220000;
      34148: inst = 32'h10408000;
      34149: inst = 32'hc404a71;
      34150: inst = 32'h8220000;
      34151: inst = 32'h10408000;
      34152: inst = 32'hc404a72;
      34153: inst = 32'h8220000;
      34154: inst = 32'h10408000;
      34155: inst = 32'hc404a73;
      34156: inst = 32'h8220000;
      34157: inst = 32'h10408000;
      34158: inst = 32'hc404a74;
      34159: inst = 32'h8220000;
      34160: inst = 32'h10408000;
      34161: inst = 32'hc404a75;
      34162: inst = 32'h8220000;
      34163: inst = 32'h10408000;
      34164: inst = 32'hc404a76;
      34165: inst = 32'h8220000;
      34166: inst = 32'h10408000;
      34167: inst = 32'hc404a77;
      34168: inst = 32'h8220000;
      34169: inst = 32'h10408000;
      34170: inst = 32'hc404a78;
      34171: inst = 32'h8220000;
      34172: inst = 32'h10408000;
      34173: inst = 32'hc404a79;
      34174: inst = 32'h8220000;
      34175: inst = 32'h10408000;
      34176: inst = 32'hc404a7a;
      34177: inst = 32'h8220000;
      34178: inst = 32'h10408000;
      34179: inst = 32'hc404a7b;
      34180: inst = 32'h8220000;
      34181: inst = 32'h10408000;
      34182: inst = 32'hc404a7c;
      34183: inst = 32'h8220000;
      34184: inst = 32'h10408000;
      34185: inst = 32'hc404a7d;
      34186: inst = 32'h8220000;
      34187: inst = 32'h10408000;
      34188: inst = 32'hc404a7e;
      34189: inst = 32'h8220000;
      34190: inst = 32'h10408000;
      34191: inst = 32'hc404a7f;
      34192: inst = 32'h8220000;
      34193: inst = 32'h10408000;
      34194: inst = 32'hc404a80;
      34195: inst = 32'h8220000;
      34196: inst = 32'h10408000;
      34197: inst = 32'hc404a81;
      34198: inst = 32'h8220000;
      34199: inst = 32'h10408000;
      34200: inst = 32'hc404a82;
      34201: inst = 32'h8220000;
      34202: inst = 32'h10408000;
      34203: inst = 32'hc404a83;
      34204: inst = 32'h8220000;
      34205: inst = 32'h10408000;
      34206: inst = 32'hc404a84;
      34207: inst = 32'h8220000;
      34208: inst = 32'h10408000;
      34209: inst = 32'hc404a85;
      34210: inst = 32'h8220000;
      34211: inst = 32'h10408000;
      34212: inst = 32'hc404a86;
      34213: inst = 32'h8220000;
      34214: inst = 32'h10408000;
      34215: inst = 32'hc404a87;
      34216: inst = 32'h8220000;
      34217: inst = 32'h10408000;
      34218: inst = 32'hc404a88;
      34219: inst = 32'h8220000;
      34220: inst = 32'h10408000;
      34221: inst = 32'hc404a89;
      34222: inst = 32'h8220000;
      34223: inst = 32'h10408000;
      34224: inst = 32'hc404a8a;
      34225: inst = 32'h8220000;
      34226: inst = 32'h10408000;
      34227: inst = 32'hc404a8b;
      34228: inst = 32'h8220000;
      34229: inst = 32'h10408000;
      34230: inst = 32'hc404a8c;
      34231: inst = 32'h8220000;
      34232: inst = 32'h10408000;
      34233: inst = 32'hc404a8d;
      34234: inst = 32'h8220000;
      34235: inst = 32'h10408000;
      34236: inst = 32'hc404a8e;
      34237: inst = 32'h8220000;
      34238: inst = 32'h10408000;
      34239: inst = 32'hc404a8f;
      34240: inst = 32'h8220000;
      34241: inst = 32'h10408000;
      34242: inst = 32'hc404a90;
      34243: inst = 32'h8220000;
      34244: inst = 32'h10408000;
      34245: inst = 32'hc404a91;
      34246: inst = 32'h8220000;
      34247: inst = 32'h10408000;
      34248: inst = 32'hc404a92;
      34249: inst = 32'h8220000;
      34250: inst = 32'h10408000;
      34251: inst = 32'hc404a93;
      34252: inst = 32'h8220000;
      34253: inst = 32'h10408000;
      34254: inst = 32'hc404a94;
      34255: inst = 32'h8220000;
      34256: inst = 32'h10408000;
      34257: inst = 32'hc404a95;
      34258: inst = 32'h8220000;
      34259: inst = 32'h10408000;
      34260: inst = 32'hc404a96;
      34261: inst = 32'h8220000;
      34262: inst = 32'h10408000;
      34263: inst = 32'hc404a97;
      34264: inst = 32'h8220000;
      34265: inst = 32'h10408000;
      34266: inst = 32'hc404a98;
      34267: inst = 32'h8220000;
      34268: inst = 32'h10408000;
      34269: inst = 32'hc404a99;
      34270: inst = 32'h8220000;
      34271: inst = 32'h10408000;
      34272: inst = 32'hc404a9a;
      34273: inst = 32'h8220000;
      34274: inst = 32'h10408000;
      34275: inst = 32'hc404a9b;
      34276: inst = 32'h8220000;
      34277: inst = 32'h10408000;
      34278: inst = 32'hc404a9c;
      34279: inst = 32'h8220000;
      34280: inst = 32'h10408000;
      34281: inst = 32'hc404a9d;
      34282: inst = 32'h8220000;
      34283: inst = 32'h10408000;
      34284: inst = 32'hc404a9e;
      34285: inst = 32'h8220000;
      34286: inst = 32'h10408000;
      34287: inst = 32'hc404a9f;
      34288: inst = 32'h8220000;
      34289: inst = 32'h10408000;
      34290: inst = 32'hc404aa0;
      34291: inst = 32'h8220000;
      34292: inst = 32'h10408000;
      34293: inst = 32'hc404aa1;
      34294: inst = 32'h8220000;
      34295: inst = 32'h10408000;
      34296: inst = 32'hc404aa2;
      34297: inst = 32'h8220000;
      34298: inst = 32'h10408000;
      34299: inst = 32'hc404aa3;
      34300: inst = 32'h8220000;
      34301: inst = 32'h10408000;
      34302: inst = 32'hc404aa4;
      34303: inst = 32'h8220000;
      34304: inst = 32'h10408000;
      34305: inst = 32'hc404aa5;
      34306: inst = 32'h8220000;
      34307: inst = 32'h10408000;
      34308: inst = 32'hc404aa6;
      34309: inst = 32'h8220000;
      34310: inst = 32'h10408000;
      34311: inst = 32'hc404aa7;
      34312: inst = 32'h8220000;
      34313: inst = 32'h10408000;
      34314: inst = 32'hc404aa8;
      34315: inst = 32'h8220000;
      34316: inst = 32'h10408000;
      34317: inst = 32'hc404aa9;
      34318: inst = 32'h8220000;
      34319: inst = 32'h10408000;
      34320: inst = 32'hc404aaa;
      34321: inst = 32'h8220000;
      34322: inst = 32'h10408000;
      34323: inst = 32'hc404aab;
      34324: inst = 32'h8220000;
      34325: inst = 32'h10408000;
      34326: inst = 32'hc404aac;
      34327: inst = 32'h8220000;
      34328: inst = 32'h10408000;
      34329: inst = 32'hc404aad;
      34330: inst = 32'h8220000;
      34331: inst = 32'h10408000;
      34332: inst = 32'hc404aae;
      34333: inst = 32'h8220000;
      34334: inst = 32'h10408000;
      34335: inst = 32'hc404aaf;
      34336: inst = 32'h8220000;
      34337: inst = 32'h10408000;
      34338: inst = 32'hc404ab0;
      34339: inst = 32'h8220000;
      34340: inst = 32'h10408000;
      34341: inst = 32'hc404ab1;
      34342: inst = 32'h8220000;
      34343: inst = 32'h10408000;
      34344: inst = 32'hc404ab2;
      34345: inst = 32'h8220000;
      34346: inst = 32'h10408000;
      34347: inst = 32'hc404ab3;
      34348: inst = 32'h8220000;
      34349: inst = 32'h10408000;
      34350: inst = 32'hc404ab4;
      34351: inst = 32'h8220000;
      34352: inst = 32'h10408000;
      34353: inst = 32'hc404ab5;
      34354: inst = 32'h8220000;
      34355: inst = 32'h10408000;
      34356: inst = 32'hc404ab6;
      34357: inst = 32'h8220000;
      34358: inst = 32'h10408000;
      34359: inst = 32'hc404ab7;
      34360: inst = 32'h8220000;
      34361: inst = 32'h10408000;
      34362: inst = 32'hc404ab8;
      34363: inst = 32'h8220000;
      34364: inst = 32'h10408000;
      34365: inst = 32'hc404ab9;
      34366: inst = 32'h8220000;
      34367: inst = 32'h10408000;
      34368: inst = 32'hc404aba;
      34369: inst = 32'h8220000;
      34370: inst = 32'h10408000;
      34371: inst = 32'hc404abb;
      34372: inst = 32'h8220000;
      34373: inst = 32'h10408000;
      34374: inst = 32'hc404abc;
      34375: inst = 32'h8220000;
      34376: inst = 32'h10408000;
      34377: inst = 32'hc404ac3;
      34378: inst = 32'h8220000;
      34379: inst = 32'h10408000;
      34380: inst = 32'hc404ac4;
      34381: inst = 32'h8220000;
      34382: inst = 32'h10408000;
      34383: inst = 32'hc404ac5;
      34384: inst = 32'h8220000;
      34385: inst = 32'h10408000;
      34386: inst = 32'hc404ac6;
      34387: inst = 32'h8220000;
      34388: inst = 32'h10408000;
      34389: inst = 32'hc404ac7;
      34390: inst = 32'h8220000;
      34391: inst = 32'h10408000;
      34392: inst = 32'hc404ac8;
      34393: inst = 32'h8220000;
      34394: inst = 32'h10408000;
      34395: inst = 32'hc404ac9;
      34396: inst = 32'h8220000;
      34397: inst = 32'h10408000;
      34398: inst = 32'hc404aca;
      34399: inst = 32'h8220000;
      34400: inst = 32'h10408000;
      34401: inst = 32'hc404acb;
      34402: inst = 32'h8220000;
      34403: inst = 32'h10408000;
      34404: inst = 32'hc404acc;
      34405: inst = 32'h8220000;
      34406: inst = 32'h10408000;
      34407: inst = 32'hc404acd;
      34408: inst = 32'h8220000;
      34409: inst = 32'h10408000;
      34410: inst = 32'hc404ad1;
      34411: inst = 32'h8220000;
      34412: inst = 32'h10408000;
      34413: inst = 32'hc404ad2;
      34414: inst = 32'h8220000;
      34415: inst = 32'h10408000;
      34416: inst = 32'hc404ad3;
      34417: inst = 32'h8220000;
      34418: inst = 32'h10408000;
      34419: inst = 32'hc404ad4;
      34420: inst = 32'h8220000;
      34421: inst = 32'h10408000;
      34422: inst = 32'hc404ad5;
      34423: inst = 32'h8220000;
      34424: inst = 32'h10408000;
      34425: inst = 32'hc404ad6;
      34426: inst = 32'h8220000;
      34427: inst = 32'h10408000;
      34428: inst = 32'hc404ad7;
      34429: inst = 32'h8220000;
      34430: inst = 32'h10408000;
      34431: inst = 32'hc404ad8;
      34432: inst = 32'h8220000;
      34433: inst = 32'h10408000;
      34434: inst = 32'hc404ad9;
      34435: inst = 32'h8220000;
      34436: inst = 32'h10408000;
      34437: inst = 32'hc404ada;
      34438: inst = 32'h8220000;
      34439: inst = 32'h10408000;
      34440: inst = 32'hc404adb;
      34441: inst = 32'h8220000;
      34442: inst = 32'h10408000;
      34443: inst = 32'hc404adc;
      34444: inst = 32'h8220000;
      34445: inst = 32'h10408000;
      34446: inst = 32'hc404add;
      34447: inst = 32'h8220000;
      34448: inst = 32'h10408000;
      34449: inst = 32'hc404ade;
      34450: inst = 32'h8220000;
      34451: inst = 32'h10408000;
      34452: inst = 32'hc404adf;
      34453: inst = 32'h8220000;
      34454: inst = 32'h10408000;
      34455: inst = 32'hc404ae0;
      34456: inst = 32'h8220000;
      34457: inst = 32'h10408000;
      34458: inst = 32'hc404ae1;
      34459: inst = 32'h8220000;
      34460: inst = 32'h10408000;
      34461: inst = 32'hc404ae2;
      34462: inst = 32'h8220000;
      34463: inst = 32'h10408000;
      34464: inst = 32'hc404ae3;
      34465: inst = 32'h8220000;
      34466: inst = 32'h10408000;
      34467: inst = 32'hc404ae4;
      34468: inst = 32'h8220000;
      34469: inst = 32'h10408000;
      34470: inst = 32'hc404ae5;
      34471: inst = 32'h8220000;
      34472: inst = 32'h10408000;
      34473: inst = 32'hc404ae6;
      34474: inst = 32'h8220000;
      34475: inst = 32'h10408000;
      34476: inst = 32'hc404ae7;
      34477: inst = 32'h8220000;
      34478: inst = 32'h10408000;
      34479: inst = 32'hc404ae8;
      34480: inst = 32'h8220000;
      34481: inst = 32'h10408000;
      34482: inst = 32'hc404ae9;
      34483: inst = 32'h8220000;
      34484: inst = 32'h10408000;
      34485: inst = 32'hc404aea;
      34486: inst = 32'h8220000;
      34487: inst = 32'h10408000;
      34488: inst = 32'hc404aeb;
      34489: inst = 32'h8220000;
      34490: inst = 32'h10408000;
      34491: inst = 32'hc404aec;
      34492: inst = 32'h8220000;
      34493: inst = 32'h10408000;
      34494: inst = 32'hc404aed;
      34495: inst = 32'h8220000;
      34496: inst = 32'h10408000;
      34497: inst = 32'hc404aee;
      34498: inst = 32'h8220000;
      34499: inst = 32'h10408000;
      34500: inst = 32'hc404aef;
      34501: inst = 32'h8220000;
      34502: inst = 32'h10408000;
      34503: inst = 32'hc404af0;
      34504: inst = 32'h8220000;
      34505: inst = 32'h10408000;
      34506: inst = 32'hc404af1;
      34507: inst = 32'h8220000;
      34508: inst = 32'h10408000;
      34509: inst = 32'hc404af2;
      34510: inst = 32'h8220000;
      34511: inst = 32'h10408000;
      34512: inst = 32'hc404af3;
      34513: inst = 32'h8220000;
      34514: inst = 32'h10408000;
      34515: inst = 32'hc404af4;
      34516: inst = 32'h8220000;
      34517: inst = 32'h10408000;
      34518: inst = 32'hc404af5;
      34519: inst = 32'h8220000;
      34520: inst = 32'h10408000;
      34521: inst = 32'hc404af6;
      34522: inst = 32'h8220000;
      34523: inst = 32'h10408000;
      34524: inst = 32'hc404af7;
      34525: inst = 32'h8220000;
      34526: inst = 32'h10408000;
      34527: inst = 32'hc404af8;
      34528: inst = 32'h8220000;
      34529: inst = 32'h10408000;
      34530: inst = 32'hc404af9;
      34531: inst = 32'h8220000;
      34532: inst = 32'h10408000;
      34533: inst = 32'hc404afa;
      34534: inst = 32'h8220000;
      34535: inst = 32'h10408000;
      34536: inst = 32'hc404afb;
      34537: inst = 32'h8220000;
      34538: inst = 32'h10408000;
      34539: inst = 32'hc404afc;
      34540: inst = 32'h8220000;
      34541: inst = 32'h10408000;
      34542: inst = 32'hc404afd;
      34543: inst = 32'h8220000;
      34544: inst = 32'h10408000;
      34545: inst = 32'hc404afe;
      34546: inst = 32'h8220000;
      34547: inst = 32'h10408000;
      34548: inst = 32'hc404aff;
      34549: inst = 32'h8220000;
      34550: inst = 32'h10408000;
      34551: inst = 32'hc404b00;
      34552: inst = 32'h8220000;
      34553: inst = 32'h10408000;
      34554: inst = 32'hc404b01;
      34555: inst = 32'h8220000;
      34556: inst = 32'h10408000;
      34557: inst = 32'hc404b02;
      34558: inst = 32'h8220000;
      34559: inst = 32'h10408000;
      34560: inst = 32'hc404b03;
      34561: inst = 32'h8220000;
      34562: inst = 32'h10408000;
      34563: inst = 32'hc404b04;
      34564: inst = 32'h8220000;
      34565: inst = 32'h10408000;
      34566: inst = 32'hc404b05;
      34567: inst = 32'h8220000;
      34568: inst = 32'h10408000;
      34569: inst = 32'hc404b06;
      34570: inst = 32'h8220000;
      34571: inst = 32'h10408000;
      34572: inst = 32'hc404b07;
      34573: inst = 32'h8220000;
      34574: inst = 32'h10408000;
      34575: inst = 32'hc404b08;
      34576: inst = 32'h8220000;
      34577: inst = 32'h10408000;
      34578: inst = 32'hc404b09;
      34579: inst = 32'h8220000;
      34580: inst = 32'h10408000;
      34581: inst = 32'hc404b0a;
      34582: inst = 32'h8220000;
      34583: inst = 32'h10408000;
      34584: inst = 32'hc404b0b;
      34585: inst = 32'h8220000;
      34586: inst = 32'h10408000;
      34587: inst = 32'hc404b0c;
      34588: inst = 32'h8220000;
      34589: inst = 32'h10408000;
      34590: inst = 32'hc404b0d;
      34591: inst = 32'h8220000;
      34592: inst = 32'h10408000;
      34593: inst = 32'hc404b0e;
      34594: inst = 32'h8220000;
      34595: inst = 32'h10408000;
      34596: inst = 32'hc404b0f;
      34597: inst = 32'h8220000;
      34598: inst = 32'h10408000;
      34599: inst = 32'hc404b10;
      34600: inst = 32'h8220000;
      34601: inst = 32'h10408000;
      34602: inst = 32'hc404b11;
      34603: inst = 32'h8220000;
      34604: inst = 32'h10408000;
      34605: inst = 32'hc404b12;
      34606: inst = 32'h8220000;
      34607: inst = 32'h10408000;
      34608: inst = 32'hc404b13;
      34609: inst = 32'h8220000;
      34610: inst = 32'h10408000;
      34611: inst = 32'hc404b14;
      34612: inst = 32'h8220000;
      34613: inst = 32'h10408000;
      34614: inst = 32'hc404b15;
      34615: inst = 32'h8220000;
      34616: inst = 32'h10408000;
      34617: inst = 32'hc404b16;
      34618: inst = 32'h8220000;
      34619: inst = 32'h10408000;
      34620: inst = 32'hc404b17;
      34621: inst = 32'h8220000;
      34622: inst = 32'h10408000;
      34623: inst = 32'hc404b18;
      34624: inst = 32'h8220000;
      34625: inst = 32'h10408000;
      34626: inst = 32'hc404b19;
      34627: inst = 32'h8220000;
      34628: inst = 32'h10408000;
      34629: inst = 32'hc404b1a;
      34630: inst = 32'h8220000;
      34631: inst = 32'h10408000;
      34632: inst = 32'hc404b1b;
      34633: inst = 32'h8220000;
      34634: inst = 32'h10408000;
      34635: inst = 32'hc404b1c;
      34636: inst = 32'h8220000;
      34637: inst = 32'h10408000;
      34638: inst = 32'hc404b31;
      34639: inst = 32'h8220000;
      34640: inst = 32'h10408000;
      34641: inst = 32'hc404b32;
      34642: inst = 32'h8220000;
      34643: inst = 32'h10408000;
      34644: inst = 32'hc404b33;
      34645: inst = 32'h8220000;
      34646: inst = 32'h10408000;
      34647: inst = 32'hc404b34;
      34648: inst = 32'h8220000;
      34649: inst = 32'h10408000;
      34650: inst = 32'hc404b35;
      34651: inst = 32'h8220000;
      34652: inst = 32'h10408000;
      34653: inst = 32'hc404b36;
      34654: inst = 32'h8220000;
      34655: inst = 32'h10408000;
      34656: inst = 32'hc404b37;
      34657: inst = 32'h8220000;
      34658: inst = 32'h10408000;
      34659: inst = 32'hc404b38;
      34660: inst = 32'h8220000;
      34661: inst = 32'h10408000;
      34662: inst = 32'hc404b39;
      34663: inst = 32'h8220000;
      34664: inst = 32'h10408000;
      34665: inst = 32'hc404b3a;
      34666: inst = 32'h8220000;
      34667: inst = 32'h10408000;
      34668: inst = 32'hc404b3b;
      34669: inst = 32'h8220000;
      34670: inst = 32'h10408000;
      34671: inst = 32'hc404b3c;
      34672: inst = 32'h8220000;
      34673: inst = 32'h10408000;
      34674: inst = 32'hc404b3d;
      34675: inst = 32'h8220000;
      34676: inst = 32'h10408000;
      34677: inst = 32'hc404b3e;
      34678: inst = 32'h8220000;
      34679: inst = 32'h10408000;
      34680: inst = 32'hc404b3f;
      34681: inst = 32'h8220000;
      34682: inst = 32'h10408000;
      34683: inst = 32'hc404b40;
      34684: inst = 32'h8220000;
      34685: inst = 32'h10408000;
      34686: inst = 32'hc404b41;
      34687: inst = 32'h8220000;
      34688: inst = 32'h10408000;
      34689: inst = 32'hc404b42;
      34690: inst = 32'h8220000;
      34691: inst = 32'h10408000;
      34692: inst = 32'hc404b43;
      34693: inst = 32'h8220000;
      34694: inst = 32'h10408000;
      34695: inst = 32'hc404b44;
      34696: inst = 32'h8220000;
      34697: inst = 32'h10408000;
      34698: inst = 32'hc404b45;
      34699: inst = 32'h8220000;
      34700: inst = 32'h10408000;
      34701: inst = 32'hc404b46;
      34702: inst = 32'h8220000;
      34703: inst = 32'h10408000;
      34704: inst = 32'hc404b47;
      34705: inst = 32'h8220000;
      34706: inst = 32'h10408000;
      34707: inst = 32'hc404b48;
      34708: inst = 32'h8220000;
      34709: inst = 32'h10408000;
      34710: inst = 32'hc404b49;
      34711: inst = 32'h8220000;
      34712: inst = 32'h10408000;
      34713: inst = 32'hc404b4a;
      34714: inst = 32'h8220000;
      34715: inst = 32'h10408000;
      34716: inst = 32'hc404b4b;
      34717: inst = 32'h8220000;
      34718: inst = 32'h10408000;
      34719: inst = 32'hc404b4c;
      34720: inst = 32'h8220000;
      34721: inst = 32'h10408000;
      34722: inst = 32'hc404b4d;
      34723: inst = 32'h8220000;
      34724: inst = 32'h10408000;
      34725: inst = 32'hc404b4e;
      34726: inst = 32'h8220000;
      34727: inst = 32'h10408000;
      34728: inst = 32'hc404b4f;
      34729: inst = 32'h8220000;
      34730: inst = 32'h10408000;
      34731: inst = 32'hc404b50;
      34732: inst = 32'h8220000;
      34733: inst = 32'h10408000;
      34734: inst = 32'hc404b51;
      34735: inst = 32'h8220000;
      34736: inst = 32'h10408000;
      34737: inst = 32'hc404b52;
      34738: inst = 32'h8220000;
      34739: inst = 32'h10408000;
      34740: inst = 32'hc404b53;
      34741: inst = 32'h8220000;
      34742: inst = 32'h10408000;
      34743: inst = 32'hc404b54;
      34744: inst = 32'h8220000;
      34745: inst = 32'h10408000;
      34746: inst = 32'hc404b55;
      34747: inst = 32'h8220000;
      34748: inst = 32'h10408000;
      34749: inst = 32'hc404b56;
      34750: inst = 32'h8220000;
      34751: inst = 32'h10408000;
      34752: inst = 32'hc404b57;
      34753: inst = 32'h8220000;
      34754: inst = 32'h10408000;
      34755: inst = 32'hc404b58;
      34756: inst = 32'h8220000;
      34757: inst = 32'h10408000;
      34758: inst = 32'hc404b59;
      34759: inst = 32'h8220000;
      34760: inst = 32'h10408000;
      34761: inst = 32'hc404b5a;
      34762: inst = 32'h8220000;
      34763: inst = 32'h10408000;
      34764: inst = 32'hc404b5b;
      34765: inst = 32'h8220000;
      34766: inst = 32'h10408000;
      34767: inst = 32'hc404b5c;
      34768: inst = 32'h8220000;
      34769: inst = 32'h10408000;
      34770: inst = 32'hc404b5d;
      34771: inst = 32'h8220000;
      34772: inst = 32'h10408000;
      34773: inst = 32'hc404b5e;
      34774: inst = 32'h8220000;
      34775: inst = 32'h10408000;
      34776: inst = 32'hc404b5f;
      34777: inst = 32'h8220000;
      34778: inst = 32'h10408000;
      34779: inst = 32'hc404b60;
      34780: inst = 32'h8220000;
      34781: inst = 32'h10408000;
      34782: inst = 32'hc404b61;
      34783: inst = 32'h8220000;
      34784: inst = 32'h10408000;
      34785: inst = 32'hc404b62;
      34786: inst = 32'h8220000;
      34787: inst = 32'h10408000;
      34788: inst = 32'hc404b63;
      34789: inst = 32'h8220000;
      34790: inst = 32'h10408000;
      34791: inst = 32'hc404b64;
      34792: inst = 32'h8220000;
      34793: inst = 32'h10408000;
      34794: inst = 32'hc404b65;
      34795: inst = 32'h8220000;
      34796: inst = 32'h10408000;
      34797: inst = 32'hc404b66;
      34798: inst = 32'h8220000;
      34799: inst = 32'h10408000;
      34800: inst = 32'hc404b67;
      34801: inst = 32'h8220000;
      34802: inst = 32'h10408000;
      34803: inst = 32'hc404b68;
      34804: inst = 32'h8220000;
      34805: inst = 32'h10408000;
      34806: inst = 32'hc404b69;
      34807: inst = 32'h8220000;
      34808: inst = 32'h10408000;
      34809: inst = 32'hc404b6a;
      34810: inst = 32'h8220000;
      34811: inst = 32'h10408000;
      34812: inst = 32'hc404b6b;
      34813: inst = 32'h8220000;
      34814: inst = 32'h10408000;
      34815: inst = 32'hc404b6c;
      34816: inst = 32'h8220000;
      34817: inst = 32'h10408000;
      34818: inst = 32'hc404b6d;
      34819: inst = 32'h8220000;
      34820: inst = 32'h10408000;
      34821: inst = 32'hc404b6e;
      34822: inst = 32'h8220000;
      34823: inst = 32'h10408000;
      34824: inst = 32'hc404b6f;
      34825: inst = 32'h8220000;
      34826: inst = 32'h10408000;
      34827: inst = 32'hc404b70;
      34828: inst = 32'h8220000;
      34829: inst = 32'h10408000;
      34830: inst = 32'hc404b71;
      34831: inst = 32'h8220000;
      34832: inst = 32'h10408000;
      34833: inst = 32'hc404b72;
      34834: inst = 32'h8220000;
      34835: inst = 32'h10408000;
      34836: inst = 32'hc404b73;
      34837: inst = 32'h8220000;
      34838: inst = 32'h10408000;
      34839: inst = 32'hc404b74;
      34840: inst = 32'h8220000;
      34841: inst = 32'h10408000;
      34842: inst = 32'hc404b75;
      34843: inst = 32'h8220000;
      34844: inst = 32'h10408000;
      34845: inst = 32'hc404b76;
      34846: inst = 32'h8220000;
      34847: inst = 32'h10408000;
      34848: inst = 32'hc404b77;
      34849: inst = 32'h8220000;
      34850: inst = 32'h10408000;
      34851: inst = 32'hc404b78;
      34852: inst = 32'h8220000;
      34853: inst = 32'h10408000;
      34854: inst = 32'hc404b79;
      34855: inst = 32'h8220000;
      34856: inst = 32'h10408000;
      34857: inst = 32'hc404b7a;
      34858: inst = 32'h8220000;
      34859: inst = 32'h10408000;
      34860: inst = 32'hc404b7b;
      34861: inst = 32'h8220000;
      34862: inst = 32'h10408000;
      34863: inst = 32'hc404b7c;
      34864: inst = 32'h8220000;
      34865: inst = 32'h10408000;
      34866: inst = 32'hc404b91;
      34867: inst = 32'h8220000;
      34868: inst = 32'h10408000;
      34869: inst = 32'hc404b92;
      34870: inst = 32'h8220000;
      34871: inst = 32'h10408000;
      34872: inst = 32'hc404b93;
      34873: inst = 32'h8220000;
      34874: inst = 32'h10408000;
      34875: inst = 32'hc404b94;
      34876: inst = 32'h8220000;
      34877: inst = 32'h10408000;
      34878: inst = 32'hc404b95;
      34879: inst = 32'h8220000;
      34880: inst = 32'h10408000;
      34881: inst = 32'hc404b96;
      34882: inst = 32'h8220000;
      34883: inst = 32'h10408000;
      34884: inst = 32'hc404b97;
      34885: inst = 32'h8220000;
      34886: inst = 32'h10408000;
      34887: inst = 32'hc404b98;
      34888: inst = 32'h8220000;
      34889: inst = 32'h10408000;
      34890: inst = 32'hc404b99;
      34891: inst = 32'h8220000;
      34892: inst = 32'h10408000;
      34893: inst = 32'hc404b9a;
      34894: inst = 32'h8220000;
      34895: inst = 32'h10408000;
      34896: inst = 32'hc404b9b;
      34897: inst = 32'h8220000;
      34898: inst = 32'h10408000;
      34899: inst = 32'hc404b9c;
      34900: inst = 32'h8220000;
      34901: inst = 32'h10408000;
      34902: inst = 32'hc404b9d;
      34903: inst = 32'h8220000;
      34904: inst = 32'h10408000;
      34905: inst = 32'hc404b9e;
      34906: inst = 32'h8220000;
      34907: inst = 32'h10408000;
      34908: inst = 32'hc404b9f;
      34909: inst = 32'h8220000;
      34910: inst = 32'h10408000;
      34911: inst = 32'hc404ba0;
      34912: inst = 32'h8220000;
      34913: inst = 32'h10408000;
      34914: inst = 32'hc404ba1;
      34915: inst = 32'h8220000;
      34916: inst = 32'h10408000;
      34917: inst = 32'hc404ba2;
      34918: inst = 32'h8220000;
      34919: inst = 32'h10408000;
      34920: inst = 32'hc404ba3;
      34921: inst = 32'h8220000;
      34922: inst = 32'h10408000;
      34923: inst = 32'hc404ba4;
      34924: inst = 32'h8220000;
      34925: inst = 32'h10408000;
      34926: inst = 32'hc404ba5;
      34927: inst = 32'h8220000;
      34928: inst = 32'h10408000;
      34929: inst = 32'hc404ba6;
      34930: inst = 32'h8220000;
      34931: inst = 32'h10408000;
      34932: inst = 32'hc404ba7;
      34933: inst = 32'h8220000;
      34934: inst = 32'h10408000;
      34935: inst = 32'hc404ba8;
      34936: inst = 32'h8220000;
      34937: inst = 32'h10408000;
      34938: inst = 32'hc404ba9;
      34939: inst = 32'h8220000;
      34940: inst = 32'h10408000;
      34941: inst = 32'hc404baa;
      34942: inst = 32'h8220000;
      34943: inst = 32'h10408000;
      34944: inst = 32'hc404bab;
      34945: inst = 32'h8220000;
      34946: inst = 32'h10408000;
      34947: inst = 32'hc404bac;
      34948: inst = 32'h8220000;
      34949: inst = 32'h10408000;
      34950: inst = 32'hc404bad;
      34951: inst = 32'h8220000;
      34952: inst = 32'h10408000;
      34953: inst = 32'hc404bae;
      34954: inst = 32'h8220000;
      34955: inst = 32'h10408000;
      34956: inst = 32'hc404baf;
      34957: inst = 32'h8220000;
      34958: inst = 32'h10408000;
      34959: inst = 32'hc404bb0;
      34960: inst = 32'h8220000;
      34961: inst = 32'h10408000;
      34962: inst = 32'hc404bb1;
      34963: inst = 32'h8220000;
      34964: inst = 32'h10408000;
      34965: inst = 32'hc404bb2;
      34966: inst = 32'h8220000;
      34967: inst = 32'h10408000;
      34968: inst = 32'hc404bb3;
      34969: inst = 32'h8220000;
      34970: inst = 32'h10408000;
      34971: inst = 32'hc404bb4;
      34972: inst = 32'h8220000;
      34973: inst = 32'h10408000;
      34974: inst = 32'hc404bb5;
      34975: inst = 32'h8220000;
      34976: inst = 32'h10408000;
      34977: inst = 32'hc404bb6;
      34978: inst = 32'h8220000;
      34979: inst = 32'h10408000;
      34980: inst = 32'hc404bb7;
      34981: inst = 32'h8220000;
      34982: inst = 32'h10408000;
      34983: inst = 32'hc404bb8;
      34984: inst = 32'h8220000;
      34985: inst = 32'h10408000;
      34986: inst = 32'hc404bb9;
      34987: inst = 32'h8220000;
      34988: inst = 32'h10408000;
      34989: inst = 32'hc404bba;
      34990: inst = 32'h8220000;
      34991: inst = 32'h10408000;
      34992: inst = 32'hc404bbb;
      34993: inst = 32'h8220000;
      34994: inst = 32'h10408000;
      34995: inst = 32'hc404bbc;
      34996: inst = 32'h8220000;
      34997: inst = 32'h10408000;
      34998: inst = 32'hc404bbd;
      34999: inst = 32'h8220000;
      35000: inst = 32'h10408000;
      35001: inst = 32'hc404bbe;
      35002: inst = 32'h8220000;
      35003: inst = 32'h10408000;
      35004: inst = 32'hc404bbf;
      35005: inst = 32'h8220000;
      35006: inst = 32'h10408000;
      35007: inst = 32'hc404bc0;
      35008: inst = 32'h8220000;
      35009: inst = 32'h10408000;
      35010: inst = 32'hc404bc1;
      35011: inst = 32'h8220000;
      35012: inst = 32'h10408000;
      35013: inst = 32'hc404bc2;
      35014: inst = 32'h8220000;
      35015: inst = 32'h10408000;
      35016: inst = 32'hc404bc3;
      35017: inst = 32'h8220000;
      35018: inst = 32'h10408000;
      35019: inst = 32'hc404bc4;
      35020: inst = 32'h8220000;
      35021: inst = 32'h10408000;
      35022: inst = 32'hc404bc5;
      35023: inst = 32'h8220000;
      35024: inst = 32'h10408000;
      35025: inst = 32'hc404bc6;
      35026: inst = 32'h8220000;
      35027: inst = 32'h10408000;
      35028: inst = 32'hc404bc7;
      35029: inst = 32'h8220000;
      35030: inst = 32'h10408000;
      35031: inst = 32'hc404bc8;
      35032: inst = 32'h8220000;
      35033: inst = 32'h10408000;
      35034: inst = 32'hc404bc9;
      35035: inst = 32'h8220000;
      35036: inst = 32'h10408000;
      35037: inst = 32'hc404bca;
      35038: inst = 32'h8220000;
      35039: inst = 32'h10408000;
      35040: inst = 32'hc404bcb;
      35041: inst = 32'h8220000;
      35042: inst = 32'h10408000;
      35043: inst = 32'hc404bcc;
      35044: inst = 32'h8220000;
      35045: inst = 32'h10408000;
      35046: inst = 32'hc404bcd;
      35047: inst = 32'h8220000;
      35048: inst = 32'h10408000;
      35049: inst = 32'hc404bce;
      35050: inst = 32'h8220000;
      35051: inst = 32'h10408000;
      35052: inst = 32'hc404bcf;
      35053: inst = 32'h8220000;
      35054: inst = 32'h10408000;
      35055: inst = 32'hc404bd0;
      35056: inst = 32'h8220000;
      35057: inst = 32'h10408000;
      35058: inst = 32'hc404bd1;
      35059: inst = 32'h8220000;
      35060: inst = 32'h10408000;
      35061: inst = 32'hc404bd2;
      35062: inst = 32'h8220000;
      35063: inst = 32'h10408000;
      35064: inst = 32'hc404bd3;
      35065: inst = 32'h8220000;
      35066: inst = 32'h10408000;
      35067: inst = 32'hc404bd4;
      35068: inst = 32'h8220000;
      35069: inst = 32'h10408000;
      35070: inst = 32'hc404bd5;
      35071: inst = 32'h8220000;
      35072: inst = 32'h10408000;
      35073: inst = 32'hc404bd6;
      35074: inst = 32'h8220000;
      35075: inst = 32'h10408000;
      35076: inst = 32'hc404bd7;
      35077: inst = 32'h8220000;
      35078: inst = 32'h10408000;
      35079: inst = 32'hc404bd8;
      35080: inst = 32'h8220000;
      35081: inst = 32'h10408000;
      35082: inst = 32'hc404bd9;
      35083: inst = 32'h8220000;
      35084: inst = 32'h10408000;
      35085: inst = 32'hc404bda;
      35086: inst = 32'h8220000;
      35087: inst = 32'h10408000;
      35088: inst = 32'hc404bdb;
      35089: inst = 32'h8220000;
      35090: inst = 32'h10408000;
      35091: inst = 32'hc404bdc;
      35092: inst = 32'h8220000;
      35093: inst = 32'h10408000;
      35094: inst = 32'hc404bf1;
      35095: inst = 32'h8220000;
      35096: inst = 32'h10408000;
      35097: inst = 32'hc404bf2;
      35098: inst = 32'h8220000;
      35099: inst = 32'h10408000;
      35100: inst = 32'hc404bf3;
      35101: inst = 32'h8220000;
      35102: inst = 32'h10408000;
      35103: inst = 32'hc404bf4;
      35104: inst = 32'h8220000;
      35105: inst = 32'h10408000;
      35106: inst = 32'hc404bf5;
      35107: inst = 32'h8220000;
      35108: inst = 32'h10408000;
      35109: inst = 32'hc404bf6;
      35110: inst = 32'h8220000;
      35111: inst = 32'h10408000;
      35112: inst = 32'hc404bf7;
      35113: inst = 32'h8220000;
      35114: inst = 32'h10408000;
      35115: inst = 32'hc404bf8;
      35116: inst = 32'h8220000;
      35117: inst = 32'h10408000;
      35118: inst = 32'hc404bf9;
      35119: inst = 32'h8220000;
      35120: inst = 32'h10408000;
      35121: inst = 32'hc404bfa;
      35122: inst = 32'h8220000;
      35123: inst = 32'h10408000;
      35124: inst = 32'hc404bfb;
      35125: inst = 32'h8220000;
      35126: inst = 32'h10408000;
      35127: inst = 32'hc404bfc;
      35128: inst = 32'h8220000;
      35129: inst = 32'h10408000;
      35130: inst = 32'hc404bfd;
      35131: inst = 32'h8220000;
      35132: inst = 32'h10408000;
      35133: inst = 32'hc404bfe;
      35134: inst = 32'h8220000;
      35135: inst = 32'h10408000;
      35136: inst = 32'hc404bff;
      35137: inst = 32'h8220000;
      35138: inst = 32'h10408000;
      35139: inst = 32'hc404c00;
      35140: inst = 32'h8220000;
      35141: inst = 32'h10408000;
      35142: inst = 32'hc404c01;
      35143: inst = 32'h8220000;
      35144: inst = 32'h10408000;
      35145: inst = 32'hc404c02;
      35146: inst = 32'h8220000;
      35147: inst = 32'h10408000;
      35148: inst = 32'hc404c03;
      35149: inst = 32'h8220000;
      35150: inst = 32'h10408000;
      35151: inst = 32'hc404c04;
      35152: inst = 32'h8220000;
      35153: inst = 32'h10408000;
      35154: inst = 32'hc404c05;
      35155: inst = 32'h8220000;
      35156: inst = 32'h10408000;
      35157: inst = 32'hc404c06;
      35158: inst = 32'h8220000;
      35159: inst = 32'h10408000;
      35160: inst = 32'hc404c07;
      35161: inst = 32'h8220000;
      35162: inst = 32'h10408000;
      35163: inst = 32'hc404c08;
      35164: inst = 32'h8220000;
      35165: inst = 32'h10408000;
      35166: inst = 32'hc404c09;
      35167: inst = 32'h8220000;
      35168: inst = 32'h10408000;
      35169: inst = 32'hc404c0a;
      35170: inst = 32'h8220000;
      35171: inst = 32'h10408000;
      35172: inst = 32'hc404c0b;
      35173: inst = 32'h8220000;
      35174: inst = 32'h10408000;
      35175: inst = 32'hc404c0c;
      35176: inst = 32'h8220000;
      35177: inst = 32'h10408000;
      35178: inst = 32'hc404c0d;
      35179: inst = 32'h8220000;
      35180: inst = 32'h10408000;
      35181: inst = 32'hc404c0e;
      35182: inst = 32'h8220000;
      35183: inst = 32'h10408000;
      35184: inst = 32'hc404c0f;
      35185: inst = 32'h8220000;
      35186: inst = 32'h10408000;
      35187: inst = 32'hc404c10;
      35188: inst = 32'h8220000;
      35189: inst = 32'h10408000;
      35190: inst = 32'hc404c11;
      35191: inst = 32'h8220000;
      35192: inst = 32'h10408000;
      35193: inst = 32'hc404c12;
      35194: inst = 32'h8220000;
      35195: inst = 32'h10408000;
      35196: inst = 32'hc404c13;
      35197: inst = 32'h8220000;
      35198: inst = 32'h10408000;
      35199: inst = 32'hc404c14;
      35200: inst = 32'h8220000;
      35201: inst = 32'h10408000;
      35202: inst = 32'hc404c15;
      35203: inst = 32'h8220000;
      35204: inst = 32'h10408000;
      35205: inst = 32'hc404c16;
      35206: inst = 32'h8220000;
      35207: inst = 32'h10408000;
      35208: inst = 32'hc404c17;
      35209: inst = 32'h8220000;
      35210: inst = 32'h10408000;
      35211: inst = 32'hc404c18;
      35212: inst = 32'h8220000;
      35213: inst = 32'h10408000;
      35214: inst = 32'hc404c19;
      35215: inst = 32'h8220000;
      35216: inst = 32'h10408000;
      35217: inst = 32'hc404c1a;
      35218: inst = 32'h8220000;
      35219: inst = 32'h10408000;
      35220: inst = 32'hc404c1b;
      35221: inst = 32'h8220000;
      35222: inst = 32'h10408000;
      35223: inst = 32'hc404c1c;
      35224: inst = 32'h8220000;
      35225: inst = 32'h10408000;
      35226: inst = 32'hc404c1d;
      35227: inst = 32'h8220000;
      35228: inst = 32'h10408000;
      35229: inst = 32'hc404c1e;
      35230: inst = 32'h8220000;
      35231: inst = 32'h10408000;
      35232: inst = 32'hc404c1f;
      35233: inst = 32'h8220000;
      35234: inst = 32'h10408000;
      35235: inst = 32'hc404c20;
      35236: inst = 32'h8220000;
      35237: inst = 32'h10408000;
      35238: inst = 32'hc404c21;
      35239: inst = 32'h8220000;
      35240: inst = 32'h10408000;
      35241: inst = 32'hc404c22;
      35242: inst = 32'h8220000;
      35243: inst = 32'h10408000;
      35244: inst = 32'hc404c23;
      35245: inst = 32'h8220000;
      35246: inst = 32'h10408000;
      35247: inst = 32'hc404c24;
      35248: inst = 32'h8220000;
      35249: inst = 32'h10408000;
      35250: inst = 32'hc404c25;
      35251: inst = 32'h8220000;
      35252: inst = 32'h10408000;
      35253: inst = 32'hc404c26;
      35254: inst = 32'h8220000;
      35255: inst = 32'h10408000;
      35256: inst = 32'hc404c27;
      35257: inst = 32'h8220000;
      35258: inst = 32'h10408000;
      35259: inst = 32'hc404c28;
      35260: inst = 32'h8220000;
      35261: inst = 32'h10408000;
      35262: inst = 32'hc404c29;
      35263: inst = 32'h8220000;
      35264: inst = 32'h10408000;
      35265: inst = 32'hc404c2a;
      35266: inst = 32'h8220000;
      35267: inst = 32'h10408000;
      35268: inst = 32'hc404c2b;
      35269: inst = 32'h8220000;
      35270: inst = 32'h10408000;
      35271: inst = 32'hc404c2c;
      35272: inst = 32'h8220000;
      35273: inst = 32'h10408000;
      35274: inst = 32'hc404c2d;
      35275: inst = 32'h8220000;
      35276: inst = 32'h10408000;
      35277: inst = 32'hc404c2e;
      35278: inst = 32'h8220000;
      35279: inst = 32'h10408000;
      35280: inst = 32'hc404c2f;
      35281: inst = 32'h8220000;
      35282: inst = 32'h10408000;
      35283: inst = 32'hc404c30;
      35284: inst = 32'h8220000;
      35285: inst = 32'h10408000;
      35286: inst = 32'hc404c31;
      35287: inst = 32'h8220000;
      35288: inst = 32'h10408000;
      35289: inst = 32'hc404c32;
      35290: inst = 32'h8220000;
      35291: inst = 32'h10408000;
      35292: inst = 32'hc404c33;
      35293: inst = 32'h8220000;
      35294: inst = 32'h10408000;
      35295: inst = 32'hc404c34;
      35296: inst = 32'h8220000;
      35297: inst = 32'h10408000;
      35298: inst = 32'hc404c35;
      35299: inst = 32'h8220000;
      35300: inst = 32'h10408000;
      35301: inst = 32'hc404c36;
      35302: inst = 32'h8220000;
      35303: inst = 32'h10408000;
      35304: inst = 32'hc404c37;
      35305: inst = 32'h8220000;
      35306: inst = 32'h10408000;
      35307: inst = 32'hc404c38;
      35308: inst = 32'h8220000;
      35309: inst = 32'h10408000;
      35310: inst = 32'hc404c39;
      35311: inst = 32'h8220000;
      35312: inst = 32'h10408000;
      35313: inst = 32'hc404c3a;
      35314: inst = 32'h8220000;
      35315: inst = 32'h10408000;
      35316: inst = 32'hc404c3b;
      35317: inst = 32'h8220000;
      35318: inst = 32'h10408000;
      35319: inst = 32'hc404c3c;
      35320: inst = 32'h8220000;
      35321: inst = 32'h10408000;
      35322: inst = 32'hc404c43;
      35323: inst = 32'h8220000;
      35324: inst = 32'h10408000;
      35325: inst = 32'hc404c44;
      35326: inst = 32'h8220000;
      35327: inst = 32'h10408000;
      35328: inst = 32'hc404c45;
      35329: inst = 32'h8220000;
      35330: inst = 32'h10408000;
      35331: inst = 32'hc404c46;
      35332: inst = 32'h8220000;
      35333: inst = 32'h10408000;
      35334: inst = 32'hc404c47;
      35335: inst = 32'h8220000;
      35336: inst = 32'h10408000;
      35337: inst = 32'hc404c48;
      35338: inst = 32'h8220000;
      35339: inst = 32'h10408000;
      35340: inst = 32'hc404c49;
      35341: inst = 32'h8220000;
      35342: inst = 32'h10408000;
      35343: inst = 32'hc404c4a;
      35344: inst = 32'h8220000;
      35345: inst = 32'h10408000;
      35346: inst = 32'hc404c4b;
      35347: inst = 32'h8220000;
      35348: inst = 32'h10408000;
      35349: inst = 32'hc404c4c;
      35350: inst = 32'h8220000;
      35351: inst = 32'h10408000;
      35352: inst = 32'hc404c4d;
      35353: inst = 32'h8220000;
      35354: inst = 32'h10408000;
      35355: inst = 32'hc404c4e;
      35356: inst = 32'h8220000;
      35357: inst = 32'h10408000;
      35358: inst = 32'hc404c4f;
      35359: inst = 32'h8220000;
      35360: inst = 32'h10408000;
      35361: inst = 32'hc404c50;
      35362: inst = 32'h8220000;
      35363: inst = 32'h10408000;
      35364: inst = 32'hc404c51;
      35365: inst = 32'h8220000;
      35366: inst = 32'h10408000;
      35367: inst = 32'hc404c52;
      35368: inst = 32'h8220000;
      35369: inst = 32'h10408000;
      35370: inst = 32'hc404c53;
      35371: inst = 32'h8220000;
      35372: inst = 32'h10408000;
      35373: inst = 32'hc404c54;
      35374: inst = 32'h8220000;
      35375: inst = 32'h10408000;
      35376: inst = 32'hc404c55;
      35377: inst = 32'h8220000;
      35378: inst = 32'h10408000;
      35379: inst = 32'hc404c56;
      35380: inst = 32'h8220000;
      35381: inst = 32'h10408000;
      35382: inst = 32'hc404c57;
      35383: inst = 32'h8220000;
      35384: inst = 32'h10408000;
      35385: inst = 32'hc404c58;
      35386: inst = 32'h8220000;
      35387: inst = 32'h10408000;
      35388: inst = 32'hc404c59;
      35389: inst = 32'h8220000;
      35390: inst = 32'h10408000;
      35391: inst = 32'hc404c5a;
      35392: inst = 32'h8220000;
      35393: inst = 32'h10408000;
      35394: inst = 32'hc404c5b;
      35395: inst = 32'h8220000;
      35396: inst = 32'h10408000;
      35397: inst = 32'hc404c5c;
      35398: inst = 32'h8220000;
      35399: inst = 32'h10408000;
      35400: inst = 32'hc404c5d;
      35401: inst = 32'h8220000;
      35402: inst = 32'h10408000;
      35403: inst = 32'hc404c5e;
      35404: inst = 32'h8220000;
      35405: inst = 32'h10408000;
      35406: inst = 32'hc404c5f;
      35407: inst = 32'h8220000;
      35408: inst = 32'h10408000;
      35409: inst = 32'hc404c60;
      35410: inst = 32'h8220000;
      35411: inst = 32'h10408000;
      35412: inst = 32'hc404c61;
      35413: inst = 32'h8220000;
      35414: inst = 32'h10408000;
      35415: inst = 32'hc404c62;
      35416: inst = 32'h8220000;
      35417: inst = 32'h10408000;
      35418: inst = 32'hc404c63;
      35419: inst = 32'h8220000;
      35420: inst = 32'h10408000;
      35421: inst = 32'hc404c64;
      35422: inst = 32'h8220000;
      35423: inst = 32'h10408000;
      35424: inst = 32'hc404c65;
      35425: inst = 32'h8220000;
      35426: inst = 32'h10408000;
      35427: inst = 32'hc404c66;
      35428: inst = 32'h8220000;
      35429: inst = 32'h10408000;
      35430: inst = 32'hc404c67;
      35431: inst = 32'h8220000;
      35432: inst = 32'h10408000;
      35433: inst = 32'hc404c68;
      35434: inst = 32'h8220000;
      35435: inst = 32'h10408000;
      35436: inst = 32'hc404c69;
      35437: inst = 32'h8220000;
      35438: inst = 32'h10408000;
      35439: inst = 32'hc404c6a;
      35440: inst = 32'h8220000;
      35441: inst = 32'h10408000;
      35442: inst = 32'hc404c6b;
      35443: inst = 32'h8220000;
      35444: inst = 32'h10408000;
      35445: inst = 32'hc404c6c;
      35446: inst = 32'h8220000;
      35447: inst = 32'h10408000;
      35448: inst = 32'hc404c6d;
      35449: inst = 32'h8220000;
      35450: inst = 32'h10408000;
      35451: inst = 32'hc404c6e;
      35452: inst = 32'h8220000;
      35453: inst = 32'h10408000;
      35454: inst = 32'hc404c6f;
      35455: inst = 32'h8220000;
      35456: inst = 32'h10408000;
      35457: inst = 32'hc404c70;
      35458: inst = 32'h8220000;
      35459: inst = 32'h10408000;
      35460: inst = 32'hc404c71;
      35461: inst = 32'h8220000;
      35462: inst = 32'h10408000;
      35463: inst = 32'hc404c72;
      35464: inst = 32'h8220000;
      35465: inst = 32'h10408000;
      35466: inst = 32'hc404c73;
      35467: inst = 32'h8220000;
      35468: inst = 32'h10408000;
      35469: inst = 32'hc404c74;
      35470: inst = 32'h8220000;
      35471: inst = 32'h10408000;
      35472: inst = 32'hc404c75;
      35473: inst = 32'h8220000;
      35474: inst = 32'h10408000;
      35475: inst = 32'hc404c76;
      35476: inst = 32'h8220000;
      35477: inst = 32'h10408000;
      35478: inst = 32'hc404c77;
      35479: inst = 32'h8220000;
      35480: inst = 32'h10408000;
      35481: inst = 32'hc404c78;
      35482: inst = 32'h8220000;
      35483: inst = 32'h10408000;
      35484: inst = 32'hc404c79;
      35485: inst = 32'h8220000;
      35486: inst = 32'h10408000;
      35487: inst = 32'hc404c7a;
      35488: inst = 32'h8220000;
      35489: inst = 32'h10408000;
      35490: inst = 32'hc404c7b;
      35491: inst = 32'h8220000;
      35492: inst = 32'h10408000;
      35493: inst = 32'hc404c7c;
      35494: inst = 32'h8220000;
      35495: inst = 32'h10408000;
      35496: inst = 32'hc404c7d;
      35497: inst = 32'h8220000;
      35498: inst = 32'h10408000;
      35499: inst = 32'hc404c7e;
      35500: inst = 32'h8220000;
      35501: inst = 32'h10408000;
      35502: inst = 32'hc404c7f;
      35503: inst = 32'h8220000;
      35504: inst = 32'h10408000;
      35505: inst = 32'hc404c80;
      35506: inst = 32'h8220000;
      35507: inst = 32'h10408000;
      35508: inst = 32'hc404c81;
      35509: inst = 32'h8220000;
      35510: inst = 32'h10408000;
      35511: inst = 32'hc404c82;
      35512: inst = 32'h8220000;
      35513: inst = 32'h10408000;
      35514: inst = 32'hc404c83;
      35515: inst = 32'h8220000;
      35516: inst = 32'h10408000;
      35517: inst = 32'hc404c84;
      35518: inst = 32'h8220000;
      35519: inst = 32'h10408000;
      35520: inst = 32'hc404c85;
      35521: inst = 32'h8220000;
      35522: inst = 32'h10408000;
      35523: inst = 32'hc404c86;
      35524: inst = 32'h8220000;
      35525: inst = 32'h10408000;
      35526: inst = 32'hc404c87;
      35527: inst = 32'h8220000;
      35528: inst = 32'h10408000;
      35529: inst = 32'hc404c88;
      35530: inst = 32'h8220000;
      35531: inst = 32'h10408000;
      35532: inst = 32'hc404c89;
      35533: inst = 32'h8220000;
      35534: inst = 32'h10408000;
      35535: inst = 32'hc404c8a;
      35536: inst = 32'h8220000;
      35537: inst = 32'h10408000;
      35538: inst = 32'hc404c8b;
      35539: inst = 32'h8220000;
      35540: inst = 32'h10408000;
      35541: inst = 32'hc404c8c;
      35542: inst = 32'h8220000;
      35543: inst = 32'h10408000;
      35544: inst = 32'hc404c8d;
      35545: inst = 32'h8220000;
      35546: inst = 32'h10408000;
      35547: inst = 32'hc404c8e;
      35548: inst = 32'h8220000;
      35549: inst = 32'h10408000;
      35550: inst = 32'hc404c8f;
      35551: inst = 32'h8220000;
      35552: inst = 32'h10408000;
      35553: inst = 32'hc404c90;
      35554: inst = 32'h8220000;
      35555: inst = 32'h10408000;
      35556: inst = 32'hc404c91;
      35557: inst = 32'h8220000;
      35558: inst = 32'h10408000;
      35559: inst = 32'hc404c92;
      35560: inst = 32'h8220000;
      35561: inst = 32'h10408000;
      35562: inst = 32'hc404c93;
      35563: inst = 32'h8220000;
      35564: inst = 32'h10408000;
      35565: inst = 32'hc404c94;
      35566: inst = 32'h8220000;
      35567: inst = 32'h10408000;
      35568: inst = 32'hc404c95;
      35569: inst = 32'h8220000;
      35570: inst = 32'h10408000;
      35571: inst = 32'hc404c96;
      35572: inst = 32'h8220000;
      35573: inst = 32'h10408000;
      35574: inst = 32'hc404c97;
      35575: inst = 32'h8220000;
      35576: inst = 32'h10408000;
      35577: inst = 32'hc404c98;
      35578: inst = 32'h8220000;
      35579: inst = 32'h10408000;
      35580: inst = 32'hc404c99;
      35581: inst = 32'h8220000;
      35582: inst = 32'h10408000;
      35583: inst = 32'hc404c9a;
      35584: inst = 32'h8220000;
      35585: inst = 32'h10408000;
      35586: inst = 32'hc404c9b;
      35587: inst = 32'h8220000;
      35588: inst = 32'h10408000;
      35589: inst = 32'hc404c9c;
      35590: inst = 32'h8220000;
      35591: inst = 32'h10408000;
      35592: inst = 32'hc404ca3;
      35593: inst = 32'h8220000;
      35594: inst = 32'h10408000;
      35595: inst = 32'hc404ca4;
      35596: inst = 32'h8220000;
      35597: inst = 32'h10408000;
      35598: inst = 32'hc404ca5;
      35599: inst = 32'h8220000;
      35600: inst = 32'h10408000;
      35601: inst = 32'hc404ca6;
      35602: inst = 32'h8220000;
      35603: inst = 32'h10408000;
      35604: inst = 32'hc404ca7;
      35605: inst = 32'h8220000;
      35606: inst = 32'h10408000;
      35607: inst = 32'hc404ca8;
      35608: inst = 32'h8220000;
      35609: inst = 32'h10408000;
      35610: inst = 32'hc404ca9;
      35611: inst = 32'h8220000;
      35612: inst = 32'h10408000;
      35613: inst = 32'hc404caa;
      35614: inst = 32'h8220000;
      35615: inst = 32'h10408000;
      35616: inst = 32'hc404cab;
      35617: inst = 32'h8220000;
      35618: inst = 32'h10408000;
      35619: inst = 32'hc404cac;
      35620: inst = 32'h8220000;
      35621: inst = 32'h10408000;
      35622: inst = 32'hc404cad;
      35623: inst = 32'h8220000;
      35624: inst = 32'h10408000;
      35625: inst = 32'hc404cae;
      35626: inst = 32'h8220000;
      35627: inst = 32'h10408000;
      35628: inst = 32'hc404caf;
      35629: inst = 32'h8220000;
      35630: inst = 32'h10408000;
      35631: inst = 32'hc404cb0;
      35632: inst = 32'h8220000;
      35633: inst = 32'h10408000;
      35634: inst = 32'hc404cb1;
      35635: inst = 32'h8220000;
      35636: inst = 32'h10408000;
      35637: inst = 32'hc404cb2;
      35638: inst = 32'h8220000;
      35639: inst = 32'h10408000;
      35640: inst = 32'hc404cb3;
      35641: inst = 32'h8220000;
      35642: inst = 32'h10408000;
      35643: inst = 32'hc404cb4;
      35644: inst = 32'h8220000;
      35645: inst = 32'h10408000;
      35646: inst = 32'hc404cb5;
      35647: inst = 32'h8220000;
      35648: inst = 32'h10408000;
      35649: inst = 32'hc404cb6;
      35650: inst = 32'h8220000;
      35651: inst = 32'h10408000;
      35652: inst = 32'hc404cb7;
      35653: inst = 32'h8220000;
      35654: inst = 32'h10408000;
      35655: inst = 32'hc404cb8;
      35656: inst = 32'h8220000;
      35657: inst = 32'h10408000;
      35658: inst = 32'hc404cb9;
      35659: inst = 32'h8220000;
      35660: inst = 32'h10408000;
      35661: inst = 32'hc404cba;
      35662: inst = 32'h8220000;
      35663: inst = 32'h10408000;
      35664: inst = 32'hc404cbb;
      35665: inst = 32'h8220000;
      35666: inst = 32'h10408000;
      35667: inst = 32'hc404cbc;
      35668: inst = 32'h8220000;
      35669: inst = 32'h10408000;
      35670: inst = 32'hc404cbd;
      35671: inst = 32'h8220000;
      35672: inst = 32'h10408000;
      35673: inst = 32'hc404cbe;
      35674: inst = 32'h8220000;
      35675: inst = 32'h10408000;
      35676: inst = 32'hc404cbf;
      35677: inst = 32'h8220000;
      35678: inst = 32'h10408000;
      35679: inst = 32'hc404cc0;
      35680: inst = 32'h8220000;
      35681: inst = 32'h10408000;
      35682: inst = 32'hc404cc1;
      35683: inst = 32'h8220000;
      35684: inst = 32'h10408000;
      35685: inst = 32'hc404cc2;
      35686: inst = 32'h8220000;
      35687: inst = 32'h10408000;
      35688: inst = 32'hc404cc3;
      35689: inst = 32'h8220000;
      35690: inst = 32'h10408000;
      35691: inst = 32'hc404cc4;
      35692: inst = 32'h8220000;
      35693: inst = 32'h10408000;
      35694: inst = 32'hc404cc5;
      35695: inst = 32'h8220000;
      35696: inst = 32'h10408000;
      35697: inst = 32'hc404cc6;
      35698: inst = 32'h8220000;
      35699: inst = 32'h10408000;
      35700: inst = 32'hc404cc7;
      35701: inst = 32'h8220000;
      35702: inst = 32'h10408000;
      35703: inst = 32'hc404cc8;
      35704: inst = 32'h8220000;
      35705: inst = 32'h10408000;
      35706: inst = 32'hc404cc9;
      35707: inst = 32'h8220000;
      35708: inst = 32'h10408000;
      35709: inst = 32'hc404cca;
      35710: inst = 32'h8220000;
      35711: inst = 32'h10408000;
      35712: inst = 32'hc404ccb;
      35713: inst = 32'h8220000;
      35714: inst = 32'h10408000;
      35715: inst = 32'hc404ccc;
      35716: inst = 32'h8220000;
      35717: inst = 32'h10408000;
      35718: inst = 32'hc404ccd;
      35719: inst = 32'h8220000;
      35720: inst = 32'h10408000;
      35721: inst = 32'hc404cce;
      35722: inst = 32'h8220000;
      35723: inst = 32'h10408000;
      35724: inst = 32'hc404ccf;
      35725: inst = 32'h8220000;
      35726: inst = 32'h10408000;
      35727: inst = 32'hc404cd0;
      35728: inst = 32'h8220000;
      35729: inst = 32'h10408000;
      35730: inst = 32'hc404cd1;
      35731: inst = 32'h8220000;
      35732: inst = 32'h10408000;
      35733: inst = 32'hc404cd2;
      35734: inst = 32'h8220000;
      35735: inst = 32'h10408000;
      35736: inst = 32'hc404cd3;
      35737: inst = 32'h8220000;
      35738: inst = 32'h10408000;
      35739: inst = 32'hc404cd4;
      35740: inst = 32'h8220000;
      35741: inst = 32'h10408000;
      35742: inst = 32'hc404cd5;
      35743: inst = 32'h8220000;
      35744: inst = 32'h10408000;
      35745: inst = 32'hc404cd6;
      35746: inst = 32'h8220000;
      35747: inst = 32'h10408000;
      35748: inst = 32'hc404cd7;
      35749: inst = 32'h8220000;
      35750: inst = 32'h10408000;
      35751: inst = 32'hc404cd8;
      35752: inst = 32'h8220000;
      35753: inst = 32'h10408000;
      35754: inst = 32'hc404cd9;
      35755: inst = 32'h8220000;
      35756: inst = 32'h10408000;
      35757: inst = 32'hc404cda;
      35758: inst = 32'h8220000;
      35759: inst = 32'h10408000;
      35760: inst = 32'hc404cdb;
      35761: inst = 32'h8220000;
      35762: inst = 32'h10408000;
      35763: inst = 32'hc404cdc;
      35764: inst = 32'h8220000;
      35765: inst = 32'h10408000;
      35766: inst = 32'hc404cdd;
      35767: inst = 32'h8220000;
      35768: inst = 32'h10408000;
      35769: inst = 32'hc404cde;
      35770: inst = 32'h8220000;
      35771: inst = 32'h10408000;
      35772: inst = 32'hc404cdf;
      35773: inst = 32'h8220000;
      35774: inst = 32'h10408000;
      35775: inst = 32'hc404ce0;
      35776: inst = 32'h8220000;
      35777: inst = 32'h10408000;
      35778: inst = 32'hc404ce1;
      35779: inst = 32'h8220000;
      35780: inst = 32'h10408000;
      35781: inst = 32'hc404ce2;
      35782: inst = 32'h8220000;
      35783: inst = 32'h10408000;
      35784: inst = 32'hc404ce3;
      35785: inst = 32'h8220000;
      35786: inst = 32'h10408000;
      35787: inst = 32'hc404ce4;
      35788: inst = 32'h8220000;
      35789: inst = 32'h10408000;
      35790: inst = 32'hc404ce5;
      35791: inst = 32'h8220000;
      35792: inst = 32'h10408000;
      35793: inst = 32'hc404ce6;
      35794: inst = 32'h8220000;
      35795: inst = 32'h10408000;
      35796: inst = 32'hc404ce7;
      35797: inst = 32'h8220000;
      35798: inst = 32'h10408000;
      35799: inst = 32'hc404ce8;
      35800: inst = 32'h8220000;
      35801: inst = 32'h10408000;
      35802: inst = 32'hc404ce9;
      35803: inst = 32'h8220000;
      35804: inst = 32'h10408000;
      35805: inst = 32'hc404cea;
      35806: inst = 32'h8220000;
      35807: inst = 32'h10408000;
      35808: inst = 32'hc404ceb;
      35809: inst = 32'h8220000;
      35810: inst = 32'h10408000;
      35811: inst = 32'hc404cec;
      35812: inst = 32'h8220000;
      35813: inst = 32'h10408000;
      35814: inst = 32'hc404ced;
      35815: inst = 32'h8220000;
      35816: inst = 32'h10408000;
      35817: inst = 32'hc404cee;
      35818: inst = 32'h8220000;
      35819: inst = 32'h10408000;
      35820: inst = 32'hc404cef;
      35821: inst = 32'h8220000;
      35822: inst = 32'h10408000;
      35823: inst = 32'hc404cf0;
      35824: inst = 32'h8220000;
      35825: inst = 32'h10408000;
      35826: inst = 32'hc404cf1;
      35827: inst = 32'h8220000;
      35828: inst = 32'h10408000;
      35829: inst = 32'hc404cf2;
      35830: inst = 32'h8220000;
      35831: inst = 32'h10408000;
      35832: inst = 32'hc404cf3;
      35833: inst = 32'h8220000;
      35834: inst = 32'h10408000;
      35835: inst = 32'hc404cf4;
      35836: inst = 32'h8220000;
      35837: inst = 32'h10408000;
      35838: inst = 32'hc404cf5;
      35839: inst = 32'h8220000;
      35840: inst = 32'h10408000;
      35841: inst = 32'hc404cf6;
      35842: inst = 32'h8220000;
      35843: inst = 32'h10408000;
      35844: inst = 32'hc404cf7;
      35845: inst = 32'h8220000;
      35846: inst = 32'h10408000;
      35847: inst = 32'hc404cf8;
      35848: inst = 32'h8220000;
      35849: inst = 32'h10408000;
      35850: inst = 32'hc404cf9;
      35851: inst = 32'h8220000;
      35852: inst = 32'h10408000;
      35853: inst = 32'hc404cfa;
      35854: inst = 32'h8220000;
      35855: inst = 32'h10408000;
      35856: inst = 32'hc404cfb;
      35857: inst = 32'h8220000;
      35858: inst = 32'h10408000;
      35859: inst = 32'hc404cfc;
      35860: inst = 32'h8220000;
      35861: inst = 32'h10408000;
      35862: inst = 32'hc404d03;
      35863: inst = 32'h8220000;
      35864: inst = 32'h10408000;
      35865: inst = 32'hc404d04;
      35866: inst = 32'h8220000;
      35867: inst = 32'h10408000;
      35868: inst = 32'hc404d05;
      35869: inst = 32'h8220000;
      35870: inst = 32'h10408000;
      35871: inst = 32'hc404d06;
      35872: inst = 32'h8220000;
      35873: inst = 32'h10408000;
      35874: inst = 32'hc404d07;
      35875: inst = 32'h8220000;
      35876: inst = 32'h10408000;
      35877: inst = 32'hc404d08;
      35878: inst = 32'h8220000;
      35879: inst = 32'h10408000;
      35880: inst = 32'hc404d09;
      35881: inst = 32'h8220000;
      35882: inst = 32'h10408000;
      35883: inst = 32'hc404d0a;
      35884: inst = 32'h8220000;
      35885: inst = 32'h10408000;
      35886: inst = 32'hc404d0b;
      35887: inst = 32'h8220000;
      35888: inst = 32'h10408000;
      35889: inst = 32'hc404d0c;
      35890: inst = 32'h8220000;
      35891: inst = 32'h10408000;
      35892: inst = 32'hc404d0d;
      35893: inst = 32'h8220000;
      35894: inst = 32'h10408000;
      35895: inst = 32'hc404d0e;
      35896: inst = 32'h8220000;
      35897: inst = 32'h10408000;
      35898: inst = 32'hc404d0f;
      35899: inst = 32'h8220000;
      35900: inst = 32'h10408000;
      35901: inst = 32'hc404d10;
      35902: inst = 32'h8220000;
      35903: inst = 32'h10408000;
      35904: inst = 32'hc404d11;
      35905: inst = 32'h8220000;
      35906: inst = 32'h10408000;
      35907: inst = 32'hc404d12;
      35908: inst = 32'h8220000;
      35909: inst = 32'h10408000;
      35910: inst = 32'hc404d13;
      35911: inst = 32'h8220000;
      35912: inst = 32'h10408000;
      35913: inst = 32'hc404d14;
      35914: inst = 32'h8220000;
      35915: inst = 32'h10408000;
      35916: inst = 32'hc404d15;
      35917: inst = 32'h8220000;
      35918: inst = 32'h10408000;
      35919: inst = 32'hc404d16;
      35920: inst = 32'h8220000;
      35921: inst = 32'h10408000;
      35922: inst = 32'hc404d17;
      35923: inst = 32'h8220000;
      35924: inst = 32'h10408000;
      35925: inst = 32'hc404d18;
      35926: inst = 32'h8220000;
      35927: inst = 32'h10408000;
      35928: inst = 32'hc404d19;
      35929: inst = 32'h8220000;
      35930: inst = 32'h10408000;
      35931: inst = 32'hc404d1a;
      35932: inst = 32'h8220000;
      35933: inst = 32'h10408000;
      35934: inst = 32'hc404d1b;
      35935: inst = 32'h8220000;
      35936: inst = 32'h10408000;
      35937: inst = 32'hc404d1c;
      35938: inst = 32'h8220000;
      35939: inst = 32'h10408000;
      35940: inst = 32'hc404d1d;
      35941: inst = 32'h8220000;
      35942: inst = 32'h10408000;
      35943: inst = 32'hc404d1e;
      35944: inst = 32'h8220000;
      35945: inst = 32'h10408000;
      35946: inst = 32'hc404d1f;
      35947: inst = 32'h8220000;
      35948: inst = 32'h10408000;
      35949: inst = 32'hc404d20;
      35950: inst = 32'h8220000;
      35951: inst = 32'h10408000;
      35952: inst = 32'hc404d21;
      35953: inst = 32'h8220000;
      35954: inst = 32'h10408000;
      35955: inst = 32'hc404d22;
      35956: inst = 32'h8220000;
      35957: inst = 32'h10408000;
      35958: inst = 32'hc404d23;
      35959: inst = 32'h8220000;
      35960: inst = 32'h10408000;
      35961: inst = 32'hc404d24;
      35962: inst = 32'h8220000;
      35963: inst = 32'h10408000;
      35964: inst = 32'hc404d3b;
      35965: inst = 32'h8220000;
      35966: inst = 32'h10408000;
      35967: inst = 32'hc404d3c;
      35968: inst = 32'h8220000;
      35969: inst = 32'h10408000;
      35970: inst = 32'hc404d3d;
      35971: inst = 32'h8220000;
      35972: inst = 32'h10408000;
      35973: inst = 32'hc404d3e;
      35974: inst = 32'h8220000;
      35975: inst = 32'h10408000;
      35976: inst = 32'hc404d3f;
      35977: inst = 32'h8220000;
      35978: inst = 32'h10408000;
      35979: inst = 32'hc404d40;
      35980: inst = 32'h8220000;
      35981: inst = 32'h10408000;
      35982: inst = 32'hc404d41;
      35983: inst = 32'h8220000;
      35984: inst = 32'h10408000;
      35985: inst = 32'hc404d42;
      35986: inst = 32'h8220000;
      35987: inst = 32'h10408000;
      35988: inst = 32'hc404d43;
      35989: inst = 32'h8220000;
      35990: inst = 32'h10408000;
      35991: inst = 32'hc404d44;
      35992: inst = 32'h8220000;
      35993: inst = 32'h10408000;
      35994: inst = 32'hc404d45;
      35995: inst = 32'h8220000;
      35996: inst = 32'h10408000;
      35997: inst = 32'hc404d46;
      35998: inst = 32'h8220000;
      35999: inst = 32'h10408000;
      36000: inst = 32'hc404d47;
      36001: inst = 32'h8220000;
      36002: inst = 32'h10408000;
      36003: inst = 32'hc404d48;
      36004: inst = 32'h8220000;
      36005: inst = 32'h10408000;
      36006: inst = 32'hc404d49;
      36007: inst = 32'h8220000;
      36008: inst = 32'h10408000;
      36009: inst = 32'hc404d4a;
      36010: inst = 32'h8220000;
      36011: inst = 32'h10408000;
      36012: inst = 32'hc404d4b;
      36013: inst = 32'h8220000;
      36014: inst = 32'h10408000;
      36015: inst = 32'hc404d4c;
      36016: inst = 32'h8220000;
      36017: inst = 32'h10408000;
      36018: inst = 32'hc404d4d;
      36019: inst = 32'h8220000;
      36020: inst = 32'h10408000;
      36021: inst = 32'hc404d4e;
      36022: inst = 32'h8220000;
      36023: inst = 32'h10408000;
      36024: inst = 32'hc404d4f;
      36025: inst = 32'h8220000;
      36026: inst = 32'h10408000;
      36027: inst = 32'hc404d50;
      36028: inst = 32'h8220000;
      36029: inst = 32'h10408000;
      36030: inst = 32'hc404d51;
      36031: inst = 32'h8220000;
      36032: inst = 32'h10408000;
      36033: inst = 32'hc404d52;
      36034: inst = 32'h8220000;
      36035: inst = 32'h10408000;
      36036: inst = 32'hc404d53;
      36037: inst = 32'h8220000;
      36038: inst = 32'h10408000;
      36039: inst = 32'hc404d54;
      36040: inst = 32'h8220000;
      36041: inst = 32'h10408000;
      36042: inst = 32'hc404d55;
      36043: inst = 32'h8220000;
      36044: inst = 32'h10408000;
      36045: inst = 32'hc404d56;
      36046: inst = 32'h8220000;
      36047: inst = 32'h10408000;
      36048: inst = 32'hc404d57;
      36049: inst = 32'h8220000;
      36050: inst = 32'h10408000;
      36051: inst = 32'hc404d58;
      36052: inst = 32'h8220000;
      36053: inst = 32'h10408000;
      36054: inst = 32'hc404d59;
      36055: inst = 32'h8220000;
      36056: inst = 32'h10408000;
      36057: inst = 32'hc404d5a;
      36058: inst = 32'h8220000;
      36059: inst = 32'h10408000;
      36060: inst = 32'hc404d5b;
      36061: inst = 32'h8220000;
      36062: inst = 32'h10408000;
      36063: inst = 32'hc404d5c;
      36064: inst = 32'h8220000;
      36065: inst = 32'h10408000;
      36066: inst = 32'hc404d63;
      36067: inst = 32'h8220000;
      36068: inst = 32'h10408000;
      36069: inst = 32'hc404d64;
      36070: inst = 32'h8220000;
      36071: inst = 32'h10408000;
      36072: inst = 32'hc404d65;
      36073: inst = 32'h8220000;
      36074: inst = 32'h10408000;
      36075: inst = 32'hc404d66;
      36076: inst = 32'h8220000;
      36077: inst = 32'h10408000;
      36078: inst = 32'hc404d67;
      36079: inst = 32'h8220000;
      36080: inst = 32'h10408000;
      36081: inst = 32'hc404d68;
      36082: inst = 32'h8220000;
      36083: inst = 32'h10408000;
      36084: inst = 32'hc404d69;
      36085: inst = 32'h8220000;
      36086: inst = 32'h10408000;
      36087: inst = 32'hc404d6a;
      36088: inst = 32'h8220000;
      36089: inst = 32'h10408000;
      36090: inst = 32'hc404d6b;
      36091: inst = 32'h8220000;
      36092: inst = 32'h10408000;
      36093: inst = 32'hc404d6c;
      36094: inst = 32'h8220000;
      36095: inst = 32'h10408000;
      36096: inst = 32'hc404d6d;
      36097: inst = 32'h8220000;
      36098: inst = 32'h10408000;
      36099: inst = 32'hc404d6e;
      36100: inst = 32'h8220000;
      36101: inst = 32'h10408000;
      36102: inst = 32'hc404d6f;
      36103: inst = 32'h8220000;
      36104: inst = 32'h10408000;
      36105: inst = 32'hc404d70;
      36106: inst = 32'h8220000;
      36107: inst = 32'h10408000;
      36108: inst = 32'hc404d71;
      36109: inst = 32'h8220000;
      36110: inst = 32'h10408000;
      36111: inst = 32'hc404d72;
      36112: inst = 32'h8220000;
      36113: inst = 32'h10408000;
      36114: inst = 32'hc404d73;
      36115: inst = 32'h8220000;
      36116: inst = 32'h10408000;
      36117: inst = 32'hc404d74;
      36118: inst = 32'h8220000;
      36119: inst = 32'h10408000;
      36120: inst = 32'hc404d75;
      36121: inst = 32'h8220000;
      36122: inst = 32'h10408000;
      36123: inst = 32'hc404d76;
      36124: inst = 32'h8220000;
      36125: inst = 32'h10408000;
      36126: inst = 32'hc404d77;
      36127: inst = 32'h8220000;
      36128: inst = 32'h10408000;
      36129: inst = 32'hc404d78;
      36130: inst = 32'h8220000;
      36131: inst = 32'h10408000;
      36132: inst = 32'hc404d79;
      36133: inst = 32'h8220000;
      36134: inst = 32'h10408000;
      36135: inst = 32'hc404d7a;
      36136: inst = 32'h8220000;
      36137: inst = 32'h10408000;
      36138: inst = 32'hc404d7b;
      36139: inst = 32'h8220000;
      36140: inst = 32'h10408000;
      36141: inst = 32'hc404d7c;
      36142: inst = 32'h8220000;
      36143: inst = 32'h10408000;
      36144: inst = 32'hc404d7d;
      36145: inst = 32'h8220000;
      36146: inst = 32'h10408000;
      36147: inst = 32'hc404d7e;
      36148: inst = 32'h8220000;
      36149: inst = 32'h10408000;
      36150: inst = 32'hc404d7f;
      36151: inst = 32'h8220000;
      36152: inst = 32'h10408000;
      36153: inst = 32'hc404d80;
      36154: inst = 32'h8220000;
      36155: inst = 32'h10408000;
      36156: inst = 32'hc404d81;
      36157: inst = 32'h8220000;
      36158: inst = 32'h10408000;
      36159: inst = 32'hc404d82;
      36160: inst = 32'h8220000;
      36161: inst = 32'h10408000;
      36162: inst = 32'hc404d83;
      36163: inst = 32'h8220000;
      36164: inst = 32'h10408000;
      36165: inst = 32'hc404d84;
      36166: inst = 32'h8220000;
      36167: inst = 32'h10408000;
      36168: inst = 32'hc404d9b;
      36169: inst = 32'h8220000;
      36170: inst = 32'h10408000;
      36171: inst = 32'hc404d9c;
      36172: inst = 32'h8220000;
      36173: inst = 32'h10408000;
      36174: inst = 32'hc404d9d;
      36175: inst = 32'h8220000;
      36176: inst = 32'h10408000;
      36177: inst = 32'hc404d9e;
      36178: inst = 32'h8220000;
      36179: inst = 32'h10408000;
      36180: inst = 32'hc404d9f;
      36181: inst = 32'h8220000;
      36182: inst = 32'h10408000;
      36183: inst = 32'hc404da0;
      36184: inst = 32'h8220000;
      36185: inst = 32'h10408000;
      36186: inst = 32'hc404da1;
      36187: inst = 32'h8220000;
      36188: inst = 32'h10408000;
      36189: inst = 32'hc404da2;
      36190: inst = 32'h8220000;
      36191: inst = 32'h10408000;
      36192: inst = 32'hc404da3;
      36193: inst = 32'h8220000;
      36194: inst = 32'h10408000;
      36195: inst = 32'hc404da4;
      36196: inst = 32'h8220000;
      36197: inst = 32'h10408000;
      36198: inst = 32'hc404da5;
      36199: inst = 32'h8220000;
      36200: inst = 32'h10408000;
      36201: inst = 32'hc404da6;
      36202: inst = 32'h8220000;
      36203: inst = 32'h10408000;
      36204: inst = 32'hc404da7;
      36205: inst = 32'h8220000;
      36206: inst = 32'h10408000;
      36207: inst = 32'hc404da8;
      36208: inst = 32'h8220000;
      36209: inst = 32'h10408000;
      36210: inst = 32'hc404da9;
      36211: inst = 32'h8220000;
      36212: inst = 32'h10408000;
      36213: inst = 32'hc404daa;
      36214: inst = 32'h8220000;
      36215: inst = 32'h10408000;
      36216: inst = 32'hc404dab;
      36217: inst = 32'h8220000;
      36218: inst = 32'h10408000;
      36219: inst = 32'hc404dac;
      36220: inst = 32'h8220000;
      36221: inst = 32'h10408000;
      36222: inst = 32'hc404dad;
      36223: inst = 32'h8220000;
      36224: inst = 32'h10408000;
      36225: inst = 32'hc404dae;
      36226: inst = 32'h8220000;
      36227: inst = 32'h10408000;
      36228: inst = 32'hc404daf;
      36229: inst = 32'h8220000;
      36230: inst = 32'h10408000;
      36231: inst = 32'hc404db0;
      36232: inst = 32'h8220000;
      36233: inst = 32'h10408000;
      36234: inst = 32'hc404db1;
      36235: inst = 32'h8220000;
      36236: inst = 32'h10408000;
      36237: inst = 32'hc404db2;
      36238: inst = 32'h8220000;
      36239: inst = 32'h10408000;
      36240: inst = 32'hc404db3;
      36241: inst = 32'h8220000;
      36242: inst = 32'h10408000;
      36243: inst = 32'hc404db4;
      36244: inst = 32'h8220000;
      36245: inst = 32'h10408000;
      36246: inst = 32'hc404db5;
      36247: inst = 32'h8220000;
      36248: inst = 32'h10408000;
      36249: inst = 32'hc404db6;
      36250: inst = 32'h8220000;
      36251: inst = 32'h10408000;
      36252: inst = 32'hc404db7;
      36253: inst = 32'h8220000;
      36254: inst = 32'h10408000;
      36255: inst = 32'hc404db8;
      36256: inst = 32'h8220000;
      36257: inst = 32'h10408000;
      36258: inst = 32'hc404db9;
      36259: inst = 32'h8220000;
      36260: inst = 32'h10408000;
      36261: inst = 32'hc404dba;
      36262: inst = 32'h8220000;
      36263: inst = 32'h10408000;
      36264: inst = 32'hc404dbb;
      36265: inst = 32'h8220000;
      36266: inst = 32'h10408000;
      36267: inst = 32'hc404dbc;
      36268: inst = 32'h8220000;
      36269: inst = 32'h10408000;
      36270: inst = 32'hc404dc3;
      36271: inst = 32'h8220000;
      36272: inst = 32'h10408000;
      36273: inst = 32'hc404dc4;
      36274: inst = 32'h8220000;
      36275: inst = 32'h10408000;
      36276: inst = 32'hc404dc5;
      36277: inst = 32'h8220000;
      36278: inst = 32'h10408000;
      36279: inst = 32'hc404dc6;
      36280: inst = 32'h8220000;
      36281: inst = 32'h10408000;
      36282: inst = 32'hc404dc7;
      36283: inst = 32'h8220000;
      36284: inst = 32'h10408000;
      36285: inst = 32'hc404dc8;
      36286: inst = 32'h8220000;
      36287: inst = 32'h10408000;
      36288: inst = 32'hc404dc9;
      36289: inst = 32'h8220000;
      36290: inst = 32'h10408000;
      36291: inst = 32'hc404dca;
      36292: inst = 32'h8220000;
      36293: inst = 32'h10408000;
      36294: inst = 32'hc404dcb;
      36295: inst = 32'h8220000;
      36296: inst = 32'h10408000;
      36297: inst = 32'hc404dcc;
      36298: inst = 32'h8220000;
      36299: inst = 32'h10408000;
      36300: inst = 32'hc404dcd;
      36301: inst = 32'h8220000;
      36302: inst = 32'h10408000;
      36303: inst = 32'hc404dce;
      36304: inst = 32'h8220000;
      36305: inst = 32'h10408000;
      36306: inst = 32'hc404dcf;
      36307: inst = 32'h8220000;
      36308: inst = 32'h10408000;
      36309: inst = 32'hc404dd0;
      36310: inst = 32'h8220000;
      36311: inst = 32'h10408000;
      36312: inst = 32'hc404dd1;
      36313: inst = 32'h8220000;
      36314: inst = 32'h10408000;
      36315: inst = 32'hc404dd2;
      36316: inst = 32'h8220000;
      36317: inst = 32'h10408000;
      36318: inst = 32'hc404dd3;
      36319: inst = 32'h8220000;
      36320: inst = 32'h10408000;
      36321: inst = 32'hc404dd4;
      36322: inst = 32'h8220000;
      36323: inst = 32'h10408000;
      36324: inst = 32'hc404dd5;
      36325: inst = 32'h8220000;
      36326: inst = 32'h10408000;
      36327: inst = 32'hc404dd6;
      36328: inst = 32'h8220000;
      36329: inst = 32'h10408000;
      36330: inst = 32'hc404dd7;
      36331: inst = 32'h8220000;
      36332: inst = 32'h10408000;
      36333: inst = 32'hc404dd8;
      36334: inst = 32'h8220000;
      36335: inst = 32'h10408000;
      36336: inst = 32'hc404dd9;
      36337: inst = 32'h8220000;
      36338: inst = 32'h10408000;
      36339: inst = 32'hc404dda;
      36340: inst = 32'h8220000;
      36341: inst = 32'h10408000;
      36342: inst = 32'hc404ddb;
      36343: inst = 32'h8220000;
      36344: inst = 32'h10408000;
      36345: inst = 32'hc404ddc;
      36346: inst = 32'h8220000;
      36347: inst = 32'h10408000;
      36348: inst = 32'hc404ddd;
      36349: inst = 32'h8220000;
      36350: inst = 32'h10408000;
      36351: inst = 32'hc404dde;
      36352: inst = 32'h8220000;
      36353: inst = 32'h10408000;
      36354: inst = 32'hc404ddf;
      36355: inst = 32'h8220000;
      36356: inst = 32'h10408000;
      36357: inst = 32'hc404de0;
      36358: inst = 32'h8220000;
      36359: inst = 32'h10408000;
      36360: inst = 32'hc404de1;
      36361: inst = 32'h8220000;
      36362: inst = 32'h10408000;
      36363: inst = 32'hc404de2;
      36364: inst = 32'h8220000;
      36365: inst = 32'h10408000;
      36366: inst = 32'hc404de3;
      36367: inst = 32'h8220000;
      36368: inst = 32'h10408000;
      36369: inst = 32'hc404de4;
      36370: inst = 32'h8220000;
      36371: inst = 32'h10408000;
      36372: inst = 32'hc404dfb;
      36373: inst = 32'h8220000;
      36374: inst = 32'h10408000;
      36375: inst = 32'hc404dfc;
      36376: inst = 32'h8220000;
      36377: inst = 32'h10408000;
      36378: inst = 32'hc404dfd;
      36379: inst = 32'h8220000;
      36380: inst = 32'h10408000;
      36381: inst = 32'hc404dfe;
      36382: inst = 32'h8220000;
      36383: inst = 32'h10408000;
      36384: inst = 32'hc404dff;
      36385: inst = 32'h8220000;
      36386: inst = 32'h10408000;
      36387: inst = 32'hc404e00;
      36388: inst = 32'h8220000;
      36389: inst = 32'h10408000;
      36390: inst = 32'hc404e01;
      36391: inst = 32'h8220000;
      36392: inst = 32'h10408000;
      36393: inst = 32'hc404e02;
      36394: inst = 32'h8220000;
      36395: inst = 32'h10408000;
      36396: inst = 32'hc404e03;
      36397: inst = 32'h8220000;
      36398: inst = 32'h10408000;
      36399: inst = 32'hc404e04;
      36400: inst = 32'h8220000;
      36401: inst = 32'h10408000;
      36402: inst = 32'hc404e05;
      36403: inst = 32'h8220000;
      36404: inst = 32'h10408000;
      36405: inst = 32'hc404e06;
      36406: inst = 32'h8220000;
      36407: inst = 32'h10408000;
      36408: inst = 32'hc404e07;
      36409: inst = 32'h8220000;
      36410: inst = 32'h10408000;
      36411: inst = 32'hc404e08;
      36412: inst = 32'h8220000;
      36413: inst = 32'h10408000;
      36414: inst = 32'hc404e09;
      36415: inst = 32'h8220000;
      36416: inst = 32'h10408000;
      36417: inst = 32'hc404e0a;
      36418: inst = 32'h8220000;
      36419: inst = 32'h10408000;
      36420: inst = 32'hc404e0b;
      36421: inst = 32'h8220000;
      36422: inst = 32'h10408000;
      36423: inst = 32'hc404e0c;
      36424: inst = 32'h8220000;
      36425: inst = 32'h10408000;
      36426: inst = 32'hc404e0d;
      36427: inst = 32'h8220000;
      36428: inst = 32'h10408000;
      36429: inst = 32'hc404e0e;
      36430: inst = 32'h8220000;
      36431: inst = 32'h10408000;
      36432: inst = 32'hc404e0f;
      36433: inst = 32'h8220000;
      36434: inst = 32'h10408000;
      36435: inst = 32'hc404e10;
      36436: inst = 32'h8220000;
      36437: inst = 32'h10408000;
      36438: inst = 32'hc404e11;
      36439: inst = 32'h8220000;
      36440: inst = 32'h10408000;
      36441: inst = 32'hc404e12;
      36442: inst = 32'h8220000;
      36443: inst = 32'h10408000;
      36444: inst = 32'hc404e13;
      36445: inst = 32'h8220000;
      36446: inst = 32'h10408000;
      36447: inst = 32'hc404e14;
      36448: inst = 32'h8220000;
      36449: inst = 32'h10408000;
      36450: inst = 32'hc404e15;
      36451: inst = 32'h8220000;
      36452: inst = 32'h10408000;
      36453: inst = 32'hc404e16;
      36454: inst = 32'h8220000;
      36455: inst = 32'h10408000;
      36456: inst = 32'hc404e17;
      36457: inst = 32'h8220000;
      36458: inst = 32'h10408000;
      36459: inst = 32'hc404e18;
      36460: inst = 32'h8220000;
      36461: inst = 32'h10408000;
      36462: inst = 32'hc404e19;
      36463: inst = 32'h8220000;
      36464: inst = 32'h10408000;
      36465: inst = 32'hc404e1a;
      36466: inst = 32'h8220000;
      36467: inst = 32'h10408000;
      36468: inst = 32'hc404e1b;
      36469: inst = 32'h8220000;
      36470: inst = 32'h10408000;
      36471: inst = 32'hc404e1c;
      36472: inst = 32'h8220000;
      36473: inst = 32'h10408000;
      36474: inst = 32'hc404e23;
      36475: inst = 32'h8220000;
      36476: inst = 32'h10408000;
      36477: inst = 32'hc404e24;
      36478: inst = 32'h8220000;
      36479: inst = 32'h10408000;
      36480: inst = 32'hc404e25;
      36481: inst = 32'h8220000;
      36482: inst = 32'h10408000;
      36483: inst = 32'hc404e26;
      36484: inst = 32'h8220000;
      36485: inst = 32'h10408000;
      36486: inst = 32'hc404e27;
      36487: inst = 32'h8220000;
      36488: inst = 32'h10408000;
      36489: inst = 32'hc404e28;
      36490: inst = 32'h8220000;
      36491: inst = 32'h10408000;
      36492: inst = 32'hc404e29;
      36493: inst = 32'h8220000;
      36494: inst = 32'h10408000;
      36495: inst = 32'hc404e2a;
      36496: inst = 32'h8220000;
      36497: inst = 32'h10408000;
      36498: inst = 32'hc404e2b;
      36499: inst = 32'h8220000;
      36500: inst = 32'h10408000;
      36501: inst = 32'hc404e2c;
      36502: inst = 32'h8220000;
      36503: inst = 32'h10408000;
      36504: inst = 32'hc404e2d;
      36505: inst = 32'h8220000;
      36506: inst = 32'h10408000;
      36507: inst = 32'hc404e2e;
      36508: inst = 32'h8220000;
      36509: inst = 32'h10408000;
      36510: inst = 32'hc404e2f;
      36511: inst = 32'h8220000;
      36512: inst = 32'h10408000;
      36513: inst = 32'hc404e30;
      36514: inst = 32'h8220000;
      36515: inst = 32'h10408000;
      36516: inst = 32'hc404e31;
      36517: inst = 32'h8220000;
      36518: inst = 32'h10408000;
      36519: inst = 32'hc404e32;
      36520: inst = 32'h8220000;
      36521: inst = 32'h10408000;
      36522: inst = 32'hc404e33;
      36523: inst = 32'h8220000;
      36524: inst = 32'h10408000;
      36525: inst = 32'hc404e34;
      36526: inst = 32'h8220000;
      36527: inst = 32'h10408000;
      36528: inst = 32'hc404e35;
      36529: inst = 32'h8220000;
      36530: inst = 32'h10408000;
      36531: inst = 32'hc404e36;
      36532: inst = 32'h8220000;
      36533: inst = 32'h10408000;
      36534: inst = 32'hc404e37;
      36535: inst = 32'h8220000;
      36536: inst = 32'h10408000;
      36537: inst = 32'hc404e38;
      36538: inst = 32'h8220000;
      36539: inst = 32'h10408000;
      36540: inst = 32'hc404e39;
      36541: inst = 32'h8220000;
      36542: inst = 32'h10408000;
      36543: inst = 32'hc404e3a;
      36544: inst = 32'h8220000;
      36545: inst = 32'h10408000;
      36546: inst = 32'hc404e3b;
      36547: inst = 32'h8220000;
      36548: inst = 32'h10408000;
      36549: inst = 32'hc404e3c;
      36550: inst = 32'h8220000;
      36551: inst = 32'h10408000;
      36552: inst = 32'hc404e3d;
      36553: inst = 32'h8220000;
      36554: inst = 32'h10408000;
      36555: inst = 32'hc404e3e;
      36556: inst = 32'h8220000;
      36557: inst = 32'h10408000;
      36558: inst = 32'hc404e3f;
      36559: inst = 32'h8220000;
      36560: inst = 32'h10408000;
      36561: inst = 32'hc404e40;
      36562: inst = 32'h8220000;
      36563: inst = 32'h10408000;
      36564: inst = 32'hc404e41;
      36565: inst = 32'h8220000;
      36566: inst = 32'h10408000;
      36567: inst = 32'hc404e42;
      36568: inst = 32'h8220000;
      36569: inst = 32'h10408000;
      36570: inst = 32'hc404e43;
      36571: inst = 32'h8220000;
      36572: inst = 32'h10408000;
      36573: inst = 32'hc404e44;
      36574: inst = 32'h8220000;
      36575: inst = 32'h10408000;
      36576: inst = 32'hc404e45;
      36577: inst = 32'h8220000;
      36578: inst = 32'h10408000;
      36579: inst = 32'hc404e46;
      36580: inst = 32'h8220000;
      36581: inst = 32'h10408000;
      36582: inst = 32'hc404e47;
      36583: inst = 32'h8220000;
      36584: inst = 32'h10408000;
      36585: inst = 32'hc404e48;
      36586: inst = 32'h8220000;
      36587: inst = 32'h10408000;
      36588: inst = 32'hc404e49;
      36589: inst = 32'h8220000;
      36590: inst = 32'h10408000;
      36591: inst = 32'hc404e4a;
      36592: inst = 32'h8220000;
      36593: inst = 32'h10408000;
      36594: inst = 32'hc404e4b;
      36595: inst = 32'h8220000;
      36596: inst = 32'h10408000;
      36597: inst = 32'hc404e4c;
      36598: inst = 32'h8220000;
      36599: inst = 32'h10408000;
      36600: inst = 32'hc404e4d;
      36601: inst = 32'h8220000;
      36602: inst = 32'h10408000;
      36603: inst = 32'hc404e4e;
      36604: inst = 32'h8220000;
      36605: inst = 32'h10408000;
      36606: inst = 32'hc404e4f;
      36607: inst = 32'h8220000;
      36608: inst = 32'h10408000;
      36609: inst = 32'hc404e50;
      36610: inst = 32'h8220000;
      36611: inst = 32'h10408000;
      36612: inst = 32'hc404e51;
      36613: inst = 32'h8220000;
      36614: inst = 32'h10408000;
      36615: inst = 32'hc404e52;
      36616: inst = 32'h8220000;
      36617: inst = 32'h10408000;
      36618: inst = 32'hc404e53;
      36619: inst = 32'h8220000;
      36620: inst = 32'h10408000;
      36621: inst = 32'hc404e54;
      36622: inst = 32'h8220000;
      36623: inst = 32'h10408000;
      36624: inst = 32'hc404e55;
      36625: inst = 32'h8220000;
      36626: inst = 32'h10408000;
      36627: inst = 32'hc404e56;
      36628: inst = 32'h8220000;
      36629: inst = 32'h10408000;
      36630: inst = 32'hc404e57;
      36631: inst = 32'h8220000;
      36632: inst = 32'h10408000;
      36633: inst = 32'hc404e5b;
      36634: inst = 32'h8220000;
      36635: inst = 32'h10408000;
      36636: inst = 32'hc404e5c;
      36637: inst = 32'h8220000;
      36638: inst = 32'h10408000;
      36639: inst = 32'hc404e5d;
      36640: inst = 32'h8220000;
      36641: inst = 32'h10408000;
      36642: inst = 32'hc404e5e;
      36643: inst = 32'h8220000;
      36644: inst = 32'h10408000;
      36645: inst = 32'hc404e5f;
      36646: inst = 32'h8220000;
      36647: inst = 32'h10408000;
      36648: inst = 32'hc404e60;
      36649: inst = 32'h8220000;
      36650: inst = 32'h10408000;
      36651: inst = 32'hc404e61;
      36652: inst = 32'h8220000;
      36653: inst = 32'h10408000;
      36654: inst = 32'hc404e62;
      36655: inst = 32'h8220000;
      36656: inst = 32'h10408000;
      36657: inst = 32'hc404e63;
      36658: inst = 32'h8220000;
      36659: inst = 32'h10408000;
      36660: inst = 32'hc404e64;
      36661: inst = 32'h8220000;
      36662: inst = 32'h10408000;
      36663: inst = 32'hc404e65;
      36664: inst = 32'h8220000;
      36665: inst = 32'h10408000;
      36666: inst = 32'hc404e66;
      36667: inst = 32'h8220000;
      36668: inst = 32'h10408000;
      36669: inst = 32'hc404e67;
      36670: inst = 32'h8220000;
      36671: inst = 32'h10408000;
      36672: inst = 32'hc404e68;
      36673: inst = 32'h8220000;
      36674: inst = 32'h10408000;
      36675: inst = 32'hc404e69;
      36676: inst = 32'h8220000;
      36677: inst = 32'h10408000;
      36678: inst = 32'hc404e6a;
      36679: inst = 32'h8220000;
      36680: inst = 32'h10408000;
      36681: inst = 32'hc404e6b;
      36682: inst = 32'h8220000;
      36683: inst = 32'h10408000;
      36684: inst = 32'hc404e6c;
      36685: inst = 32'h8220000;
      36686: inst = 32'h10408000;
      36687: inst = 32'hc404e6d;
      36688: inst = 32'h8220000;
      36689: inst = 32'h10408000;
      36690: inst = 32'hc404e6e;
      36691: inst = 32'h8220000;
      36692: inst = 32'h10408000;
      36693: inst = 32'hc404e6f;
      36694: inst = 32'h8220000;
      36695: inst = 32'h10408000;
      36696: inst = 32'hc404e70;
      36697: inst = 32'h8220000;
      36698: inst = 32'h10408000;
      36699: inst = 32'hc404e71;
      36700: inst = 32'h8220000;
      36701: inst = 32'h10408000;
      36702: inst = 32'hc404e72;
      36703: inst = 32'h8220000;
      36704: inst = 32'h10408000;
      36705: inst = 32'hc404e73;
      36706: inst = 32'h8220000;
      36707: inst = 32'h10408000;
      36708: inst = 32'hc404e74;
      36709: inst = 32'h8220000;
      36710: inst = 32'h10408000;
      36711: inst = 32'hc404e75;
      36712: inst = 32'h8220000;
      36713: inst = 32'h10408000;
      36714: inst = 32'hc404e76;
      36715: inst = 32'h8220000;
      36716: inst = 32'h10408000;
      36717: inst = 32'hc404e77;
      36718: inst = 32'h8220000;
      36719: inst = 32'h10408000;
      36720: inst = 32'hc404e78;
      36721: inst = 32'h8220000;
      36722: inst = 32'h10408000;
      36723: inst = 32'hc404e79;
      36724: inst = 32'h8220000;
      36725: inst = 32'h10408000;
      36726: inst = 32'hc404e7a;
      36727: inst = 32'h8220000;
      36728: inst = 32'h10408000;
      36729: inst = 32'hc404e7b;
      36730: inst = 32'h8220000;
      36731: inst = 32'h10408000;
      36732: inst = 32'hc404e7c;
      36733: inst = 32'h8220000;
      36734: inst = 32'h10408000;
      36735: inst = 32'hc404e83;
      36736: inst = 32'h8220000;
      36737: inst = 32'h10408000;
      36738: inst = 32'hc404e84;
      36739: inst = 32'h8220000;
      36740: inst = 32'h10408000;
      36741: inst = 32'hc404e85;
      36742: inst = 32'h8220000;
      36743: inst = 32'h10408000;
      36744: inst = 32'hc404e86;
      36745: inst = 32'h8220000;
      36746: inst = 32'h10408000;
      36747: inst = 32'hc404e87;
      36748: inst = 32'h8220000;
      36749: inst = 32'h10408000;
      36750: inst = 32'hc404e88;
      36751: inst = 32'h8220000;
      36752: inst = 32'h10408000;
      36753: inst = 32'hc404e89;
      36754: inst = 32'h8220000;
      36755: inst = 32'h10408000;
      36756: inst = 32'hc404e8a;
      36757: inst = 32'h8220000;
      36758: inst = 32'h10408000;
      36759: inst = 32'hc404e8b;
      36760: inst = 32'h8220000;
      36761: inst = 32'h10408000;
      36762: inst = 32'hc404e8c;
      36763: inst = 32'h8220000;
      36764: inst = 32'h10408000;
      36765: inst = 32'hc404e8d;
      36766: inst = 32'h8220000;
      36767: inst = 32'h10408000;
      36768: inst = 32'hc404e8e;
      36769: inst = 32'h8220000;
      36770: inst = 32'h10408000;
      36771: inst = 32'hc404e8f;
      36772: inst = 32'h8220000;
      36773: inst = 32'h10408000;
      36774: inst = 32'hc404e90;
      36775: inst = 32'h8220000;
      36776: inst = 32'h10408000;
      36777: inst = 32'hc404e91;
      36778: inst = 32'h8220000;
      36779: inst = 32'h10408000;
      36780: inst = 32'hc404e92;
      36781: inst = 32'h8220000;
      36782: inst = 32'h10408000;
      36783: inst = 32'hc404e93;
      36784: inst = 32'h8220000;
      36785: inst = 32'h10408000;
      36786: inst = 32'hc404e94;
      36787: inst = 32'h8220000;
      36788: inst = 32'h10408000;
      36789: inst = 32'hc404e95;
      36790: inst = 32'h8220000;
      36791: inst = 32'h10408000;
      36792: inst = 32'hc404e96;
      36793: inst = 32'h8220000;
      36794: inst = 32'h10408000;
      36795: inst = 32'hc404e97;
      36796: inst = 32'h8220000;
      36797: inst = 32'h10408000;
      36798: inst = 32'hc404e98;
      36799: inst = 32'h8220000;
      36800: inst = 32'h10408000;
      36801: inst = 32'hc404e99;
      36802: inst = 32'h8220000;
      36803: inst = 32'h10408000;
      36804: inst = 32'hc404e9a;
      36805: inst = 32'h8220000;
      36806: inst = 32'h10408000;
      36807: inst = 32'hc404e9b;
      36808: inst = 32'h8220000;
      36809: inst = 32'h10408000;
      36810: inst = 32'hc404e9c;
      36811: inst = 32'h8220000;
      36812: inst = 32'h10408000;
      36813: inst = 32'hc404e9d;
      36814: inst = 32'h8220000;
      36815: inst = 32'h10408000;
      36816: inst = 32'hc404e9e;
      36817: inst = 32'h8220000;
      36818: inst = 32'h10408000;
      36819: inst = 32'hc404e9f;
      36820: inst = 32'h8220000;
      36821: inst = 32'h10408000;
      36822: inst = 32'hc404ea0;
      36823: inst = 32'h8220000;
      36824: inst = 32'h10408000;
      36825: inst = 32'hc404ea1;
      36826: inst = 32'h8220000;
      36827: inst = 32'h10408000;
      36828: inst = 32'hc404ea2;
      36829: inst = 32'h8220000;
      36830: inst = 32'h10408000;
      36831: inst = 32'hc404ea3;
      36832: inst = 32'h8220000;
      36833: inst = 32'h10408000;
      36834: inst = 32'hc404ea4;
      36835: inst = 32'h8220000;
      36836: inst = 32'h10408000;
      36837: inst = 32'hc404ea5;
      36838: inst = 32'h8220000;
      36839: inst = 32'h10408000;
      36840: inst = 32'hc404ea6;
      36841: inst = 32'h8220000;
      36842: inst = 32'h10408000;
      36843: inst = 32'hc404ea7;
      36844: inst = 32'h8220000;
      36845: inst = 32'h10408000;
      36846: inst = 32'hc404ea8;
      36847: inst = 32'h8220000;
      36848: inst = 32'h10408000;
      36849: inst = 32'hc404ea9;
      36850: inst = 32'h8220000;
      36851: inst = 32'h10408000;
      36852: inst = 32'hc404eaa;
      36853: inst = 32'h8220000;
      36854: inst = 32'h10408000;
      36855: inst = 32'hc404eab;
      36856: inst = 32'h8220000;
      36857: inst = 32'h10408000;
      36858: inst = 32'hc404eac;
      36859: inst = 32'h8220000;
      36860: inst = 32'h10408000;
      36861: inst = 32'hc404ead;
      36862: inst = 32'h8220000;
      36863: inst = 32'h10408000;
      36864: inst = 32'hc404eae;
      36865: inst = 32'h8220000;
      36866: inst = 32'h10408000;
      36867: inst = 32'hc404eaf;
      36868: inst = 32'h8220000;
      36869: inst = 32'h10408000;
      36870: inst = 32'hc404eb0;
      36871: inst = 32'h8220000;
      36872: inst = 32'h10408000;
      36873: inst = 32'hc404eb1;
      36874: inst = 32'h8220000;
      36875: inst = 32'h10408000;
      36876: inst = 32'hc404eb2;
      36877: inst = 32'h8220000;
      36878: inst = 32'h10408000;
      36879: inst = 32'hc404eb3;
      36880: inst = 32'h8220000;
      36881: inst = 32'h10408000;
      36882: inst = 32'hc404eb4;
      36883: inst = 32'h8220000;
      36884: inst = 32'h10408000;
      36885: inst = 32'hc404eb5;
      36886: inst = 32'h8220000;
      36887: inst = 32'h10408000;
      36888: inst = 32'hc404eb6;
      36889: inst = 32'h8220000;
      36890: inst = 32'h10408000;
      36891: inst = 32'hc404eb7;
      36892: inst = 32'h8220000;
      36893: inst = 32'h10408000;
      36894: inst = 32'hc404ebb;
      36895: inst = 32'h8220000;
      36896: inst = 32'h10408000;
      36897: inst = 32'hc404ebc;
      36898: inst = 32'h8220000;
      36899: inst = 32'h10408000;
      36900: inst = 32'hc404ebd;
      36901: inst = 32'h8220000;
      36902: inst = 32'h10408000;
      36903: inst = 32'hc404ebe;
      36904: inst = 32'h8220000;
      36905: inst = 32'h10408000;
      36906: inst = 32'hc404ebf;
      36907: inst = 32'h8220000;
      36908: inst = 32'h10408000;
      36909: inst = 32'hc404ec0;
      36910: inst = 32'h8220000;
      36911: inst = 32'h10408000;
      36912: inst = 32'hc404ec1;
      36913: inst = 32'h8220000;
      36914: inst = 32'h10408000;
      36915: inst = 32'hc404ec2;
      36916: inst = 32'h8220000;
      36917: inst = 32'h10408000;
      36918: inst = 32'hc404ec3;
      36919: inst = 32'h8220000;
      36920: inst = 32'h10408000;
      36921: inst = 32'hc404ec4;
      36922: inst = 32'h8220000;
      36923: inst = 32'h10408000;
      36924: inst = 32'hc404ec5;
      36925: inst = 32'h8220000;
      36926: inst = 32'h10408000;
      36927: inst = 32'hc404ec6;
      36928: inst = 32'h8220000;
      36929: inst = 32'h10408000;
      36930: inst = 32'hc404ec7;
      36931: inst = 32'h8220000;
      36932: inst = 32'h10408000;
      36933: inst = 32'hc404ec8;
      36934: inst = 32'h8220000;
      36935: inst = 32'h10408000;
      36936: inst = 32'hc404ec9;
      36937: inst = 32'h8220000;
      36938: inst = 32'h10408000;
      36939: inst = 32'hc404eca;
      36940: inst = 32'h8220000;
      36941: inst = 32'h10408000;
      36942: inst = 32'hc404ecb;
      36943: inst = 32'h8220000;
      36944: inst = 32'h10408000;
      36945: inst = 32'hc404ecc;
      36946: inst = 32'h8220000;
      36947: inst = 32'h10408000;
      36948: inst = 32'hc404ecd;
      36949: inst = 32'h8220000;
      36950: inst = 32'h10408000;
      36951: inst = 32'hc404ece;
      36952: inst = 32'h8220000;
      36953: inst = 32'h10408000;
      36954: inst = 32'hc404ecf;
      36955: inst = 32'h8220000;
      36956: inst = 32'h10408000;
      36957: inst = 32'hc404ed0;
      36958: inst = 32'h8220000;
      36959: inst = 32'h10408000;
      36960: inst = 32'hc404ed1;
      36961: inst = 32'h8220000;
      36962: inst = 32'h10408000;
      36963: inst = 32'hc404ed2;
      36964: inst = 32'h8220000;
      36965: inst = 32'h10408000;
      36966: inst = 32'hc404ed3;
      36967: inst = 32'h8220000;
      36968: inst = 32'h10408000;
      36969: inst = 32'hc404ed4;
      36970: inst = 32'h8220000;
      36971: inst = 32'h10408000;
      36972: inst = 32'hc404ed5;
      36973: inst = 32'h8220000;
      36974: inst = 32'h10408000;
      36975: inst = 32'hc404ed6;
      36976: inst = 32'h8220000;
      36977: inst = 32'h10408000;
      36978: inst = 32'hc404ed7;
      36979: inst = 32'h8220000;
      36980: inst = 32'h10408000;
      36981: inst = 32'hc404ed8;
      36982: inst = 32'h8220000;
      36983: inst = 32'h10408000;
      36984: inst = 32'hc404ed9;
      36985: inst = 32'h8220000;
      36986: inst = 32'h10408000;
      36987: inst = 32'hc404eda;
      36988: inst = 32'h8220000;
      36989: inst = 32'h10408000;
      36990: inst = 32'hc404edb;
      36991: inst = 32'h8220000;
      36992: inst = 32'h10408000;
      36993: inst = 32'hc404edc;
      36994: inst = 32'h8220000;
      36995: inst = 32'h10408000;
      36996: inst = 32'hc404ee3;
      36997: inst = 32'h8220000;
      36998: inst = 32'h10408000;
      36999: inst = 32'hc404ee4;
      37000: inst = 32'h8220000;
      37001: inst = 32'h10408000;
      37002: inst = 32'hc404ee5;
      37003: inst = 32'h8220000;
      37004: inst = 32'h10408000;
      37005: inst = 32'hc404ee6;
      37006: inst = 32'h8220000;
      37007: inst = 32'h10408000;
      37008: inst = 32'hc404ee7;
      37009: inst = 32'h8220000;
      37010: inst = 32'h10408000;
      37011: inst = 32'hc404ee8;
      37012: inst = 32'h8220000;
      37013: inst = 32'h10408000;
      37014: inst = 32'hc404ee9;
      37015: inst = 32'h8220000;
      37016: inst = 32'h10408000;
      37017: inst = 32'hc404eea;
      37018: inst = 32'h8220000;
      37019: inst = 32'h10408000;
      37020: inst = 32'hc404eeb;
      37021: inst = 32'h8220000;
      37022: inst = 32'h10408000;
      37023: inst = 32'hc404eec;
      37024: inst = 32'h8220000;
      37025: inst = 32'h10408000;
      37026: inst = 32'hc404eed;
      37027: inst = 32'h8220000;
      37028: inst = 32'h10408000;
      37029: inst = 32'hc404eee;
      37030: inst = 32'h8220000;
      37031: inst = 32'h10408000;
      37032: inst = 32'hc404eef;
      37033: inst = 32'h8220000;
      37034: inst = 32'h10408000;
      37035: inst = 32'hc404ef0;
      37036: inst = 32'h8220000;
      37037: inst = 32'h10408000;
      37038: inst = 32'hc404ef1;
      37039: inst = 32'h8220000;
      37040: inst = 32'h10408000;
      37041: inst = 32'hc404ef2;
      37042: inst = 32'h8220000;
      37043: inst = 32'h10408000;
      37044: inst = 32'hc404ef3;
      37045: inst = 32'h8220000;
      37046: inst = 32'h10408000;
      37047: inst = 32'hc404ef4;
      37048: inst = 32'h8220000;
      37049: inst = 32'h10408000;
      37050: inst = 32'hc404ef5;
      37051: inst = 32'h8220000;
      37052: inst = 32'h10408000;
      37053: inst = 32'hc404ef6;
      37054: inst = 32'h8220000;
      37055: inst = 32'h10408000;
      37056: inst = 32'hc404ef7;
      37057: inst = 32'h8220000;
      37058: inst = 32'h10408000;
      37059: inst = 32'hc404ef8;
      37060: inst = 32'h8220000;
      37061: inst = 32'h10408000;
      37062: inst = 32'hc404ef9;
      37063: inst = 32'h8220000;
      37064: inst = 32'h10408000;
      37065: inst = 32'hc404efa;
      37066: inst = 32'h8220000;
      37067: inst = 32'h10408000;
      37068: inst = 32'hc404efb;
      37069: inst = 32'h8220000;
      37070: inst = 32'h10408000;
      37071: inst = 32'hc404efc;
      37072: inst = 32'h8220000;
      37073: inst = 32'h10408000;
      37074: inst = 32'hc404efd;
      37075: inst = 32'h8220000;
      37076: inst = 32'h10408000;
      37077: inst = 32'hc404efe;
      37078: inst = 32'h8220000;
      37079: inst = 32'h10408000;
      37080: inst = 32'hc404eff;
      37081: inst = 32'h8220000;
      37082: inst = 32'h10408000;
      37083: inst = 32'hc404f00;
      37084: inst = 32'h8220000;
      37085: inst = 32'h10408000;
      37086: inst = 32'hc404f01;
      37087: inst = 32'h8220000;
      37088: inst = 32'h10408000;
      37089: inst = 32'hc404f02;
      37090: inst = 32'h8220000;
      37091: inst = 32'h10408000;
      37092: inst = 32'hc404f03;
      37093: inst = 32'h8220000;
      37094: inst = 32'h10408000;
      37095: inst = 32'hc404f04;
      37096: inst = 32'h8220000;
      37097: inst = 32'h10408000;
      37098: inst = 32'hc404f05;
      37099: inst = 32'h8220000;
      37100: inst = 32'h10408000;
      37101: inst = 32'hc404f06;
      37102: inst = 32'h8220000;
      37103: inst = 32'h10408000;
      37104: inst = 32'hc404f07;
      37105: inst = 32'h8220000;
      37106: inst = 32'h10408000;
      37107: inst = 32'hc404f08;
      37108: inst = 32'h8220000;
      37109: inst = 32'h10408000;
      37110: inst = 32'hc404f09;
      37111: inst = 32'h8220000;
      37112: inst = 32'h10408000;
      37113: inst = 32'hc404f0a;
      37114: inst = 32'h8220000;
      37115: inst = 32'h10408000;
      37116: inst = 32'hc404f0b;
      37117: inst = 32'h8220000;
      37118: inst = 32'h10408000;
      37119: inst = 32'hc404f0c;
      37120: inst = 32'h8220000;
      37121: inst = 32'h10408000;
      37122: inst = 32'hc404f0d;
      37123: inst = 32'h8220000;
      37124: inst = 32'h10408000;
      37125: inst = 32'hc404f0e;
      37126: inst = 32'h8220000;
      37127: inst = 32'h10408000;
      37128: inst = 32'hc404f0f;
      37129: inst = 32'h8220000;
      37130: inst = 32'h10408000;
      37131: inst = 32'hc404f10;
      37132: inst = 32'h8220000;
      37133: inst = 32'h10408000;
      37134: inst = 32'hc404f11;
      37135: inst = 32'h8220000;
      37136: inst = 32'h10408000;
      37137: inst = 32'hc404f12;
      37138: inst = 32'h8220000;
      37139: inst = 32'h10408000;
      37140: inst = 32'hc404f13;
      37141: inst = 32'h8220000;
      37142: inst = 32'h10408000;
      37143: inst = 32'hc404f14;
      37144: inst = 32'h8220000;
      37145: inst = 32'h10408000;
      37146: inst = 32'hc404f15;
      37147: inst = 32'h8220000;
      37148: inst = 32'h10408000;
      37149: inst = 32'hc404f16;
      37150: inst = 32'h8220000;
      37151: inst = 32'h10408000;
      37152: inst = 32'hc404f17;
      37153: inst = 32'h8220000;
      37154: inst = 32'h10408000;
      37155: inst = 32'hc404f1b;
      37156: inst = 32'h8220000;
      37157: inst = 32'h10408000;
      37158: inst = 32'hc404f1c;
      37159: inst = 32'h8220000;
      37160: inst = 32'h10408000;
      37161: inst = 32'hc404f1d;
      37162: inst = 32'h8220000;
      37163: inst = 32'h10408000;
      37164: inst = 32'hc404f1e;
      37165: inst = 32'h8220000;
      37166: inst = 32'h10408000;
      37167: inst = 32'hc404f1f;
      37168: inst = 32'h8220000;
      37169: inst = 32'h10408000;
      37170: inst = 32'hc404f20;
      37171: inst = 32'h8220000;
      37172: inst = 32'h10408000;
      37173: inst = 32'hc404f21;
      37174: inst = 32'h8220000;
      37175: inst = 32'h10408000;
      37176: inst = 32'hc404f22;
      37177: inst = 32'h8220000;
      37178: inst = 32'h10408000;
      37179: inst = 32'hc404f23;
      37180: inst = 32'h8220000;
      37181: inst = 32'h10408000;
      37182: inst = 32'hc404f24;
      37183: inst = 32'h8220000;
      37184: inst = 32'h10408000;
      37185: inst = 32'hc404f25;
      37186: inst = 32'h8220000;
      37187: inst = 32'h10408000;
      37188: inst = 32'hc404f26;
      37189: inst = 32'h8220000;
      37190: inst = 32'h10408000;
      37191: inst = 32'hc404f27;
      37192: inst = 32'h8220000;
      37193: inst = 32'h10408000;
      37194: inst = 32'hc404f28;
      37195: inst = 32'h8220000;
      37196: inst = 32'h10408000;
      37197: inst = 32'hc404f29;
      37198: inst = 32'h8220000;
      37199: inst = 32'h10408000;
      37200: inst = 32'hc404f2a;
      37201: inst = 32'h8220000;
      37202: inst = 32'h10408000;
      37203: inst = 32'hc404f2b;
      37204: inst = 32'h8220000;
      37205: inst = 32'h10408000;
      37206: inst = 32'hc404f2c;
      37207: inst = 32'h8220000;
      37208: inst = 32'h10408000;
      37209: inst = 32'hc404f2d;
      37210: inst = 32'h8220000;
      37211: inst = 32'h10408000;
      37212: inst = 32'hc404f2e;
      37213: inst = 32'h8220000;
      37214: inst = 32'h10408000;
      37215: inst = 32'hc404f2f;
      37216: inst = 32'h8220000;
      37217: inst = 32'h10408000;
      37218: inst = 32'hc404f30;
      37219: inst = 32'h8220000;
      37220: inst = 32'h10408000;
      37221: inst = 32'hc404f31;
      37222: inst = 32'h8220000;
      37223: inst = 32'h10408000;
      37224: inst = 32'hc404f32;
      37225: inst = 32'h8220000;
      37226: inst = 32'h10408000;
      37227: inst = 32'hc404f33;
      37228: inst = 32'h8220000;
      37229: inst = 32'h10408000;
      37230: inst = 32'hc404f34;
      37231: inst = 32'h8220000;
      37232: inst = 32'h10408000;
      37233: inst = 32'hc404f35;
      37234: inst = 32'h8220000;
      37235: inst = 32'h10408000;
      37236: inst = 32'hc404f36;
      37237: inst = 32'h8220000;
      37238: inst = 32'h10408000;
      37239: inst = 32'hc404f37;
      37240: inst = 32'h8220000;
      37241: inst = 32'h10408000;
      37242: inst = 32'hc404f38;
      37243: inst = 32'h8220000;
      37244: inst = 32'h10408000;
      37245: inst = 32'hc404f39;
      37246: inst = 32'h8220000;
      37247: inst = 32'h10408000;
      37248: inst = 32'hc404f3a;
      37249: inst = 32'h8220000;
      37250: inst = 32'h10408000;
      37251: inst = 32'hc404f3b;
      37252: inst = 32'h8220000;
      37253: inst = 32'h10408000;
      37254: inst = 32'hc404f3c;
      37255: inst = 32'h8220000;
      37256: inst = 32'h10408000;
      37257: inst = 32'hc404f43;
      37258: inst = 32'h8220000;
      37259: inst = 32'h10408000;
      37260: inst = 32'hc404f44;
      37261: inst = 32'h8220000;
      37262: inst = 32'h10408000;
      37263: inst = 32'hc404f45;
      37264: inst = 32'h8220000;
      37265: inst = 32'h10408000;
      37266: inst = 32'hc404f46;
      37267: inst = 32'h8220000;
      37268: inst = 32'h10408000;
      37269: inst = 32'hc404f47;
      37270: inst = 32'h8220000;
      37271: inst = 32'h10408000;
      37272: inst = 32'hc404f48;
      37273: inst = 32'h8220000;
      37274: inst = 32'h10408000;
      37275: inst = 32'hc404f49;
      37276: inst = 32'h8220000;
      37277: inst = 32'h10408000;
      37278: inst = 32'hc404f4a;
      37279: inst = 32'h8220000;
      37280: inst = 32'h10408000;
      37281: inst = 32'hc404f4b;
      37282: inst = 32'h8220000;
      37283: inst = 32'h10408000;
      37284: inst = 32'hc404f4c;
      37285: inst = 32'h8220000;
      37286: inst = 32'h10408000;
      37287: inst = 32'hc404f4d;
      37288: inst = 32'h8220000;
      37289: inst = 32'h10408000;
      37290: inst = 32'hc404f4e;
      37291: inst = 32'h8220000;
      37292: inst = 32'h10408000;
      37293: inst = 32'hc404f4f;
      37294: inst = 32'h8220000;
      37295: inst = 32'h10408000;
      37296: inst = 32'hc404f50;
      37297: inst = 32'h8220000;
      37298: inst = 32'h10408000;
      37299: inst = 32'hc404f51;
      37300: inst = 32'h8220000;
      37301: inst = 32'h10408000;
      37302: inst = 32'hc404f52;
      37303: inst = 32'h8220000;
      37304: inst = 32'h10408000;
      37305: inst = 32'hc404f53;
      37306: inst = 32'h8220000;
      37307: inst = 32'h10408000;
      37308: inst = 32'hc404f54;
      37309: inst = 32'h8220000;
      37310: inst = 32'h10408000;
      37311: inst = 32'hc404f55;
      37312: inst = 32'h8220000;
      37313: inst = 32'h10408000;
      37314: inst = 32'hc404f56;
      37315: inst = 32'h8220000;
      37316: inst = 32'h10408000;
      37317: inst = 32'hc404f57;
      37318: inst = 32'h8220000;
      37319: inst = 32'h10408000;
      37320: inst = 32'hc404f58;
      37321: inst = 32'h8220000;
      37322: inst = 32'h10408000;
      37323: inst = 32'hc404f59;
      37324: inst = 32'h8220000;
      37325: inst = 32'h10408000;
      37326: inst = 32'hc404f5a;
      37327: inst = 32'h8220000;
      37328: inst = 32'h10408000;
      37329: inst = 32'hc404f5b;
      37330: inst = 32'h8220000;
      37331: inst = 32'h10408000;
      37332: inst = 32'hc404f5c;
      37333: inst = 32'h8220000;
      37334: inst = 32'h10408000;
      37335: inst = 32'hc404f5d;
      37336: inst = 32'h8220000;
      37337: inst = 32'h10408000;
      37338: inst = 32'hc404f5e;
      37339: inst = 32'h8220000;
      37340: inst = 32'h10408000;
      37341: inst = 32'hc404f5f;
      37342: inst = 32'h8220000;
      37343: inst = 32'h10408000;
      37344: inst = 32'hc404f60;
      37345: inst = 32'h8220000;
      37346: inst = 32'h10408000;
      37347: inst = 32'hc404f61;
      37348: inst = 32'h8220000;
      37349: inst = 32'h10408000;
      37350: inst = 32'hc404f62;
      37351: inst = 32'h8220000;
      37352: inst = 32'h10408000;
      37353: inst = 32'hc404f63;
      37354: inst = 32'h8220000;
      37355: inst = 32'h10408000;
      37356: inst = 32'hc404f64;
      37357: inst = 32'h8220000;
      37358: inst = 32'h10408000;
      37359: inst = 32'hc404f65;
      37360: inst = 32'h8220000;
      37361: inst = 32'h10408000;
      37362: inst = 32'hc404f66;
      37363: inst = 32'h8220000;
      37364: inst = 32'h10408000;
      37365: inst = 32'hc404f67;
      37366: inst = 32'h8220000;
      37367: inst = 32'h10408000;
      37368: inst = 32'hc404f68;
      37369: inst = 32'h8220000;
      37370: inst = 32'h10408000;
      37371: inst = 32'hc404f69;
      37372: inst = 32'h8220000;
      37373: inst = 32'h10408000;
      37374: inst = 32'hc404f6a;
      37375: inst = 32'h8220000;
      37376: inst = 32'h10408000;
      37377: inst = 32'hc404f6b;
      37378: inst = 32'h8220000;
      37379: inst = 32'h10408000;
      37380: inst = 32'hc404f6c;
      37381: inst = 32'h8220000;
      37382: inst = 32'h10408000;
      37383: inst = 32'hc404f6d;
      37384: inst = 32'h8220000;
      37385: inst = 32'h10408000;
      37386: inst = 32'hc404f6e;
      37387: inst = 32'h8220000;
      37388: inst = 32'h10408000;
      37389: inst = 32'hc404f6f;
      37390: inst = 32'h8220000;
      37391: inst = 32'h10408000;
      37392: inst = 32'hc404f70;
      37393: inst = 32'h8220000;
      37394: inst = 32'h10408000;
      37395: inst = 32'hc404f71;
      37396: inst = 32'h8220000;
      37397: inst = 32'h10408000;
      37398: inst = 32'hc404f72;
      37399: inst = 32'h8220000;
      37400: inst = 32'h10408000;
      37401: inst = 32'hc404f73;
      37402: inst = 32'h8220000;
      37403: inst = 32'h10408000;
      37404: inst = 32'hc404f74;
      37405: inst = 32'h8220000;
      37406: inst = 32'h10408000;
      37407: inst = 32'hc404f75;
      37408: inst = 32'h8220000;
      37409: inst = 32'h10408000;
      37410: inst = 32'hc404f76;
      37411: inst = 32'h8220000;
      37412: inst = 32'h10408000;
      37413: inst = 32'hc404f77;
      37414: inst = 32'h8220000;
      37415: inst = 32'h10408000;
      37416: inst = 32'hc404f7b;
      37417: inst = 32'h8220000;
      37418: inst = 32'h10408000;
      37419: inst = 32'hc404f7c;
      37420: inst = 32'h8220000;
      37421: inst = 32'h10408000;
      37422: inst = 32'hc404f7d;
      37423: inst = 32'h8220000;
      37424: inst = 32'h10408000;
      37425: inst = 32'hc404f7e;
      37426: inst = 32'h8220000;
      37427: inst = 32'h10408000;
      37428: inst = 32'hc404f7f;
      37429: inst = 32'h8220000;
      37430: inst = 32'h10408000;
      37431: inst = 32'hc404f80;
      37432: inst = 32'h8220000;
      37433: inst = 32'h10408000;
      37434: inst = 32'hc404f81;
      37435: inst = 32'h8220000;
      37436: inst = 32'h10408000;
      37437: inst = 32'hc404f82;
      37438: inst = 32'h8220000;
      37439: inst = 32'h10408000;
      37440: inst = 32'hc404f83;
      37441: inst = 32'h8220000;
      37442: inst = 32'h10408000;
      37443: inst = 32'hc404f84;
      37444: inst = 32'h8220000;
      37445: inst = 32'h10408000;
      37446: inst = 32'hc404f85;
      37447: inst = 32'h8220000;
      37448: inst = 32'h10408000;
      37449: inst = 32'hc404f86;
      37450: inst = 32'h8220000;
      37451: inst = 32'h10408000;
      37452: inst = 32'hc404f87;
      37453: inst = 32'h8220000;
      37454: inst = 32'h10408000;
      37455: inst = 32'hc404f88;
      37456: inst = 32'h8220000;
      37457: inst = 32'h10408000;
      37458: inst = 32'hc404f89;
      37459: inst = 32'h8220000;
      37460: inst = 32'h10408000;
      37461: inst = 32'hc404f8a;
      37462: inst = 32'h8220000;
      37463: inst = 32'h10408000;
      37464: inst = 32'hc404f8b;
      37465: inst = 32'h8220000;
      37466: inst = 32'h10408000;
      37467: inst = 32'hc404f8c;
      37468: inst = 32'h8220000;
      37469: inst = 32'h10408000;
      37470: inst = 32'hc404f8d;
      37471: inst = 32'h8220000;
      37472: inst = 32'h10408000;
      37473: inst = 32'hc404f8e;
      37474: inst = 32'h8220000;
      37475: inst = 32'h10408000;
      37476: inst = 32'hc404f8f;
      37477: inst = 32'h8220000;
      37478: inst = 32'h10408000;
      37479: inst = 32'hc404f90;
      37480: inst = 32'h8220000;
      37481: inst = 32'h10408000;
      37482: inst = 32'hc404f91;
      37483: inst = 32'h8220000;
      37484: inst = 32'h10408000;
      37485: inst = 32'hc404f92;
      37486: inst = 32'h8220000;
      37487: inst = 32'h10408000;
      37488: inst = 32'hc404f93;
      37489: inst = 32'h8220000;
      37490: inst = 32'h10408000;
      37491: inst = 32'hc404f94;
      37492: inst = 32'h8220000;
      37493: inst = 32'h10408000;
      37494: inst = 32'hc404f95;
      37495: inst = 32'h8220000;
      37496: inst = 32'h10408000;
      37497: inst = 32'hc404f96;
      37498: inst = 32'h8220000;
      37499: inst = 32'h10408000;
      37500: inst = 32'hc404f97;
      37501: inst = 32'h8220000;
      37502: inst = 32'h10408000;
      37503: inst = 32'hc404f98;
      37504: inst = 32'h8220000;
      37505: inst = 32'h10408000;
      37506: inst = 32'hc404f99;
      37507: inst = 32'h8220000;
      37508: inst = 32'h10408000;
      37509: inst = 32'hc404f9a;
      37510: inst = 32'h8220000;
      37511: inst = 32'h10408000;
      37512: inst = 32'hc404f9b;
      37513: inst = 32'h8220000;
      37514: inst = 32'h10408000;
      37515: inst = 32'hc404f9c;
      37516: inst = 32'h8220000;
      37517: inst = 32'h10408000;
      37518: inst = 32'hc404fa3;
      37519: inst = 32'h8220000;
      37520: inst = 32'h10408000;
      37521: inst = 32'hc404fa4;
      37522: inst = 32'h8220000;
      37523: inst = 32'h10408000;
      37524: inst = 32'hc404fa5;
      37525: inst = 32'h8220000;
      37526: inst = 32'h10408000;
      37527: inst = 32'hc404fa6;
      37528: inst = 32'h8220000;
      37529: inst = 32'h10408000;
      37530: inst = 32'hc404fa7;
      37531: inst = 32'h8220000;
      37532: inst = 32'h10408000;
      37533: inst = 32'hc404fa8;
      37534: inst = 32'h8220000;
      37535: inst = 32'h10408000;
      37536: inst = 32'hc404fa9;
      37537: inst = 32'h8220000;
      37538: inst = 32'h10408000;
      37539: inst = 32'hc404faa;
      37540: inst = 32'h8220000;
      37541: inst = 32'h10408000;
      37542: inst = 32'hc404fab;
      37543: inst = 32'h8220000;
      37544: inst = 32'h10408000;
      37545: inst = 32'hc404fac;
      37546: inst = 32'h8220000;
      37547: inst = 32'h10408000;
      37548: inst = 32'hc404fad;
      37549: inst = 32'h8220000;
      37550: inst = 32'h10408000;
      37551: inst = 32'hc404fae;
      37552: inst = 32'h8220000;
      37553: inst = 32'h10408000;
      37554: inst = 32'hc404faf;
      37555: inst = 32'h8220000;
      37556: inst = 32'h10408000;
      37557: inst = 32'hc404fb0;
      37558: inst = 32'h8220000;
      37559: inst = 32'h10408000;
      37560: inst = 32'hc404fb1;
      37561: inst = 32'h8220000;
      37562: inst = 32'h10408000;
      37563: inst = 32'hc404fb2;
      37564: inst = 32'h8220000;
      37565: inst = 32'h10408000;
      37566: inst = 32'hc404fb3;
      37567: inst = 32'h8220000;
      37568: inst = 32'h10408000;
      37569: inst = 32'hc404fb4;
      37570: inst = 32'h8220000;
      37571: inst = 32'h10408000;
      37572: inst = 32'hc404fb5;
      37573: inst = 32'h8220000;
      37574: inst = 32'h10408000;
      37575: inst = 32'hc404fb6;
      37576: inst = 32'h8220000;
      37577: inst = 32'h10408000;
      37578: inst = 32'hc404fb7;
      37579: inst = 32'h8220000;
      37580: inst = 32'h10408000;
      37581: inst = 32'hc404fb8;
      37582: inst = 32'h8220000;
      37583: inst = 32'h10408000;
      37584: inst = 32'hc404fb9;
      37585: inst = 32'h8220000;
      37586: inst = 32'h10408000;
      37587: inst = 32'hc404fba;
      37588: inst = 32'h8220000;
      37589: inst = 32'h10408000;
      37590: inst = 32'hc404fbb;
      37591: inst = 32'h8220000;
      37592: inst = 32'h10408000;
      37593: inst = 32'hc404fbc;
      37594: inst = 32'h8220000;
      37595: inst = 32'h10408000;
      37596: inst = 32'hc404fbd;
      37597: inst = 32'h8220000;
      37598: inst = 32'h10408000;
      37599: inst = 32'hc404fbe;
      37600: inst = 32'h8220000;
      37601: inst = 32'h10408000;
      37602: inst = 32'hc404fbf;
      37603: inst = 32'h8220000;
      37604: inst = 32'h10408000;
      37605: inst = 32'hc404fc0;
      37606: inst = 32'h8220000;
      37607: inst = 32'h10408000;
      37608: inst = 32'hc404fc1;
      37609: inst = 32'h8220000;
      37610: inst = 32'h10408000;
      37611: inst = 32'hc404fc2;
      37612: inst = 32'h8220000;
      37613: inst = 32'h10408000;
      37614: inst = 32'hc404fc3;
      37615: inst = 32'h8220000;
      37616: inst = 32'h10408000;
      37617: inst = 32'hc404fc4;
      37618: inst = 32'h8220000;
      37619: inst = 32'h10408000;
      37620: inst = 32'hc404fc5;
      37621: inst = 32'h8220000;
      37622: inst = 32'h10408000;
      37623: inst = 32'hc404fc6;
      37624: inst = 32'h8220000;
      37625: inst = 32'h10408000;
      37626: inst = 32'hc404fc7;
      37627: inst = 32'h8220000;
      37628: inst = 32'h10408000;
      37629: inst = 32'hc404fc8;
      37630: inst = 32'h8220000;
      37631: inst = 32'h10408000;
      37632: inst = 32'hc404fc9;
      37633: inst = 32'h8220000;
      37634: inst = 32'h10408000;
      37635: inst = 32'hc404fca;
      37636: inst = 32'h8220000;
      37637: inst = 32'h10408000;
      37638: inst = 32'hc404fcb;
      37639: inst = 32'h8220000;
      37640: inst = 32'h10408000;
      37641: inst = 32'hc404fcc;
      37642: inst = 32'h8220000;
      37643: inst = 32'h10408000;
      37644: inst = 32'hc404fcd;
      37645: inst = 32'h8220000;
      37646: inst = 32'h10408000;
      37647: inst = 32'hc404fce;
      37648: inst = 32'h8220000;
      37649: inst = 32'h10408000;
      37650: inst = 32'hc404fcf;
      37651: inst = 32'h8220000;
      37652: inst = 32'h10408000;
      37653: inst = 32'hc404fd0;
      37654: inst = 32'h8220000;
      37655: inst = 32'h10408000;
      37656: inst = 32'hc404fd1;
      37657: inst = 32'h8220000;
      37658: inst = 32'h10408000;
      37659: inst = 32'hc404fd2;
      37660: inst = 32'h8220000;
      37661: inst = 32'h10408000;
      37662: inst = 32'hc404fd3;
      37663: inst = 32'h8220000;
      37664: inst = 32'h10408000;
      37665: inst = 32'hc404fd4;
      37666: inst = 32'h8220000;
      37667: inst = 32'h10408000;
      37668: inst = 32'hc404fd5;
      37669: inst = 32'h8220000;
      37670: inst = 32'h10408000;
      37671: inst = 32'hc404fd6;
      37672: inst = 32'h8220000;
      37673: inst = 32'h10408000;
      37674: inst = 32'hc404fd7;
      37675: inst = 32'h8220000;
      37676: inst = 32'h10408000;
      37677: inst = 32'hc404fdb;
      37678: inst = 32'h8220000;
      37679: inst = 32'h10408000;
      37680: inst = 32'hc404fdc;
      37681: inst = 32'h8220000;
      37682: inst = 32'h10408000;
      37683: inst = 32'hc404fdd;
      37684: inst = 32'h8220000;
      37685: inst = 32'h10408000;
      37686: inst = 32'hc404fde;
      37687: inst = 32'h8220000;
      37688: inst = 32'h10408000;
      37689: inst = 32'hc404fdf;
      37690: inst = 32'h8220000;
      37691: inst = 32'h10408000;
      37692: inst = 32'hc404fe0;
      37693: inst = 32'h8220000;
      37694: inst = 32'h10408000;
      37695: inst = 32'hc404fe1;
      37696: inst = 32'h8220000;
      37697: inst = 32'h10408000;
      37698: inst = 32'hc404fe2;
      37699: inst = 32'h8220000;
      37700: inst = 32'h10408000;
      37701: inst = 32'hc404fe3;
      37702: inst = 32'h8220000;
      37703: inst = 32'h10408000;
      37704: inst = 32'hc404fe4;
      37705: inst = 32'h8220000;
      37706: inst = 32'h10408000;
      37707: inst = 32'hc404fe5;
      37708: inst = 32'h8220000;
      37709: inst = 32'h10408000;
      37710: inst = 32'hc404fe6;
      37711: inst = 32'h8220000;
      37712: inst = 32'h10408000;
      37713: inst = 32'hc404fe7;
      37714: inst = 32'h8220000;
      37715: inst = 32'h10408000;
      37716: inst = 32'hc404fe8;
      37717: inst = 32'h8220000;
      37718: inst = 32'h10408000;
      37719: inst = 32'hc404fe9;
      37720: inst = 32'h8220000;
      37721: inst = 32'h10408000;
      37722: inst = 32'hc404fea;
      37723: inst = 32'h8220000;
      37724: inst = 32'h10408000;
      37725: inst = 32'hc404feb;
      37726: inst = 32'h8220000;
      37727: inst = 32'h10408000;
      37728: inst = 32'hc404fec;
      37729: inst = 32'h8220000;
      37730: inst = 32'h10408000;
      37731: inst = 32'hc404fed;
      37732: inst = 32'h8220000;
      37733: inst = 32'h10408000;
      37734: inst = 32'hc404fee;
      37735: inst = 32'h8220000;
      37736: inst = 32'h10408000;
      37737: inst = 32'hc404fef;
      37738: inst = 32'h8220000;
      37739: inst = 32'h10408000;
      37740: inst = 32'hc404ff0;
      37741: inst = 32'h8220000;
      37742: inst = 32'h10408000;
      37743: inst = 32'hc404ff1;
      37744: inst = 32'h8220000;
      37745: inst = 32'h10408000;
      37746: inst = 32'hc404ff2;
      37747: inst = 32'h8220000;
      37748: inst = 32'h10408000;
      37749: inst = 32'hc404ff3;
      37750: inst = 32'h8220000;
      37751: inst = 32'h10408000;
      37752: inst = 32'hc404ff4;
      37753: inst = 32'h8220000;
      37754: inst = 32'h10408000;
      37755: inst = 32'hc404ff5;
      37756: inst = 32'h8220000;
      37757: inst = 32'h10408000;
      37758: inst = 32'hc404ff6;
      37759: inst = 32'h8220000;
      37760: inst = 32'h10408000;
      37761: inst = 32'hc404ff7;
      37762: inst = 32'h8220000;
      37763: inst = 32'h10408000;
      37764: inst = 32'hc404ff8;
      37765: inst = 32'h8220000;
      37766: inst = 32'h10408000;
      37767: inst = 32'hc404ff9;
      37768: inst = 32'h8220000;
      37769: inst = 32'h10408000;
      37770: inst = 32'hc404ffa;
      37771: inst = 32'h8220000;
      37772: inst = 32'h10408000;
      37773: inst = 32'hc404ffb;
      37774: inst = 32'h8220000;
      37775: inst = 32'h10408000;
      37776: inst = 32'hc404ffc;
      37777: inst = 32'h8220000;
      37778: inst = 32'h10408000;
      37779: inst = 32'hc405003;
      37780: inst = 32'h8220000;
      37781: inst = 32'h10408000;
      37782: inst = 32'hc405004;
      37783: inst = 32'h8220000;
      37784: inst = 32'h10408000;
      37785: inst = 32'hc405005;
      37786: inst = 32'h8220000;
      37787: inst = 32'h10408000;
      37788: inst = 32'hc405006;
      37789: inst = 32'h8220000;
      37790: inst = 32'h10408000;
      37791: inst = 32'hc405007;
      37792: inst = 32'h8220000;
      37793: inst = 32'h10408000;
      37794: inst = 32'hc405008;
      37795: inst = 32'h8220000;
      37796: inst = 32'h10408000;
      37797: inst = 32'hc405009;
      37798: inst = 32'h8220000;
      37799: inst = 32'h10408000;
      37800: inst = 32'hc40500a;
      37801: inst = 32'h8220000;
      37802: inst = 32'h10408000;
      37803: inst = 32'hc40500b;
      37804: inst = 32'h8220000;
      37805: inst = 32'h10408000;
      37806: inst = 32'hc40500c;
      37807: inst = 32'h8220000;
      37808: inst = 32'h10408000;
      37809: inst = 32'hc40500d;
      37810: inst = 32'h8220000;
      37811: inst = 32'h10408000;
      37812: inst = 32'hc40500e;
      37813: inst = 32'h8220000;
      37814: inst = 32'h10408000;
      37815: inst = 32'hc40500f;
      37816: inst = 32'h8220000;
      37817: inst = 32'h10408000;
      37818: inst = 32'hc405010;
      37819: inst = 32'h8220000;
      37820: inst = 32'h10408000;
      37821: inst = 32'hc405011;
      37822: inst = 32'h8220000;
      37823: inst = 32'h10408000;
      37824: inst = 32'hc405012;
      37825: inst = 32'h8220000;
      37826: inst = 32'h10408000;
      37827: inst = 32'hc405013;
      37828: inst = 32'h8220000;
      37829: inst = 32'h10408000;
      37830: inst = 32'hc405014;
      37831: inst = 32'h8220000;
      37832: inst = 32'h10408000;
      37833: inst = 32'hc405015;
      37834: inst = 32'h8220000;
      37835: inst = 32'h10408000;
      37836: inst = 32'hc405016;
      37837: inst = 32'h8220000;
      37838: inst = 32'h10408000;
      37839: inst = 32'hc405017;
      37840: inst = 32'h8220000;
      37841: inst = 32'h10408000;
      37842: inst = 32'hc405018;
      37843: inst = 32'h8220000;
      37844: inst = 32'h10408000;
      37845: inst = 32'hc405019;
      37846: inst = 32'h8220000;
      37847: inst = 32'h10408000;
      37848: inst = 32'hc40501a;
      37849: inst = 32'h8220000;
      37850: inst = 32'h10408000;
      37851: inst = 32'hc40501b;
      37852: inst = 32'h8220000;
      37853: inst = 32'h10408000;
      37854: inst = 32'hc40501c;
      37855: inst = 32'h8220000;
      37856: inst = 32'h10408000;
      37857: inst = 32'hc40501d;
      37858: inst = 32'h8220000;
      37859: inst = 32'h10408000;
      37860: inst = 32'hc40501e;
      37861: inst = 32'h8220000;
      37862: inst = 32'h10408000;
      37863: inst = 32'hc40501f;
      37864: inst = 32'h8220000;
      37865: inst = 32'h10408000;
      37866: inst = 32'hc405020;
      37867: inst = 32'h8220000;
      37868: inst = 32'h10408000;
      37869: inst = 32'hc405021;
      37870: inst = 32'h8220000;
      37871: inst = 32'h10408000;
      37872: inst = 32'hc405022;
      37873: inst = 32'h8220000;
      37874: inst = 32'h10408000;
      37875: inst = 32'hc405023;
      37876: inst = 32'h8220000;
      37877: inst = 32'h10408000;
      37878: inst = 32'hc405024;
      37879: inst = 32'h8220000;
      37880: inst = 32'h10408000;
      37881: inst = 32'hc405025;
      37882: inst = 32'h8220000;
      37883: inst = 32'h10408000;
      37884: inst = 32'hc405026;
      37885: inst = 32'h8220000;
      37886: inst = 32'h10408000;
      37887: inst = 32'hc405027;
      37888: inst = 32'h8220000;
      37889: inst = 32'h10408000;
      37890: inst = 32'hc405028;
      37891: inst = 32'h8220000;
      37892: inst = 32'h10408000;
      37893: inst = 32'hc405029;
      37894: inst = 32'h8220000;
      37895: inst = 32'h10408000;
      37896: inst = 32'hc40502a;
      37897: inst = 32'h8220000;
      37898: inst = 32'h10408000;
      37899: inst = 32'hc40502b;
      37900: inst = 32'h8220000;
      37901: inst = 32'h10408000;
      37902: inst = 32'hc40502c;
      37903: inst = 32'h8220000;
      37904: inst = 32'h10408000;
      37905: inst = 32'hc40502d;
      37906: inst = 32'h8220000;
      37907: inst = 32'h10408000;
      37908: inst = 32'hc40502e;
      37909: inst = 32'h8220000;
      37910: inst = 32'h10408000;
      37911: inst = 32'hc40502f;
      37912: inst = 32'h8220000;
      37913: inst = 32'h10408000;
      37914: inst = 32'hc405030;
      37915: inst = 32'h8220000;
      37916: inst = 32'h10408000;
      37917: inst = 32'hc405031;
      37918: inst = 32'h8220000;
      37919: inst = 32'h10408000;
      37920: inst = 32'hc405032;
      37921: inst = 32'h8220000;
      37922: inst = 32'h10408000;
      37923: inst = 32'hc405033;
      37924: inst = 32'h8220000;
      37925: inst = 32'h10408000;
      37926: inst = 32'hc405034;
      37927: inst = 32'h8220000;
      37928: inst = 32'h10408000;
      37929: inst = 32'hc405035;
      37930: inst = 32'h8220000;
      37931: inst = 32'h10408000;
      37932: inst = 32'hc405036;
      37933: inst = 32'h8220000;
      37934: inst = 32'h10408000;
      37935: inst = 32'hc405037;
      37936: inst = 32'h8220000;
      37937: inst = 32'h10408000;
      37938: inst = 32'hc40503b;
      37939: inst = 32'h8220000;
      37940: inst = 32'h10408000;
      37941: inst = 32'hc40503c;
      37942: inst = 32'h8220000;
      37943: inst = 32'h10408000;
      37944: inst = 32'hc40503d;
      37945: inst = 32'h8220000;
      37946: inst = 32'h10408000;
      37947: inst = 32'hc40503e;
      37948: inst = 32'h8220000;
      37949: inst = 32'h10408000;
      37950: inst = 32'hc40503f;
      37951: inst = 32'h8220000;
      37952: inst = 32'h10408000;
      37953: inst = 32'hc405040;
      37954: inst = 32'h8220000;
      37955: inst = 32'h10408000;
      37956: inst = 32'hc405041;
      37957: inst = 32'h8220000;
      37958: inst = 32'h10408000;
      37959: inst = 32'hc405042;
      37960: inst = 32'h8220000;
      37961: inst = 32'h10408000;
      37962: inst = 32'hc405043;
      37963: inst = 32'h8220000;
      37964: inst = 32'h10408000;
      37965: inst = 32'hc405044;
      37966: inst = 32'h8220000;
      37967: inst = 32'h10408000;
      37968: inst = 32'hc405045;
      37969: inst = 32'h8220000;
      37970: inst = 32'h10408000;
      37971: inst = 32'hc405046;
      37972: inst = 32'h8220000;
      37973: inst = 32'h10408000;
      37974: inst = 32'hc405047;
      37975: inst = 32'h8220000;
      37976: inst = 32'h10408000;
      37977: inst = 32'hc405048;
      37978: inst = 32'h8220000;
      37979: inst = 32'h10408000;
      37980: inst = 32'hc405049;
      37981: inst = 32'h8220000;
      37982: inst = 32'h10408000;
      37983: inst = 32'hc40504a;
      37984: inst = 32'h8220000;
      37985: inst = 32'h10408000;
      37986: inst = 32'hc40504b;
      37987: inst = 32'h8220000;
      37988: inst = 32'h10408000;
      37989: inst = 32'hc40504c;
      37990: inst = 32'h8220000;
      37991: inst = 32'h10408000;
      37992: inst = 32'hc40504d;
      37993: inst = 32'h8220000;
      37994: inst = 32'h10408000;
      37995: inst = 32'hc40504e;
      37996: inst = 32'h8220000;
      37997: inst = 32'h10408000;
      37998: inst = 32'hc40504f;
      37999: inst = 32'h8220000;
      38000: inst = 32'h10408000;
      38001: inst = 32'hc405050;
      38002: inst = 32'h8220000;
      38003: inst = 32'h10408000;
      38004: inst = 32'hc405051;
      38005: inst = 32'h8220000;
      38006: inst = 32'h10408000;
      38007: inst = 32'hc405052;
      38008: inst = 32'h8220000;
      38009: inst = 32'h10408000;
      38010: inst = 32'hc405053;
      38011: inst = 32'h8220000;
      38012: inst = 32'h10408000;
      38013: inst = 32'hc405054;
      38014: inst = 32'h8220000;
      38015: inst = 32'h10408000;
      38016: inst = 32'hc405055;
      38017: inst = 32'h8220000;
      38018: inst = 32'h10408000;
      38019: inst = 32'hc405056;
      38020: inst = 32'h8220000;
      38021: inst = 32'h10408000;
      38022: inst = 32'hc405057;
      38023: inst = 32'h8220000;
      38024: inst = 32'h10408000;
      38025: inst = 32'hc405058;
      38026: inst = 32'h8220000;
      38027: inst = 32'h10408000;
      38028: inst = 32'hc405059;
      38029: inst = 32'h8220000;
      38030: inst = 32'h10408000;
      38031: inst = 32'hc40505a;
      38032: inst = 32'h8220000;
      38033: inst = 32'h10408000;
      38034: inst = 32'hc40505b;
      38035: inst = 32'h8220000;
      38036: inst = 32'h10408000;
      38037: inst = 32'hc40505c;
      38038: inst = 32'h8220000;
      38039: inst = 32'h10408000;
      38040: inst = 32'hc405063;
      38041: inst = 32'h8220000;
      38042: inst = 32'h10408000;
      38043: inst = 32'hc405064;
      38044: inst = 32'h8220000;
      38045: inst = 32'h10408000;
      38046: inst = 32'hc405065;
      38047: inst = 32'h8220000;
      38048: inst = 32'h10408000;
      38049: inst = 32'hc405066;
      38050: inst = 32'h8220000;
      38051: inst = 32'h10408000;
      38052: inst = 32'hc405067;
      38053: inst = 32'h8220000;
      38054: inst = 32'h10408000;
      38055: inst = 32'hc405068;
      38056: inst = 32'h8220000;
      38057: inst = 32'h10408000;
      38058: inst = 32'hc405069;
      38059: inst = 32'h8220000;
      38060: inst = 32'h10408000;
      38061: inst = 32'hc40506a;
      38062: inst = 32'h8220000;
      38063: inst = 32'h10408000;
      38064: inst = 32'hc40506b;
      38065: inst = 32'h8220000;
      38066: inst = 32'h10408000;
      38067: inst = 32'hc40506c;
      38068: inst = 32'h8220000;
      38069: inst = 32'h10408000;
      38070: inst = 32'hc40506d;
      38071: inst = 32'h8220000;
      38072: inst = 32'h10408000;
      38073: inst = 32'hc40506e;
      38074: inst = 32'h8220000;
      38075: inst = 32'h10408000;
      38076: inst = 32'hc40506f;
      38077: inst = 32'h8220000;
      38078: inst = 32'h10408000;
      38079: inst = 32'hc405070;
      38080: inst = 32'h8220000;
      38081: inst = 32'h10408000;
      38082: inst = 32'hc405071;
      38083: inst = 32'h8220000;
      38084: inst = 32'h10408000;
      38085: inst = 32'hc405072;
      38086: inst = 32'h8220000;
      38087: inst = 32'h10408000;
      38088: inst = 32'hc405073;
      38089: inst = 32'h8220000;
      38090: inst = 32'h10408000;
      38091: inst = 32'hc405074;
      38092: inst = 32'h8220000;
      38093: inst = 32'h10408000;
      38094: inst = 32'hc405075;
      38095: inst = 32'h8220000;
      38096: inst = 32'h10408000;
      38097: inst = 32'hc405076;
      38098: inst = 32'h8220000;
      38099: inst = 32'h10408000;
      38100: inst = 32'hc405077;
      38101: inst = 32'h8220000;
      38102: inst = 32'h10408000;
      38103: inst = 32'hc405078;
      38104: inst = 32'h8220000;
      38105: inst = 32'h10408000;
      38106: inst = 32'hc405079;
      38107: inst = 32'h8220000;
      38108: inst = 32'h10408000;
      38109: inst = 32'hc40507a;
      38110: inst = 32'h8220000;
      38111: inst = 32'h10408000;
      38112: inst = 32'hc40507b;
      38113: inst = 32'h8220000;
      38114: inst = 32'h10408000;
      38115: inst = 32'hc40507c;
      38116: inst = 32'h8220000;
      38117: inst = 32'h10408000;
      38118: inst = 32'hc40507d;
      38119: inst = 32'h8220000;
      38120: inst = 32'h10408000;
      38121: inst = 32'hc40507e;
      38122: inst = 32'h8220000;
      38123: inst = 32'h10408000;
      38124: inst = 32'hc40507f;
      38125: inst = 32'h8220000;
      38126: inst = 32'h10408000;
      38127: inst = 32'hc405080;
      38128: inst = 32'h8220000;
      38129: inst = 32'h10408000;
      38130: inst = 32'hc405081;
      38131: inst = 32'h8220000;
      38132: inst = 32'h10408000;
      38133: inst = 32'hc405082;
      38134: inst = 32'h8220000;
      38135: inst = 32'h10408000;
      38136: inst = 32'hc405083;
      38137: inst = 32'h8220000;
      38138: inst = 32'h10408000;
      38139: inst = 32'hc405084;
      38140: inst = 32'h8220000;
      38141: inst = 32'h10408000;
      38142: inst = 32'hc405085;
      38143: inst = 32'h8220000;
      38144: inst = 32'h10408000;
      38145: inst = 32'hc405086;
      38146: inst = 32'h8220000;
      38147: inst = 32'h10408000;
      38148: inst = 32'hc405087;
      38149: inst = 32'h8220000;
      38150: inst = 32'h10408000;
      38151: inst = 32'hc405088;
      38152: inst = 32'h8220000;
      38153: inst = 32'h10408000;
      38154: inst = 32'hc405089;
      38155: inst = 32'h8220000;
      38156: inst = 32'h10408000;
      38157: inst = 32'hc40508a;
      38158: inst = 32'h8220000;
      38159: inst = 32'h10408000;
      38160: inst = 32'hc40508b;
      38161: inst = 32'h8220000;
      38162: inst = 32'h10408000;
      38163: inst = 32'hc40508c;
      38164: inst = 32'h8220000;
      38165: inst = 32'h10408000;
      38166: inst = 32'hc40508d;
      38167: inst = 32'h8220000;
      38168: inst = 32'h10408000;
      38169: inst = 32'hc40508e;
      38170: inst = 32'h8220000;
      38171: inst = 32'h10408000;
      38172: inst = 32'hc40508f;
      38173: inst = 32'h8220000;
      38174: inst = 32'h10408000;
      38175: inst = 32'hc405090;
      38176: inst = 32'h8220000;
      38177: inst = 32'h10408000;
      38178: inst = 32'hc405091;
      38179: inst = 32'h8220000;
      38180: inst = 32'h10408000;
      38181: inst = 32'hc405092;
      38182: inst = 32'h8220000;
      38183: inst = 32'h10408000;
      38184: inst = 32'hc405093;
      38185: inst = 32'h8220000;
      38186: inst = 32'h10408000;
      38187: inst = 32'hc405094;
      38188: inst = 32'h8220000;
      38189: inst = 32'h10408000;
      38190: inst = 32'hc405095;
      38191: inst = 32'h8220000;
      38192: inst = 32'h10408000;
      38193: inst = 32'hc405096;
      38194: inst = 32'h8220000;
      38195: inst = 32'h10408000;
      38196: inst = 32'hc405097;
      38197: inst = 32'h8220000;
      38198: inst = 32'h10408000;
      38199: inst = 32'hc4050c3;
      38200: inst = 32'h8220000;
      38201: inst = 32'h10408000;
      38202: inst = 32'hc4050c4;
      38203: inst = 32'h8220000;
      38204: inst = 32'h10408000;
      38205: inst = 32'hc4050c5;
      38206: inst = 32'h8220000;
      38207: inst = 32'h10408000;
      38208: inst = 32'hc4050c6;
      38209: inst = 32'h8220000;
      38210: inst = 32'h10408000;
      38211: inst = 32'hc4050c7;
      38212: inst = 32'h8220000;
      38213: inst = 32'h10408000;
      38214: inst = 32'hc4050c8;
      38215: inst = 32'h8220000;
      38216: inst = 32'h10408000;
      38217: inst = 32'hc4050c9;
      38218: inst = 32'h8220000;
      38219: inst = 32'h10408000;
      38220: inst = 32'hc4050ca;
      38221: inst = 32'h8220000;
      38222: inst = 32'h10408000;
      38223: inst = 32'hc4050cb;
      38224: inst = 32'h8220000;
      38225: inst = 32'h10408000;
      38226: inst = 32'hc4050cc;
      38227: inst = 32'h8220000;
      38228: inst = 32'h10408000;
      38229: inst = 32'hc4050cd;
      38230: inst = 32'h8220000;
      38231: inst = 32'h10408000;
      38232: inst = 32'hc4050ce;
      38233: inst = 32'h8220000;
      38234: inst = 32'h10408000;
      38235: inst = 32'hc4050cf;
      38236: inst = 32'h8220000;
      38237: inst = 32'h10408000;
      38238: inst = 32'hc4050d0;
      38239: inst = 32'h8220000;
      38240: inst = 32'h10408000;
      38241: inst = 32'hc4050d1;
      38242: inst = 32'h8220000;
      38243: inst = 32'h10408000;
      38244: inst = 32'hc4050d2;
      38245: inst = 32'h8220000;
      38246: inst = 32'h10408000;
      38247: inst = 32'hc4050d3;
      38248: inst = 32'h8220000;
      38249: inst = 32'h10408000;
      38250: inst = 32'hc4050d4;
      38251: inst = 32'h8220000;
      38252: inst = 32'h10408000;
      38253: inst = 32'hc4050d5;
      38254: inst = 32'h8220000;
      38255: inst = 32'h10408000;
      38256: inst = 32'hc4050d6;
      38257: inst = 32'h8220000;
      38258: inst = 32'h10408000;
      38259: inst = 32'hc4050d7;
      38260: inst = 32'h8220000;
      38261: inst = 32'h10408000;
      38262: inst = 32'hc4050d8;
      38263: inst = 32'h8220000;
      38264: inst = 32'h10408000;
      38265: inst = 32'hc4050d9;
      38266: inst = 32'h8220000;
      38267: inst = 32'h10408000;
      38268: inst = 32'hc4050da;
      38269: inst = 32'h8220000;
      38270: inst = 32'h10408000;
      38271: inst = 32'hc4050db;
      38272: inst = 32'h8220000;
      38273: inst = 32'h10408000;
      38274: inst = 32'hc4050dc;
      38275: inst = 32'h8220000;
      38276: inst = 32'h10408000;
      38277: inst = 32'hc4050dd;
      38278: inst = 32'h8220000;
      38279: inst = 32'h10408000;
      38280: inst = 32'hc4050de;
      38281: inst = 32'h8220000;
      38282: inst = 32'h10408000;
      38283: inst = 32'hc4050df;
      38284: inst = 32'h8220000;
      38285: inst = 32'h10408000;
      38286: inst = 32'hc4050e0;
      38287: inst = 32'h8220000;
      38288: inst = 32'h10408000;
      38289: inst = 32'hc4050e1;
      38290: inst = 32'h8220000;
      38291: inst = 32'h10408000;
      38292: inst = 32'hc4050e2;
      38293: inst = 32'h8220000;
      38294: inst = 32'h10408000;
      38295: inst = 32'hc4050e3;
      38296: inst = 32'h8220000;
      38297: inst = 32'h10408000;
      38298: inst = 32'hc4050e4;
      38299: inst = 32'h8220000;
      38300: inst = 32'h10408000;
      38301: inst = 32'hc4050e5;
      38302: inst = 32'h8220000;
      38303: inst = 32'h10408000;
      38304: inst = 32'hc4050e6;
      38305: inst = 32'h8220000;
      38306: inst = 32'h10408000;
      38307: inst = 32'hc4050e7;
      38308: inst = 32'h8220000;
      38309: inst = 32'h10408000;
      38310: inst = 32'hc4050e8;
      38311: inst = 32'h8220000;
      38312: inst = 32'h10408000;
      38313: inst = 32'hc4050e9;
      38314: inst = 32'h8220000;
      38315: inst = 32'h10408000;
      38316: inst = 32'hc4050ea;
      38317: inst = 32'h8220000;
      38318: inst = 32'h10408000;
      38319: inst = 32'hc4050eb;
      38320: inst = 32'h8220000;
      38321: inst = 32'h10408000;
      38322: inst = 32'hc4050ec;
      38323: inst = 32'h8220000;
      38324: inst = 32'h10408000;
      38325: inst = 32'hc4050ed;
      38326: inst = 32'h8220000;
      38327: inst = 32'h10408000;
      38328: inst = 32'hc4050ee;
      38329: inst = 32'h8220000;
      38330: inst = 32'h10408000;
      38331: inst = 32'hc4050ef;
      38332: inst = 32'h8220000;
      38333: inst = 32'h10408000;
      38334: inst = 32'hc4050f0;
      38335: inst = 32'h8220000;
      38336: inst = 32'h10408000;
      38337: inst = 32'hc4050f1;
      38338: inst = 32'h8220000;
      38339: inst = 32'h10408000;
      38340: inst = 32'hc4050f2;
      38341: inst = 32'h8220000;
      38342: inst = 32'h10408000;
      38343: inst = 32'hc4050f3;
      38344: inst = 32'h8220000;
      38345: inst = 32'h10408000;
      38346: inst = 32'hc4050f4;
      38347: inst = 32'h8220000;
      38348: inst = 32'h10408000;
      38349: inst = 32'hc4050f5;
      38350: inst = 32'h8220000;
      38351: inst = 32'h10408000;
      38352: inst = 32'hc4050f6;
      38353: inst = 32'h8220000;
      38354: inst = 32'h10408000;
      38355: inst = 32'hc4050f7;
      38356: inst = 32'h8220000;
      38357: inst = 32'h10408000;
      38358: inst = 32'hc405123;
      38359: inst = 32'h8220000;
      38360: inst = 32'h10408000;
      38361: inst = 32'hc405124;
      38362: inst = 32'h8220000;
      38363: inst = 32'h10408000;
      38364: inst = 32'hc405125;
      38365: inst = 32'h8220000;
      38366: inst = 32'h10408000;
      38367: inst = 32'hc405126;
      38368: inst = 32'h8220000;
      38369: inst = 32'h10408000;
      38370: inst = 32'hc405127;
      38371: inst = 32'h8220000;
      38372: inst = 32'h10408000;
      38373: inst = 32'hc405128;
      38374: inst = 32'h8220000;
      38375: inst = 32'h10408000;
      38376: inst = 32'hc405129;
      38377: inst = 32'h8220000;
      38378: inst = 32'h10408000;
      38379: inst = 32'hc40512a;
      38380: inst = 32'h8220000;
      38381: inst = 32'h10408000;
      38382: inst = 32'hc40512b;
      38383: inst = 32'h8220000;
      38384: inst = 32'h10408000;
      38385: inst = 32'hc40512c;
      38386: inst = 32'h8220000;
      38387: inst = 32'h10408000;
      38388: inst = 32'hc40512d;
      38389: inst = 32'h8220000;
      38390: inst = 32'h10408000;
      38391: inst = 32'hc40512e;
      38392: inst = 32'h8220000;
      38393: inst = 32'h10408000;
      38394: inst = 32'hc40512f;
      38395: inst = 32'h8220000;
      38396: inst = 32'h10408000;
      38397: inst = 32'hc405130;
      38398: inst = 32'h8220000;
      38399: inst = 32'h10408000;
      38400: inst = 32'hc405131;
      38401: inst = 32'h8220000;
      38402: inst = 32'h10408000;
      38403: inst = 32'hc405132;
      38404: inst = 32'h8220000;
      38405: inst = 32'h10408000;
      38406: inst = 32'hc405133;
      38407: inst = 32'h8220000;
      38408: inst = 32'h10408000;
      38409: inst = 32'hc405134;
      38410: inst = 32'h8220000;
      38411: inst = 32'h10408000;
      38412: inst = 32'hc405135;
      38413: inst = 32'h8220000;
      38414: inst = 32'h10408000;
      38415: inst = 32'hc405139;
      38416: inst = 32'h8220000;
      38417: inst = 32'h10408000;
      38418: inst = 32'hc40513a;
      38419: inst = 32'h8220000;
      38420: inst = 32'h10408000;
      38421: inst = 32'hc40513b;
      38422: inst = 32'h8220000;
      38423: inst = 32'h10408000;
      38424: inst = 32'hc40513c;
      38425: inst = 32'h8220000;
      38426: inst = 32'h10408000;
      38427: inst = 32'hc40513d;
      38428: inst = 32'h8220000;
      38429: inst = 32'h10408000;
      38430: inst = 32'hc40513e;
      38431: inst = 32'h8220000;
      38432: inst = 32'h10408000;
      38433: inst = 32'hc40513f;
      38434: inst = 32'h8220000;
      38435: inst = 32'h10408000;
      38436: inst = 32'hc405140;
      38437: inst = 32'h8220000;
      38438: inst = 32'h10408000;
      38439: inst = 32'hc405141;
      38440: inst = 32'h8220000;
      38441: inst = 32'h10408000;
      38442: inst = 32'hc405142;
      38443: inst = 32'h8220000;
      38444: inst = 32'h10408000;
      38445: inst = 32'hc405143;
      38446: inst = 32'h8220000;
      38447: inst = 32'h10408000;
      38448: inst = 32'hc405144;
      38449: inst = 32'h8220000;
      38450: inst = 32'h10408000;
      38451: inst = 32'hc405145;
      38452: inst = 32'h8220000;
      38453: inst = 32'h10408000;
      38454: inst = 32'hc405146;
      38455: inst = 32'h8220000;
      38456: inst = 32'h10408000;
      38457: inst = 32'hc405147;
      38458: inst = 32'h8220000;
      38459: inst = 32'h10408000;
      38460: inst = 32'hc405148;
      38461: inst = 32'h8220000;
      38462: inst = 32'h10408000;
      38463: inst = 32'hc405149;
      38464: inst = 32'h8220000;
      38465: inst = 32'h10408000;
      38466: inst = 32'hc40514a;
      38467: inst = 32'h8220000;
      38468: inst = 32'h10408000;
      38469: inst = 32'hc40514b;
      38470: inst = 32'h8220000;
      38471: inst = 32'h10408000;
      38472: inst = 32'hc40514c;
      38473: inst = 32'h8220000;
      38474: inst = 32'h10408000;
      38475: inst = 32'hc40514d;
      38476: inst = 32'h8220000;
      38477: inst = 32'h10408000;
      38478: inst = 32'hc40514e;
      38479: inst = 32'h8220000;
      38480: inst = 32'h10408000;
      38481: inst = 32'hc40514f;
      38482: inst = 32'h8220000;
      38483: inst = 32'h10408000;
      38484: inst = 32'hc405150;
      38485: inst = 32'h8220000;
      38486: inst = 32'h10408000;
      38487: inst = 32'hc405151;
      38488: inst = 32'h8220000;
      38489: inst = 32'h10408000;
      38490: inst = 32'hc405152;
      38491: inst = 32'h8220000;
      38492: inst = 32'h10408000;
      38493: inst = 32'hc405153;
      38494: inst = 32'h8220000;
      38495: inst = 32'h10408000;
      38496: inst = 32'hc405154;
      38497: inst = 32'h8220000;
      38498: inst = 32'h10408000;
      38499: inst = 32'hc405155;
      38500: inst = 32'h8220000;
      38501: inst = 32'h10408000;
      38502: inst = 32'hc405156;
      38503: inst = 32'h8220000;
      38504: inst = 32'h10408000;
      38505: inst = 32'hc405157;
      38506: inst = 32'h8220000;
      38507: inst = 32'h10408000;
      38508: inst = 32'hc405183;
      38509: inst = 32'h8220000;
      38510: inst = 32'h10408000;
      38511: inst = 32'hc405184;
      38512: inst = 32'h8220000;
      38513: inst = 32'h10408000;
      38514: inst = 32'hc405185;
      38515: inst = 32'h8220000;
      38516: inst = 32'h10408000;
      38517: inst = 32'hc405186;
      38518: inst = 32'h8220000;
      38519: inst = 32'h10408000;
      38520: inst = 32'hc405187;
      38521: inst = 32'h8220000;
      38522: inst = 32'h10408000;
      38523: inst = 32'hc405188;
      38524: inst = 32'h8220000;
      38525: inst = 32'h10408000;
      38526: inst = 32'hc405189;
      38527: inst = 32'h8220000;
      38528: inst = 32'h10408000;
      38529: inst = 32'hc40518a;
      38530: inst = 32'h8220000;
      38531: inst = 32'h10408000;
      38532: inst = 32'hc40518b;
      38533: inst = 32'h8220000;
      38534: inst = 32'h10408000;
      38535: inst = 32'hc40518c;
      38536: inst = 32'h8220000;
      38537: inst = 32'h10408000;
      38538: inst = 32'hc40518d;
      38539: inst = 32'h8220000;
      38540: inst = 32'h10408000;
      38541: inst = 32'hc40518e;
      38542: inst = 32'h8220000;
      38543: inst = 32'h10408000;
      38544: inst = 32'hc40518f;
      38545: inst = 32'h8220000;
      38546: inst = 32'h10408000;
      38547: inst = 32'hc405190;
      38548: inst = 32'h8220000;
      38549: inst = 32'h10408000;
      38550: inst = 32'hc405191;
      38551: inst = 32'h8220000;
      38552: inst = 32'h10408000;
      38553: inst = 32'hc405192;
      38554: inst = 32'h8220000;
      38555: inst = 32'h10408000;
      38556: inst = 32'hc405193;
      38557: inst = 32'h8220000;
      38558: inst = 32'h10408000;
      38559: inst = 32'hc405194;
      38560: inst = 32'h8220000;
      38561: inst = 32'h10408000;
      38562: inst = 32'hc405195;
      38563: inst = 32'h8220000;
      38564: inst = 32'h10408000;
      38565: inst = 32'hc405199;
      38566: inst = 32'h8220000;
      38567: inst = 32'h10408000;
      38568: inst = 32'hc40519a;
      38569: inst = 32'h8220000;
      38570: inst = 32'h10408000;
      38571: inst = 32'hc40519b;
      38572: inst = 32'h8220000;
      38573: inst = 32'h10408000;
      38574: inst = 32'hc40519c;
      38575: inst = 32'h8220000;
      38576: inst = 32'h10408000;
      38577: inst = 32'hc40519d;
      38578: inst = 32'h8220000;
      38579: inst = 32'h10408000;
      38580: inst = 32'hc40519e;
      38581: inst = 32'h8220000;
      38582: inst = 32'h10408000;
      38583: inst = 32'hc40519f;
      38584: inst = 32'h8220000;
      38585: inst = 32'h10408000;
      38586: inst = 32'hc4051a0;
      38587: inst = 32'h8220000;
      38588: inst = 32'h10408000;
      38589: inst = 32'hc4051a1;
      38590: inst = 32'h8220000;
      38591: inst = 32'h10408000;
      38592: inst = 32'hc4051a2;
      38593: inst = 32'h8220000;
      38594: inst = 32'h10408000;
      38595: inst = 32'hc4051a3;
      38596: inst = 32'h8220000;
      38597: inst = 32'h10408000;
      38598: inst = 32'hc4051a4;
      38599: inst = 32'h8220000;
      38600: inst = 32'h10408000;
      38601: inst = 32'hc4051a5;
      38602: inst = 32'h8220000;
      38603: inst = 32'h10408000;
      38604: inst = 32'hc4051a6;
      38605: inst = 32'h8220000;
      38606: inst = 32'h10408000;
      38607: inst = 32'hc4051a7;
      38608: inst = 32'h8220000;
      38609: inst = 32'h10408000;
      38610: inst = 32'hc4051a8;
      38611: inst = 32'h8220000;
      38612: inst = 32'h10408000;
      38613: inst = 32'hc4051a9;
      38614: inst = 32'h8220000;
      38615: inst = 32'h10408000;
      38616: inst = 32'hc4051aa;
      38617: inst = 32'h8220000;
      38618: inst = 32'h10408000;
      38619: inst = 32'hc4051ab;
      38620: inst = 32'h8220000;
      38621: inst = 32'h10408000;
      38622: inst = 32'hc4051ac;
      38623: inst = 32'h8220000;
      38624: inst = 32'h10408000;
      38625: inst = 32'hc4051ad;
      38626: inst = 32'h8220000;
      38627: inst = 32'h10408000;
      38628: inst = 32'hc4051ae;
      38629: inst = 32'h8220000;
      38630: inst = 32'h10408000;
      38631: inst = 32'hc4051af;
      38632: inst = 32'h8220000;
      38633: inst = 32'h10408000;
      38634: inst = 32'hc4051b0;
      38635: inst = 32'h8220000;
      38636: inst = 32'h10408000;
      38637: inst = 32'hc4051b1;
      38638: inst = 32'h8220000;
      38639: inst = 32'h10408000;
      38640: inst = 32'hc4051b2;
      38641: inst = 32'h8220000;
      38642: inst = 32'h10408000;
      38643: inst = 32'hc4051b3;
      38644: inst = 32'h8220000;
      38645: inst = 32'h10408000;
      38646: inst = 32'hc4051b4;
      38647: inst = 32'h8220000;
      38648: inst = 32'h10408000;
      38649: inst = 32'hc4051b5;
      38650: inst = 32'h8220000;
      38651: inst = 32'h10408000;
      38652: inst = 32'hc4051b6;
      38653: inst = 32'h8220000;
      38654: inst = 32'h10408000;
      38655: inst = 32'hc4051b7;
      38656: inst = 32'h8220000;
      38657: inst = 32'h10408000;
      38658: inst = 32'hc4051b8;
      38659: inst = 32'h8220000;
      38660: inst = 32'h10408000;
      38661: inst = 32'hc4051b9;
      38662: inst = 32'h8220000;
      38663: inst = 32'h10408000;
      38664: inst = 32'hc4051ba;
      38665: inst = 32'h8220000;
      38666: inst = 32'h10408000;
      38667: inst = 32'hc4051bb;
      38668: inst = 32'h8220000;
      38669: inst = 32'h10408000;
      38670: inst = 32'hc4051bc;
      38671: inst = 32'h8220000;
      38672: inst = 32'h10408000;
      38673: inst = 32'hc4051bd;
      38674: inst = 32'h8220000;
      38675: inst = 32'h10408000;
      38676: inst = 32'hc4051be;
      38677: inst = 32'h8220000;
      38678: inst = 32'h10408000;
      38679: inst = 32'hc4051bf;
      38680: inst = 32'h8220000;
      38681: inst = 32'h10408000;
      38682: inst = 32'hc4051c0;
      38683: inst = 32'h8220000;
      38684: inst = 32'h10408000;
      38685: inst = 32'hc4051c1;
      38686: inst = 32'h8220000;
      38687: inst = 32'h10408000;
      38688: inst = 32'hc4051c2;
      38689: inst = 32'h8220000;
      38690: inst = 32'h10408000;
      38691: inst = 32'hc4051c3;
      38692: inst = 32'h8220000;
      38693: inst = 32'h10408000;
      38694: inst = 32'hc4051c4;
      38695: inst = 32'h8220000;
      38696: inst = 32'h10408000;
      38697: inst = 32'hc4051c5;
      38698: inst = 32'h8220000;
      38699: inst = 32'h10408000;
      38700: inst = 32'hc4051c6;
      38701: inst = 32'h8220000;
      38702: inst = 32'h10408000;
      38703: inst = 32'hc4051c7;
      38704: inst = 32'h8220000;
      38705: inst = 32'h10408000;
      38706: inst = 32'hc4051c8;
      38707: inst = 32'h8220000;
      38708: inst = 32'h10408000;
      38709: inst = 32'hc4051c9;
      38710: inst = 32'h8220000;
      38711: inst = 32'h10408000;
      38712: inst = 32'hc4051ca;
      38713: inst = 32'h8220000;
      38714: inst = 32'h10408000;
      38715: inst = 32'hc4051cb;
      38716: inst = 32'h8220000;
      38717: inst = 32'h10408000;
      38718: inst = 32'hc4051cc;
      38719: inst = 32'h8220000;
      38720: inst = 32'h10408000;
      38721: inst = 32'hc4051cd;
      38722: inst = 32'h8220000;
      38723: inst = 32'h10408000;
      38724: inst = 32'hc4051ce;
      38725: inst = 32'h8220000;
      38726: inst = 32'h10408000;
      38727: inst = 32'hc4051cf;
      38728: inst = 32'h8220000;
      38729: inst = 32'h10408000;
      38730: inst = 32'hc4051d0;
      38731: inst = 32'h8220000;
      38732: inst = 32'h10408000;
      38733: inst = 32'hc4051d1;
      38734: inst = 32'h8220000;
      38735: inst = 32'h10408000;
      38736: inst = 32'hc4051d2;
      38737: inst = 32'h8220000;
      38738: inst = 32'h10408000;
      38739: inst = 32'hc4051d3;
      38740: inst = 32'h8220000;
      38741: inst = 32'h10408000;
      38742: inst = 32'hc4051d4;
      38743: inst = 32'h8220000;
      38744: inst = 32'h10408000;
      38745: inst = 32'hc4051d5;
      38746: inst = 32'h8220000;
      38747: inst = 32'h10408000;
      38748: inst = 32'hc4051d6;
      38749: inst = 32'h8220000;
      38750: inst = 32'h10408000;
      38751: inst = 32'hc4051d7;
      38752: inst = 32'h8220000;
      38753: inst = 32'h10408000;
      38754: inst = 32'hc4051d8;
      38755: inst = 32'h8220000;
      38756: inst = 32'h10408000;
      38757: inst = 32'hc4051d9;
      38758: inst = 32'h8220000;
      38759: inst = 32'h10408000;
      38760: inst = 32'hc4051da;
      38761: inst = 32'h8220000;
      38762: inst = 32'h10408000;
      38763: inst = 32'hc4051db;
      38764: inst = 32'h8220000;
      38765: inst = 32'h10408000;
      38766: inst = 32'hc4051dc;
      38767: inst = 32'h8220000;
      38768: inst = 32'h10408000;
      38769: inst = 32'hc4051e3;
      38770: inst = 32'h8220000;
      38771: inst = 32'h10408000;
      38772: inst = 32'hc4051e4;
      38773: inst = 32'h8220000;
      38774: inst = 32'h10408000;
      38775: inst = 32'hc4051e5;
      38776: inst = 32'h8220000;
      38777: inst = 32'h10408000;
      38778: inst = 32'hc4051e6;
      38779: inst = 32'h8220000;
      38780: inst = 32'h10408000;
      38781: inst = 32'hc4051e7;
      38782: inst = 32'h8220000;
      38783: inst = 32'h10408000;
      38784: inst = 32'hc4051e8;
      38785: inst = 32'h8220000;
      38786: inst = 32'h10408000;
      38787: inst = 32'hc4051e9;
      38788: inst = 32'h8220000;
      38789: inst = 32'h10408000;
      38790: inst = 32'hc4051ea;
      38791: inst = 32'h8220000;
      38792: inst = 32'h10408000;
      38793: inst = 32'hc4051eb;
      38794: inst = 32'h8220000;
      38795: inst = 32'h10408000;
      38796: inst = 32'hc4051ec;
      38797: inst = 32'h8220000;
      38798: inst = 32'h10408000;
      38799: inst = 32'hc4051ed;
      38800: inst = 32'h8220000;
      38801: inst = 32'h10408000;
      38802: inst = 32'hc4051ee;
      38803: inst = 32'h8220000;
      38804: inst = 32'h10408000;
      38805: inst = 32'hc4051ef;
      38806: inst = 32'h8220000;
      38807: inst = 32'h10408000;
      38808: inst = 32'hc4051f0;
      38809: inst = 32'h8220000;
      38810: inst = 32'h10408000;
      38811: inst = 32'hc4051f1;
      38812: inst = 32'h8220000;
      38813: inst = 32'h10408000;
      38814: inst = 32'hc4051f2;
      38815: inst = 32'h8220000;
      38816: inst = 32'h10408000;
      38817: inst = 32'hc4051f3;
      38818: inst = 32'h8220000;
      38819: inst = 32'h10408000;
      38820: inst = 32'hc4051f4;
      38821: inst = 32'h8220000;
      38822: inst = 32'h10408000;
      38823: inst = 32'hc4051f5;
      38824: inst = 32'h8220000;
      38825: inst = 32'h10408000;
      38826: inst = 32'hc4051f9;
      38827: inst = 32'h8220000;
      38828: inst = 32'h10408000;
      38829: inst = 32'hc4051fa;
      38830: inst = 32'h8220000;
      38831: inst = 32'h10408000;
      38832: inst = 32'hc4051fb;
      38833: inst = 32'h8220000;
      38834: inst = 32'h10408000;
      38835: inst = 32'hc4051fc;
      38836: inst = 32'h8220000;
      38837: inst = 32'h10408000;
      38838: inst = 32'hc4051fd;
      38839: inst = 32'h8220000;
      38840: inst = 32'h10408000;
      38841: inst = 32'hc4051fe;
      38842: inst = 32'h8220000;
      38843: inst = 32'h10408000;
      38844: inst = 32'hc4051ff;
      38845: inst = 32'h8220000;
      38846: inst = 32'h10408000;
      38847: inst = 32'hc405200;
      38848: inst = 32'h8220000;
      38849: inst = 32'h10408000;
      38850: inst = 32'hc405201;
      38851: inst = 32'h8220000;
      38852: inst = 32'h10408000;
      38853: inst = 32'hc405202;
      38854: inst = 32'h8220000;
      38855: inst = 32'h10408000;
      38856: inst = 32'hc405203;
      38857: inst = 32'h8220000;
      38858: inst = 32'h10408000;
      38859: inst = 32'hc405204;
      38860: inst = 32'h8220000;
      38861: inst = 32'h10408000;
      38862: inst = 32'hc405205;
      38863: inst = 32'h8220000;
      38864: inst = 32'h10408000;
      38865: inst = 32'hc405206;
      38866: inst = 32'h8220000;
      38867: inst = 32'h10408000;
      38868: inst = 32'hc405207;
      38869: inst = 32'h8220000;
      38870: inst = 32'h10408000;
      38871: inst = 32'hc405208;
      38872: inst = 32'h8220000;
      38873: inst = 32'h10408000;
      38874: inst = 32'hc405209;
      38875: inst = 32'h8220000;
      38876: inst = 32'h10408000;
      38877: inst = 32'hc40520a;
      38878: inst = 32'h8220000;
      38879: inst = 32'h10408000;
      38880: inst = 32'hc40520b;
      38881: inst = 32'h8220000;
      38882: inst = 32'h10408000;
      38883: inst = 32'hc40520c;
      38884: inst = 32'h8220000;
      38885: inst = 32'h10408000;
      38886: inst = 32'hc40520d;
      38887: inst = 32'h8220000;
      38888: inst = 32'h10408000;
      38889: inst = 32'hc40520e;
      38890: inst = 32'h8220000;
      38891: inst = 32'h10408000;
      38892: inst = 32'hc40520f;
      38893: inst = 32'h8220000;
      38894: inst = 32'h10408000;
      38895: inst = 32'hc405210;
      38896: inst = 32'h8220000;
      38897: inst = 32'h10408000;
      38898: inst = 32'hc405211;
      38899: inst = 32'h8220000;
      38900: inst = 32'h10408000;
      38901: inst = 32'hc405212;
      38902: inst = 32'h8220000;
      38903: inst = 32'h10408000;
      38904: inst = 32'hc405213;
      38905: inst = 32'h8220000;
      38906: inst = 32'h10408000;
      38907: inst = 32'hc405214;
      38908: inst = 32'h8220000;
      38909: inst = 32'h10408000;
      38910: inst = 32'hc405215;
      38911: inst = 32'h8220000;
      38912: inst = 32'h10408000;
      38913: inst = 32'hc405216;
      38914: inst = 32'h8220000;
      38915: inst = 32'h10408000;
      38916: inst = 32'hc405217;
      38917: inst = 32'h8220000;
      38918: inst = 32'h10408000;
      38919: inst = 32'hc405218;
      38920: inst = 32'h8220000;
      38921: inst = 32'h10408000;
      38922: inst = 32'hc405219;
      38923: inst = 32'h8220000;
      38924: inst = 32'h10408000;
      38925: inst = 32'hc40521a;
      38926: inst = 32'h8220000;
      38927: inst = 32'h10408000;
      38928: inst = 32'hc40521b;
      38929: inst = 32'h8220000;
      38930: inst = 32'h10408000;
      38931: inst = 32'hc40521c;
      38932: inst = 32'h8220000;
      38933: inst = 32'h10408000;
      38934: inst = 32'hc40521d;
      38935: inst = 32'h8220000;
      38936: inst = 32'h10408000;
      38937: inst = 32'hc40521e;
      38938: inst = 32'h8220000;
      38939: inst = 32'h10408000;
      38940: inst = 32'hc40521f;
      38941: inst = 32'h8220000;
      38942: inst = 32'h10408000;
      38943: inst = 32'hc405220;
      38944: inst = 32'h8220000;
      38945: inst = 32'h10408000;
      38946: inst = 32'hc405221;
      38947: inst = 32'h8220000;
      38948: inst = 32'h10408000;
      38949: inst = 32'hc405222;
      38950: inst = 32'h8220000;
      38951: inst = 32'h10408000;
      38952: inst = 32'hc405223;
      38953: inst = 32'h8220000;
      38954: inst = 32'h10408000;
      38955: inst = 32'hc405224;
      38956: inst = 32'h8220000;
      38957: inst = 32'h10408000;
      38958: inst = 32'hc405225;
      38959: inst = 32'h8220000;
      38960: inst = 32'h10408000;
      38961: inst = 32'hc405226;
      38962: inst = 32'h8220000;
      38963: inst = 32'h10408000;
      38964: inst = 32'hc405227;
      38965: inst = 32'h8220000;
      38966: inst = 32'h10408000;
      38967: inst = 32'hc405228;
      38968: inst = 32'h8220000;
      38969: inst = 32'h10408000;
      38970: inst = 32'hc405229;
      38971: inst = 32'h8220000;
      38972: inst = 32'h10408000;
      38973: inst = 32'hc40522a;
      38974: inst = 32'h8220000;
      38975: inst = 32'h10408000;
      38976: inst = 32'hc40522b;
      38977: inst = 32'h8220000;
      38978: inst = 32'h10408000;
      38979: inst = 32'hc40522c;
      38980: inst = 32'h8220000;
      38981: inst = 32'h10408000;
      38982: inst = 32'hc40522d;
      38983: inst = 32'h8220000;
      38984: inst = 32'h10408000;
      38985: inst = 32'hc40522e;
      38986: inst = 32'h8220000;
      38987: inst = 32'h10408000;
      38988: inst = 32'hc40522f;
      38989: inst = 32'h8220000;
      38990: inst = 32'h10408000;
      38991: inst = 32'hc405230;
      38992: inst = 32'h8220000;
      38993: inst = 32'h10408000;
      38994: inst = 32'hc405231;
      38995: inst = 32'h8220000;
      38996: inst = 32'h10408000;
      38997: inst = 32'hc405232;
      38998: inst = 32'h8220000;
      38999: inst = 32'h10408000;
      39000: inst = 32'hc405233;
      39001: inst = 32'h8220000;
      39002: inst = 32'h10408000;
      39003: inst = 32'hc405234;
      39004: inst = 32'h8220000;
      39005: inst = 32'h10408000;
      39006: inst = 32'hc405235;
      39007: inst = 32'h8220000;
      39008: inst = 32'h10408000;
      39009: inst = 32'hc405236;
      39010: inst = 32'h8220000;
      39011: inst = 32'h10408000;
      39012: inst = 32'hc405237;
      39013: inst = 32'h8220000;
      39014: inst = 32'h10408000;
      39015: inst = 32'hc405238;
      39016: inst = 32'h8220000;
      39017: inst = 32'h10408000;
      39018: inst = 32'hc405239;
      39019: inst = 32'h8220000;
      39020: inst = 32'h10408000;
      39021: inst = 32'hc40523a;
      39022: inst = 32'h8220000;
      39023: inst = 32'h10408000;
      39024: inst = 32'hc40523b;
      39025: inst = 32'h8220000;
      39026: inst = 32'h10408000;
      39027: inst = 32'hc40523c;
      39028: inst = 32'h8220000;
      39029: inst = 32'h10408000;
      39030: inst = 32'hc405243;
      39031: inst = 32'h8220000;
      39032: inst = 32'h10408000;
      39033: inst = 32'hc405244;
      39034: inst = 32'h8220000;
      39035: inst = 32'h10408000;
      39036: inst = 32'hc405245;
      39037: inst = 32'h8220000;
      39038: inst = 32'h10408000;
      39039: inst = 32'hc405246;
      39040: inst = 32'h8220000;
      39041: inst = 32'h10408000;
      39042: inst = 32'hc405247;
      39043: inst = 32'h8220000;
      39044: inst = 32'h10408000;
      39045: inst = 32'hc405248;
      39046: inst = 32'h8220000;
      39047: inst = 32'h10408000;
      39048: inst = 32'hc405249;
      39049: inst = 32'h8220000;
      39050: inst = 32'h10408000;
      39051: inst = 32'hc40524a;
      39052: inst = 32'h8220000;
      39053: inst = 32'h10408000;
      39054: inst = 32'hc40524b;
      39055: inst = 32'h8220000;
      39056: inst = 32'h10408000;
      39057: inst = 32'hc40524c;
      39058: inst = 32'h8220000;
      39059: inst = 32'h10408000;
      39060: inst = 32'hc40524d;
      39061: inst = 32'h8220000;
      39062: inst = 32'h10408000;
      39063: inst = 32'hc40524e;
      39064: inst = 32'h8220000;
      39065: inst = 32'h10408000;
      39066: inst = 32'hc40524f;
      39067: inst = 32'h8220000;
      39068: inst = 32'h10408000;
      39069: inst = 32'hc405250;
      39070: inst = 32'h8220000;
      39071: inst = 32'h10408000;
      39072: inst = 32'hc405251;
      39073: inst = 32'h8220000;
      39074: inst = 32'h10408000;
      39075: inst = 32'hc405252;
      39076: inst = 32'h8220000;
      39077: inst = 32'h10408000;
      39078: inst = 32'hc405253;
      39079: inst = 32'h8220000;
      39080: inst = 32'h10408000;
      39081: inst = 32'hc405254;
      39082: inst = 32'h8220000;
      39083: inst = 32'h10408000;
      39084: inst = 32'hc405255;
      39085: inst = 32'h8220000;
      39086: inst = 32'h10408000;
      39087: inst = 32'hc405259;
      39088: inst = 32'h8220000;
      39089: inst = 32'h10408000;
      39090: inst = 32'hc40525a;
      39091: inst = 32'h8220000;
      39092: inst = 32'h10408000;
      39093: inst = 32'hc40525b;
      39094: inst = 32'h8220000;
      39095: inst = 32'h10408000;
      39096: inst = 32'hc40525c;
      39097: inst = 32'h8220000;
      39098: inst = 32'h10408000;
      39099: inst = 32'hc40525d;
      39100: inst = 32'h8220000;
      39101: inst = 32'h10408000;
      39102: inst = 32'hc40525e;
      39103: inst = 32'h8220000;
      39104: inst = 32'h10408000;
      39105: inst = 32'hc40525f;
      39106: inst = 32'h8220000;
      39107: inst = 32'h10408000;
      39108: inst = 32'hc405260;
      39109: inst = 32'h8220000;
      39110: inst = 32'h10408000;
      39111: inst = 32'hc405261;
      39112: inst = 32'h8220000;
      39113: inst = 32'h10408000;
      39114: inst = 32'hc405262;
      39115: inst = 32'h8220000;
      39116: inst = 32'h10408000;
      39117: inst = 32'hc405263;
      39118: inst = 32'h8220000;
      39119: inst = 32'h10408000;
      39120: inst = 32'hc405264;
      39121: inst = 32'h8220000;
      39122: inst = 32'h10408000;
      39123: inst = 32'hc405265;
      39124: inst = 32'h8220000;
      39125: inst = 32'h10408000;
      39126: inst = 32'hc405266;
      39127: inst = 32'h8220000;
      39128: inst = 32'h10408000;
      39129: inst = 32'hc405267;
      39130: inst = 32'h8220000;
      39131: inst = 32'h10408000;
      39132: inst = 32'hc405268;
      39133: inst = 32'h8220000;
      39134: inst = 32'h10408000;
      39135: inst = 32'hc405269;
      39136: inst = 32'h8220000;
      39137: inst = 32'h10408000;
      39138: inst = 32'hc40526a;
      39139: inst = 32'h8220000;
      39140: inst = 32'h10408000;
      39141: inst = 32'hc40526b;
      39142: inst = 32'h8220000;
      39143: inst = 32'h10408000;
      39144: inst = 32'hc40526c;
      39145: inst = 32'h8220000;
      39146: inst = 32'h10408000;
      39147: inst = 32'hc40526d;
      39148: inst = 32'h8220000;
      39149: inst = 32'h10408000;
      39150: inst = 32'hc40526e;
      39151: inst = 32'h8220000;
      39152: inst = 32'h10408000;
      39153: inst = 32'hc40526f;
      39154: inst = 32'h8220000;
      39155: inst = 32'h10408000;
      39156: inst = 32'hc405270;
      39157: inst = 32'h8220000;
      39158: inst = 32'h10408000;
      39159: inst = 32'hc405271;
      39160: inst = 32'h8220000;
      39161: inst = 32'h10408000;
      39162: inst = 32'hc405272;
      39163: inst = 32'h8220000;
      39164: inst = 32'h10408000;
      39165: inst = 32'hc405273;
      39166: inst = 32'h8220000;
      39167: inst = 32'h10408000;
      39168: inst = 32'hc405274;
      39169: inst = 32'h8220000;
      39170: inst = 32'h10408000;
      39171: inst = 32'hc405275;
      39172: inst = 32'h8220000;
      39173: inst = 32'h10408000;
      39174: inst = 32'hc405276;
      39175: inst = 32'h8220000;
      39176: inst = 32'h10408000;
      39177: inst = 32'hc405277;
      39178: inst = 32'h8220000;
      39179: inst = 32'h10408000;
      39180: inst = 32'hc405278;
      39181: inst = 32'h8220000;
      39182: inst = 32'h10408000;
      39183: inst = 32'hc405279;
      39184: inst = 32'h8220000;
      39185: inst = 32'h10408000;
      39186: inst = 32'hc40527a;
      39187: inst = 32'h8220000;
      39188: inst = 32'h10408000;
      39189: inst = 32'hc40527b;
      39190: inst = 32'h8220000;
      39191: inst = 32'h10408000;
      39192: inst = 32'hc40527c;
      39193: inst = 32'h8220000;
      39194: inst = 32'h10408000;
      39195: inst = 32'hc40527d;
      39196: inst = 32'h8220000;
      39197: inst = 32'h10408000;
      39198: inst = 32'hc40527e;
      39199: inst = 32'h8220000;
      39200: inst = 32'h10408000;
      39201: inst = 32'hc40527f;
      39202: inst = 32'h8220000;
      39203: inst = 32'h10408000;
      39204: inst = 32'hc405280;
      39205: inst = 32'h8220000;
      39206: inst = 32'h10408000;
      39207: inst = 32'hc405281;
      39208: inst = 32'h8220000;
      39209: inst = 32'h10408000;
      39210: inst = 32'hc405282;
      39211: inst = 32'h8220000;
      39212: inst = 32'h10408000;
      39213: inst = 32'hc405283;
      39214: inst = 32'h8220000;
      39215: inst = 32'h10408000;
      39216: inst = 32'hc405284;
      39217: inst = 32'h8220000;
      39218: inst = 32'h10408000;
      39219: inst = 32'hc405285;
      39220: inst = 32'h8220000;
      39221: inst = 32'h10408000;
      39222: inst = 32'hc405286;
      39223: inst = 32'h8220000;
      39224: inst = 32'h10408000;
      39225: inst = 32'hc405287;
      39226: inst = 32'h8220000;
      39227: inst = 32'h10408000;
      39228: inst = 32'hc405288;
      39229: inst = 32'h8220000;
      39230: inst = 32'h10408000;
      39231: inst = 32'hc405289;
      39232: inst = 32'h8220000;
      39233: inst = 32'h10408000;
      39234: inst = 32'hc40528a;
      39235: inst = 32'h8220000;
      39236: inst = 32'h10408000;
      39237: inst = 32'hc40528b;
      39238: inst = 32'h8220000;
      39239: inst = 32'h10408000;
      39240: inst = 32'hc40528c;
      39241: inst = 32'h8220000;
      39242: inst = 32'h10408000;
      39243: inst = 32'hc40528d;
      39244: inst = 32'h8220000;
      39245: inst = 32'h10408000;
      39246: inst = 32'hc40528e;
      39247: inst = 32'h8220000;
      39248: inst = 32'h10408000;
      39249: inst = 32'hc40528f;
      39250: inst = 32'h8220000;
      39251: inst = 32'h10408000;
      39252: inst = 32'hc405290;
      39253: inst = 32'h8220000;
      39254: inst = 32'h10408000;
      39255: inst = 32'hc405291;
      39256: inst = 32'h8220000;
      39257: inst = 32'h10408000;
      39258: inst = 32'hc405292;
      39259: inst = 32'h8220000;
      39260: inst = 32'h10408000;
      39261: inst = 32'hc405293;
      39262: inst = 32'h8220000;
      39263: inst = 32'h10408000;
      39264: inst = 32'hc405294;
      39265: inst = 32'h8220000;
      39266: inst = 32'h10408000;
      39267: inst = 32'hc405295;
      39268: inst = 32'h8220000;
      39269: inst = 32'h10408000;
      39270: inst = 32'hc405296;
      39271: inst = 32'h8220000;
      39272: inst = 32'h10408000;
      39273: inst = 32'hc405297;
      39274: inst = 32'h8220000;
      39275: inst = 32'h10408000;
      39276: inst = 32'hc405298;
      39277: inst = 32'h8220000;
      39278: inst = 32'h10408000;
      39279: inst = 32'hc405299;
      39280: inst = 32'h8220000;
      39281: inst = 32'h10408000;
      39282: inst = 32'hc40529a;
      39283: inst = 32'h8220000;
      39284: inst = 32'h10408000;
      39285: inst = 32'hc40529b;
      39286: inst = 32'h8220000;
      39287: inst = 32'h10408000;
      39288: inst = 32'hc40529c;
      39289: inst = 32'h8220000;
      39290: inst = 32'h10408000;
      39291: inst = 32'hc4052a3;
      39292: inst = 32'h8220000;
      39293: inst = 32'h10408000;
      39294: inst = 32'hc4052a4;
      39295: inst = 32'h8220000;
      39296: inst = 32'h10408000;
      39297: inst = 32'hc4052a5;
      39298: inst = 32'h8220000;
      39299: inst = 32'h10408000;
      39300: inst = 32'hc4052a6;
      39301: inst = 32'h8220000;
      39302: inst = 32'h10408000;
      39303: inst = 32'hc4052a7;
      39304: inst = 32'h8220000;
      39305: inst = 32'h10408000;
      39306: inst = 32'hc4052a8;
      39307: inst = 32'h8220000;
      39308: inst = 32'h10408000;
      39309: inst = 32'hc4052a9;
      39310: inst = 32'h8220000;
      39311: inst = 32'h10408000;
      39312: inst = 32'hc4052aa;
      39313: inst = 32'h8220000;
      39314: inst = 32'h10408000;
      39315: inst = 32'hc4052ab;
      39316: inst = 32'h8220000;
      39317: inst = 32'h10408000;
      39318: inst = 32'hc4052ac;
      39319: inst = 32'h8220000;
      39320: inst = 32'h10408000;
      39321: inst = 32'hc4052ad;
      39322: inst = 32'h8220000;
      39323: inst = 32'h10408000;
      39324: inst = 32'hc4052ae;
      39325: inst = 32'h8220000;
      39326: inst = 32'h10408000;
      39327: inst = 32'hc4052af;
      39328: inst = 32'h8220000;
      39329: inst = 32'h10408000;
      39330: inst = 32'hc4052b0;
      39331: inst = 32'h8220000;
      39332: inst = 32'h10408000;
      39333: inst = 32'hc4052b1;
      39334: inst = 32'h8220000;
      39335: inst = 32'h10408000;
      39336: inst = 32'hc4052b2;
      39337: inst = 32'h8220000;
      39338: inst = 32'h10408000;
      39339: inst = 32'hc4052b3;
      39340: inst = 32'h8220000;
      39341: inst = 32'h10408000;
      39342: inst = 32'hc4052b4;
      39343: inst = 32'h8220000;
      39344: inst = 32'h10408000;
      39345: inst = 32'hc4052b5;
      39346: inst = 32'h8220000;
      39347: inst = 32'h10408000;
      39348: inst = 32'hc4052b9;
      39349: inst = 32'h8220000;
      39350: inst = 32'h10408000;
      39351: inst = 32'hc4052ba;
      39352: inst = 32'h8220000;
      39353: inst = 32'h10408000;
      39354: inst = 32'hc4052bb;
      39355: inst = 32'h8220000;
      39356: inst = 32'h10408000;
      39357: inst = 32'hc4052bc;
      39358: inst = 32'h8220000;
      39359: inst = 32'h10408000;
      39360: inst = 32'hc4052bd;
      39361: inst = 32'h8220000;
      39362: inst = 32'h10408000;
      39363: inst = 32'hc4052be;
      39364: inst = 32'h8220000;
      39365: inst = 32'h10408000;
      39366: inst = 32'hc4052bf;
      39367: inst = 32'h8220000;
      39368: inst = 32'h10408000;
      39369: inst = 32'hc4052c0;
      39370: inst = 32'h8220000;
      39371: inst = 32'h10408000;
      39372: inst = 32'hc4052c1;
      39373: inst = 32'h8220000;
      39374: inst = 32'h10408000;
      39375: inst = 32'hc4052c2;
      39376: inst = 32'h8220000;
      39377: inst = 32'h10408000;
      39378: inst = 32'hc4052c3;
      39379: inst = 32'h8220000;
      39380: inst = 32'h10408000;
      39381: inst = 32'hc4052c4;
      39382: inst = 32'h8220000;
      39383: inst = 32'h10408000;
      39384: inst = 32'hc4052c5;
      39385: inst = 32'h8220000;
      39386: inst = 32'h10408000;
      39387: inst = 32'hc4052c6;
      39388: inst = 32'h8220000;
      39389: inst = 32'h10408000;
      39390: inst = 32'hc4052c7;
      39391: inst = 32'h8220000;
      39392: inst = 32'h10408000;
      39393: inst = 32'hc4052c8;
      39394: inst = 32'h8220000;
      39395: inst = 32'h10408000;
      39396: inst = 32'hc4052c9;
      39397: inst = 32'h8220000;
      39398: inst = 32'h10408000;
      39399: inst = 32'hc4052ca;
      39400: inst = 32'h8220000;
      39401: inst = 32'h10408000;
      39402: inst = 32'hc4052cb;
      39403: inst = 32'h8220000;
      39404: inst = 32'h10408000;
      39405: inst = 32'hc4052cc;
      39406: inst = 32'h8220000;
      39407: inst = 32'h10408000;
      39408: inst = 32'hc4052cd;
      39409: inst = 32'h8220000;
      39410: inst = 32'h10408000;
      39411: inst = 32'hc4052ce;
      39412: inst = 32'h8220000;
      39413: inst = 32'h10408000;
      39414: inst = 32'hc4052cf;
      39415: inst = 32'h8220000;
      39416: inst = 32'h10408000;
      39417: inst = 32'hc4052d0;
      39418: inst = 32'h8220000;
      39419: inst = 32'h10408000;
      39420: inst = 32'hc4052d1;
      39421: inst = 32'h8220000;
      39422: inst = 32'h10408000;
      39423: inst = 32'hc4052d2;
      39424: inst = 32'h8220000;
      39425: inst = 32'h10408000;
      39426: inst = 32'hc4052d3;
      39427: inst = 32'h8220000;
      39428: inst = 32'h10408000;
      39429: inst = 32'hc4052d4;
      39430: inst = 32'h8220000;
      39431: inst = 32'h10408000;
      39432: inst = 32'hc4052d5;
      39433: inst = 32'h8220000;
      39434: inst = 32'h10408000;
      39435: inst = 32'hc4052d6;
      39436: inst = 32'h8220000;
      39437: inst = 32'h10408000;
      39438: inst = 32'hc4052d7;
      39439: inst = 32'h8220000;
      39440: inst = 32'h10408000;
      39441: inst = 32'hc4052d8;
      39442: inst = 32'h8220000;
      39443: inst = 32'h10408000;
      39444: inst = 32'hc4052d9;
      39445: inst = 32'h8220000;
      39446: inst = 32'h10408000;
      39447: inst = 32'hc4052da;
      39448: inst = 32'h8220000;
      39449: inst = 32'h10408000;
      39450: inst = 32'hc4052db;
      39451: inst = 32'h8220000;
      39452: inst = 32'h10408000;
      39453: inst = 32'hc4052dc;
      39454: inst = 32'h8220000;
      39455: inst = 32'h10408000;
      39456: inst = 32'hc4052dd;
      39457: inst = 32'h8220000;
      39458: inst = 32'h10408000;
      39459: inst = 32'hc4052de;
      39460: inst = 32'h8220000;
      39461: inst = 32'h10408000;
      39462: inst = 32'hc4052df;
      39463: inst = 32'h8220000;
      39464: inst = 32'h10408000;
      39465: inst = 32'hc4052e0;
      39466: inst = 32'h8220000;
      39467: inst = 32'h10408000;
      39468: inst = 32'hc4052e1;
      39469: inst = 32'h8220000;
      39470: inst = 32'h10408000;
      39471: inst = 32'hc4052e2;
      39472: inst = 32'h8220000;
      39473: inst = 32'h10408000;
      39474: inst = 32'hc4052e3;
      39475: inst = 32'h8220000;
      39476: inst = 32'h10408000;
      39477: inst = 32'hc4052e4;
      39478: inst = 32'h8220000;
      39479: inst = 32'h10408000;
      39480: inst = 32'hc4052e5;
      39481: inst = 32'h8220000;
      39482: inst = 32'h10408000;
      39483: inst = 32'hc4052e6;
      39484: inst = 32'h8220000;
      39485: inst = 32'h10408000;
      39486: inst = 32'hc4052e7;
      39487: inst = 32'h8220000;
      39488: inst = 32'h10408000;
      39489: inst = 32'hc4052e8;
      39490: inst = 32'h8220000;
      39491: inst = 32'h10408000;
      39492: inst = 32'hc4052e9;
      39493: inst = 32'h8220000;
      39494: inst = 32'h10408000;
      39495: inst = 32'hc4052ea;
      39496: inst = 32'h8220000;
      39497: inst = 32'h10408000;
      39498: inst = 32'hc4052eb;
      39499: inst = 32'h8220000;
      39500: inst = 32'h10408000;
      39501: inst = 32'hc4052ec;
      39502: inst = 32'h8220000;
      39503: inst = 32'h10408000;
      39504: inst = 32'hc4052ed;
      39505: inst = 32'h8220000;
      39506: inst = 32'h10408000;
      39507: inst = 32'hc4052ee;
      39508: inst = 32'h8220000;
      39509: inst = 32'h10408000;
      39510: inst = 32'hc4052ef;
      39511: inst = 32'h8220000;
      39512: inst = 32'h10408000;
      39513: inst = 32'hc4052f0;
      39514: inst = 32'h8220000;
      39515: inst = 32'h10408000;
      39516: inst = 32'hc4052f1;
      39517: inst = 32'h8220000;
      39518: inst = 32'h10408000;
      39519: inst = 32'hc4052f2;
      39520: inst = 32'h8220000;
      39521: inst = 32'h10408000;
      39522: inst = 32'hc4052f3;
      39523: inst = 32'h8220000;
      39524: inst = 32'h10408000;
      39525: inst = 32'hc4052f4;
      39526: inst = 32'h8220000;
      39527: inst = 32'h10408000;
      39528: inst = 32'hc4052f5;
      39529: inst = 32'h8220000;
      39530: inst = 32'h10408000;
      39531: inst = 32'hc4052f6;
      39532: inst = 32'h8220000;
      39533: inst = 32'h10408000;
      39534: inst = 32'hc4052f7;
      39535: inst = 32'h8220000;
      39536: inst = 32'h10408000;
      39537: inst = 32'hc4052f8;
      39538: inst = 32'h8220000;
      39539: inst = 32'h10408000;
      39540: inst = 32'hc4052f9;
      39541: inst = 32'h8220000;
      39542: inst = 32'h10408000;
      39543: inst = 32'hc4052fa;
      39544: inst = 32'h8220000;
      39545: inst = 32'h10408000;
      39546: inst = 32'hc4052fb;
      39547: inst = 32'h8220000;
      39548: inst = 32'h10408000;
      39549: inst = 32'hc4052fc;
      39550: inst = 32'h8220000;
      39551: inst = 32'h10408000;
      39552: inst = 32'hc405303;
      39553: inst = 32'h8220000;
      39554: inst = 32'h10408000;
      39555: inst = 32'hc405304;
      39556: inst = 32'h8220000;
      39557: inst = 32'h10408000;
      39558: inst = 32'hc405305;
      39559: inst = 32'h8220000;
      39560: inst = 32'h10408000;
      39561: inst = 32'hc405306;
      39562: inst = 32'h8220000;
      39563: inst = 32'h10408000;
      39564: inst = 32'hc405307;
      39565: inst = 32'h8220000;
      39566: inst = 32'h10408000;
      39567: inst = 32'hc405308;
      39568: inst = 32'h8220000;
      39569: inst = 32'h10408000;
      39570: inst = 32'hc405309;
      39571: inst = 32'h8220000;
      39572: inst = 32'h10408000;
      39573: inst = 32'hc40530a;
      39574: inst = 32'h8220000;
      39575: inst = 32'h10408000;
      39576: inst = 32'hc40530b;
      39577: inst = 32'h8220000;
      39578: inst = 32'h10408000;
      39579: inst = 32'hc40530c;
      39580: inst = 32'h8220000;
      39581: inst = 32'h10408000;
      39582: inst = 32'hc40530d;
      39583: inst = 32'h8220000;
      39584: inst = 32'h10408000;
      39585: inst = 32'hc40530e;
      39586: inst = 32'h8220000;
      39587: inst = 32'h10408000;
      39588: inst = 32'hc40530f;
      39589: inst = 32'h8220000;
      39590: inst = 32'h10408000;
      39591: inst = 32'hc405310;
      39592: inst = 32'h8220000;
      39593: inst = 32'h10408000;
      39594: inst = 32'hc405311;
      39595: inst = 32'h8220000;
      39596: inst = 32'h10408000;
      39597: inst = 32'hc405312;
      39598: inst = 32'h8220000;
      39599: inst = 32'h10408000;
      39600: inst = 32'hc405313;
      39601: inst = 32'h8220000;
      39602: inst = 32'h10408000;
      39603: inst = 32'hc405314;
      39604: inst = 32'h8220000;
      39605: inst = 32'h10408000;
      39606: inst = 32'hc405315;
      39607: inst = 32'h8220000;
      39608: inst = 32'h10408000;
      39609: inst = 32'hc405319;
      39610: inst = 32'h8220000;
      39611: inst = 32'h10408000;
      39612: inst = 32'hc40531a;
      39613: inst = 32'h8220000;
      39614: inst = 32'h10408000;
      39615: inst = 32'hc40531b;
      39616: inst = 32'h8220000;
      39617: inst = 32'h10408000;
      39618: inst = 32'hc40531c;
      39619: inst = 32'h8220000;
      39620: inst = 32'h10408000;
      39621: inst = 32'hc40531d;
      39622: inst = 32'h8220000;
      39623: inst = 32'h10408000;
      39624: inst = 32'hc40531e;
      39625: inst = 32'h8220000;
      39626: inst = 32'h10408000;
      39627: inst = 32'hc40531f;
      39628: inst = 32'h8220000;
      39629: inst = 32'h10408000;
      39630: inst = 32'hc405320;
      39631: inst = 32'h8220000;
      39632: inst = 32'h10408000;
      39633: inst = 32'hc405321;
      39634: inst = 32'h8220000;
      39635: inst = 32'h10408000;
      39636: inst = 32'hc405322;
      39637: inst = 32'h8220000;
      39638: inst = 32'h10408000;
      39639: inst = 32'hc405323;
      39640: inst = 32'h8220000;
      39641: inst = 32'h10408000;
      39642: inst = 32'hc405324;
      39643: inst = 32'h8220000;
      39644: inst = 32'h10408000;
      39645: inst = 32'hc405325;
      39646: inst = 32'h8220000;
      39647: inst = 32'h10408000;
      39648: inst = 32'hc405326;
      39649: inst = 32'h8220000;
      39650: inst = 32'h10408000;
      39651: inst = 32'hc405327;
      39652: inst = 32'h8220000;
      39653: inst = 32'h10408000;
      39654: inst = 32'hc405328;
      39655: inst = 32'h8220000;
      39656: inst = 32'h10408000;
      39657: inst = 32'hc405329;
      39658: inst = 32'h8220000;
      39659: inst = 32'h10408000;
      39660: inst = 32'hc40532a;
      39661: inst = 32'h8220000;
      39662: inst = 32'h10408000;
      39663: inst = 32'hc40532b;
      39664: inst = 32'h8220000;
      39665: inst = 32'h10408000;
      39666: inst = 32'hc40532c;
      39667: inst = 32'h8220000;
      39668: inst = 32'h10408000;
      39669: inst = 32'hc40532d;
      39670: inst = 32'h8220000;
      39671: inst = 32'h10408000;
      39672: inst = 32'hc40532e;
      39673: inst = 32'h8220000;
      39674: inst = 32'h10408000;
      39675: inst = 32'hc40532f;
      39676: inst = 32'h8220000;
      39677: inst = 32'h10408000;
      39678: inst = 32'hc405330;
      39679: inst = 32'h8220000;
      39680: inst = 32'h10408000;
      39681: inst = 32'hc405331;
      39682: inst = 32'h8220000;
      39683: inst = 32'h10408000;
      39684: inst = 32'hc405332;
      39685: inst = 32'h8220000;
      39686: inst = 32'h10408000;
      39687: inst = 32'hc405333;
      39688: inst = 32'h8220000;
      39689: inst = 32'h10408000;
      39690: inst = 32'hc405334;
      39691: inst = 32'h8220000;
      39692: inst = 32'h10408000;
      39693: inst = 32'hc405335;
      39694: inst = 32'h8220000;
      39695: inst = 32'h10408000;
      39696: inst = 32'hc405336;
      39697: inst = 32'h8220000;
      39698: inst = 32'h10408000;
      39699: inst = 32'hc405337;
      39700: inst = 32'h8220000;
      39701: inst = 32'h10408000;
      39702: inst = 32'hc405338;
      39703: inst = 32'h8220000;
      39704: inst = 32'h10408000;
      39705: inst = 32'hc405339;
      39706: inst = 32'h8220000;
      39707: inst = 32'h10408000;
      39708: inst = 32'hc40533a;
      39709: inst = 32'h8220000;
      39710: inst = 32'h10408000;
      39711: inst = 32'hc40533b;
      39712: inst = 32'h8220000;
      39713: inst = 32'h10408000;
      39714: inst = 32'hc40533c;
      39715: inst = 32'h8220000;
      39716: inst = 32'h10408000;
      39717: inst = 32'hc40533d;
      39718: inst = 32'h8220000;
      39719: inst = 32'h10408000;
      39720: inst = 32'hc40533e;
      39721: inst = 32'h8220000;
      39722: inst = 32'h10408000;
      39723: inst = 32'hc40533f;
      39724: inst = 32'h8220000;
      39725: inst = 32'h10408000;
      39726: inst = 32'hc405340;
      39727: inst = 32'h8220000;
      39728: inst = 32'h10408000;
      39729: inst = 32'hc405341;
      39730: inst = 32'h8220000;
      39731: inst = 32'h10408000;
      39732: inst = 32'hc405342;
      39733: inst = 32'h8220000;
      39734: inst = 32'h10408000;
      39735: inst = 32'hc405343;
      39736: inst = 32'h8220000;
      39737: inst = 32'h10408000;
      39738: inst = 32'hc405344;
      39739: inst = 32'h8220000;
      39740: inst = 32'h10408000;
      39741: inst = 32'hc405345;
      39742: inst = 32'h8220000;
      39743: inst = 32'h10408000;
      39744: inst = 32'hc405346;
      39745: inst = 32'h8220000;
      39746: inst = 32'h10408000;
      39747: inst = 32'hc405347;
      39748: inst = 32'h8220000;
      39749: inst = 32'h10408000;
      39750: inst = 32'hc405348;
      39751: inst = 32'h8220000;
      39752: inst = 32'h10408000;
      39753: inst = 32'hc405349;
      39754: inst = 32'h8220000;
      39755: inst = 32'h10408000;
      39756: inst = 32'hc40534a;
      39757: inst = 32'h8220000;
      39758: inst = 32'h10408000;
      39759: inst = 32'hc40534b;
      39760: inst = 32'h8220000;
      39761: inst = 32'h10408000;
      39762: inst = 32'hc40534c;
      39763: inst = 32'h8220000;
      39764: inst = 32'h10408000;
      39765: inst = 32'hc40534d;
      39766: inst = 32'h8220000;
      39767: inst = 32'h10408000;
      39768: inst = 32'hc40534e;
      39769: inst = 32'h8220000;
      39770: inst = 32'h10408000;
      39771: inst = 32'hc40534f;
      39772: inst = 32'h8220000;
      39773: inst = 32'h10408000;
      39774: inst = 32'hc405350;
      39775: inst = 32'h8220000;
      39776: inst = 32'h10408000;
      39777: inst = 32'hc405351;
      39778: inst = 32'h8220000;
      39779: inst = 32'h10408000;
      39780: inst = 32'hc40535c;
      39781: inst = 32'h8220000;
      39782: inst = 32'h10408000;
      39783: inst = 32'hc405363;
      39784: inst = 32'h8220000;
      39785: inst = 32'h10408000;
      39786: inst = 32'hc405364;
      39787: inst = 32'h8220000;
      39788: inst = 32'h10408000;
      39789: inst = 32'hc405365;
      39790: inst = 32'h8220000;
      39791: inst = 32'h10408000;
      39792: inst = 32'hc405366;
      39793: inst = 32'h8220000;
      39794: inst = 32'h10408000;
      39795: inst = 32'hc405367;
      39796: inst = 32'h8220000;
      39797: inst = 32'h10408000;
      39798: inst = 32'hc405368;
      39799: inst = 32'h8220000;
      39800: inst = 32'h10408000;
      39801: inst = 32'hc405369;
      39802: inst = 32'h8220000;
      39803: inst = 32'h10408000;
      39804: inst = 32'hc40536a;
      39805: inst = 32'h8220000;
      39806: inst = 32'h10408000;
      39807: inst = 32'hc40536b;
      39808: inst = 32'h8220000;
      39809: inst = 32'h10408000;
      39810: inst = 32'hc40536c;
      39811: inst = 32'h8220000;
      39812: inst = 32'h10408000;
      39813: inst = 32'hc40536d;
      39814: inst = 32'h8220000;
      39815: inst = 32'h10408000;
      39816: inst = 32'hc40536e;
      39817: inst = 32'h8220000;
      39818: inst = 32'h10408000;
      39819: inst = 32'hc40536f;
      39820: inst = 32'h8220000;
      39821: inst = 32'h10408000;
      39822: inst = 32'hc405370;
      39823: inst = 32'h8220000;
      39824: inst = 32'h10408000;
      39825: inst = 32'hc405371;
      39826: inst = 32'h8220000;
      39827: inst = 32'h10408000;
      39828: inst = 32'hc405372;
      39829: inst = 32'h8220000;
      39830: inst = 32'h10408000;
      39831: inst = 32'hc405373;
      39832: inst = 32'h8220000;
      39833: inst = 32'h10408000;
      39834: inst = 32'hc405374;
      39835: inst = 32'h8220000;
      39836: inst = 32'h10408000;
      39837: inst = 32'hc405375;
      39838: inst = 32'h8220000;
      39839: inst = 32'h10408000;
      39840: inst = 32'hc405379;
      39841: inst = 32'h8220000;
      39842: inst = 32'h10408000;
      39843: inst = 32'hc40537a;
      39844: inst = 32'h8220000;
      39845: inst = 32'h10408000;
      39846: inst = 32'hc40537b;
      39847: inst = 32'h8220000;
      39848: inst = 32'h10408000;
      39849: inst = 32'hc40537c;
      39850: inst = 32'h8220000;
      39851: inst = 32'h10408000;
      39852: inst = 32'hc40537d;
      39853: inst = 32'h8220000;
      39854: inst = 32'h10408000;
      39855: inst = 32'hc40537e;
      39856: inst = 32'h8220000;
      39857: inst = 32'h10408000;
      39858: inst = 32'hc40537f;
      39859: inst = 32'h8220000;
      39860: inst = 32'h10408000;
      39861: inst = 32'hc405380;
      39862: inst = 32'h8220000;
      39863: inst = 32'h10408000;
      39864: inst = 32'hc405381;
      39865: inst = 32'h8220000;
      39866: inst = 32'h10408000;
      39867: inst = 32'hc405382;
      39868: inst = 32'h8220000;
      39869: inst = 32'h10408000;
      39870: inst = 32'hc405383;
      39871: inst = 32'h8220000;
      39872: inst = 32'h10408000;
      39873: inst = 32'hc405384;
      39874: inst = 32'h8220000;
      39875: inst = 32'h10408000;
      39876: inst = 32'hc405385;
      39877: inst = 32'h8220000;
      39878: inst = 32'h10408000;
      39879: inst = 32'hc405386;
      39880: inst = 32'h8220000;
      39881: inst = 32'h10408000;
      39882: inst = 32'hc405387;
      39883: inst = 32'h8220000;
      39884: inst = 32'h10408000;
      39885: inst = 32'hc405388;
      39886: inst = 32'h8220000;
      39887: inst = 32'h10408000;
      39888: inst = 32'hc405389;
      39889: inst = 32'h8220000;
      39890: inst = 32'h10408000;
      39891: inst = 32'hc40538a;
      39892: inst = 32'h8220000;
      39893: inst = 32'h10408000;
      39894: inst = 32'hc40538b;
      39895: inst = 32'h8220000;
      39896: inst = 32'h10408000;
      39897: inst = 32'hc40538c;
      39898: inst = 32'h8220000;
      39899: inst = 32'h10408000;
      39900: inst = 32'hc40538d;
      39901: inst = 32'h8220000;
      39902: inst = 32'h10408000;
      39903: inst = 32'hc40538e;
      39904: inst = 32'h8220000;
      39905: inst = 32'h10408000;
      39906: inst = 32'hc40538f;
      39907: inst = 32'h8220000;
      39908: inst = 32'h10408000;
      39909: inst = 32'hc405390;
      39910: inst = 32'h8220000;
      39911: inst = 32'h10408000;
      39912: inst = 32'hc405391;
      39913: inst = 32'h8220000;
      39914: inst = 32'h10408000;
      39915: inst = 32'hc405392;
      39916: inst = 32'h8220000;
      39917: inst = 32'h10408000;
      39918: inst = 32'hc405393;
      39919: inst = 32'h8220000;
      39920: inst = 32'h10408000;
      39921: inst = 32'hc405394;
      39922: inst = 32'h8220000;
      39923: inst = 32'h10408000;
      39924: inst = 32'hc405395;
      39925: inst = 32'h8220000;
      39926: inst = 32'h10408000;
      39927: inst = 32'hc405396;
      39928: inst = 32'h8220000;
      39929: inst = 32'h10408000;
      39930: inst = 32'hc405397;
      39931: inst = 32'h8220000;
      39932: inst = 32'h10408000;
      39933: inst = 32'hc405398;
      39934: inst = 32'h8220000;
      39935: inst = 32'h10408000;
      39936: inst = 32'hc405399;
      39937: inst = 32'h8220000;
      39938: inst = 32'h10408000;
      39939: inst = 32'hc40539a;
      39940: inst = 32'h8220000;
      39941: inst = 32'h10408000;
      39942: inst = 32'hc40539b;
      39943: inst = 32'h8220000;
      39944: inst = 32'h10408000;
      39945: inst = 32'hc40539c;
      39946: inst = 32'h8220000;
      39947: inst = 32'h10408000;
      39948: inst = 32'hc40539d;
      39949: inst = 32'h8220000;
      39950: inst = 32'h10408000;
      39951: inst = 32'hc40539e;
      39952: inst = 32'h8220000;
      39953: inst = 32'h10408000;
      39954: inst = 32'hc40539f;
      39955: inst = 32'h8220000;
      39956: inst = 32'h10408000;
      39957: inst = 32'hc4053a0;
      39958: inst = 32'h8220000;
      39959: inst = 32'h10408000;
      39960: inst = 32'hc4053a1;
      39961: inst = 32'h8220000;
      39962: inst = 32'h10408000;
      39963: inst = 32'hc4053a2;
      39964: inst = 32'h8220000;
      39965: inst = 32'h10408000;
      39966: inst = 32'hc4053a3;
      39967: inst = 32'h8220000;
      39968: inst = 32'h10408000;
      39969: inst = 32'hc4053a4;
      39970: inst = 32'h8220000;
      39971: inst = 32'h10408000;
      39972: inst = 32'hc4053a5;
      39973: inst = 32'h8220000;
      39974: inst = 32'h10408000;
      39975: inst = 32'hc4053a6;
      39976: inst = 32'h8220000;
      39977: inst = 32'h10408000;
      39978: inst = 32'hc4053a7;
      39979: inst = 32'h8220000;
      39980: inst = 32'h10408000;
      39981: inst = 32'hc4053a8;
      39982: inst = 32'h8220000;
      39983: inst = 32'h10408000;
      39984: inst = 32'hc4053a9;
      39985: inst = 32'h8220000;
      39986: inst = 32'h10408000;
      39987: inst = 32'hc4053aa;
      39988: inst = 32'h8220000;
      39989: inst = 32'h10408000;
      39990: inst = 32'hc4053ab;
      39991: inst = 32'h8220000;
      39992: inst = 32'h10408000;
      39993: inst = 32'hc4053ac;
      39994: inst = 32'h8220000;
      39995: inst = 32'h10408000;
      39996: inst = 32'hc4053ad;
      39997: inst = 32'h8220000;
      39998: inst = 32'h10408000;
      39999: inst = 32'hc4053ae;
      40000: inst = 32'h8220000;
      40001: inst = 32'h10408000;
      40002: inst = 32'hc4053af;
      40003: inst = 32'h8220000;
      40004: inst = 32'h10408000;
      40005: inst = 32'hc4053b0;
      40006: inst = 32'h8220000;
      40007: inst = 32'h10408000;
      40008: inst = 32'hc4053b1;
      40009: inst = 32'h8220000;
      40010: inst = 32'h10408000;
      40011: inst = 32'hc4053bc;
      40012: inst = 32'h8220000;
      40013: inst = 32'h10408000;
      40014: inst = 32'hc4053c3;
      40015: inst = 32'h8220000;
      40016: inst = 32'h10408000;
      40017: inst = 32'hc4053c4;
      40018: inst = 32'h8220000;
      40019: inst = 32'h10408000;
      40020: inst = 32'hc4053c5;
      40021: inst = 32'h8220000;
      40022: inst = 32'h10408000;
      40023: inst = 32'hc4053c6;
      40024: inst = 32'h8220000;
      40025: inst = 32'h10408000;
      40026: inst = 32'hc4053c7;
      40027: inst = 32'h8220000;
      40028: inst = 32'h10408000;
      40029: inst = 32'hc4053cf;
      40030: inst = 32'h8220000;
      40031: inst = 32'h10408000;
      40032: inst = 32'hc4053d0;
      40033: inst = 32'h8220000;
      40034: inst = 32'h10408000;
      40035: inst = 32'hc4053d1;
      40036: inst = 32'h8220000;
      40037: inst = 32'h10408000;
      40038: inst = 32'hc4053d2;
      40039: inst = 32'h8220000;
      40040: inst = 32'h10408000;
      40041: inst = 32'hc4053d3;
      40042: inst = 32'h8220000;
      40043: inst = 32'h10408000;
      40044: inst = 32'hc4053d4;
      40045: inst = 32'h8220000;
      40046: inst = 32'h10408000;
      40047: inst = 32'hc4053d5;
      40048: inst = 32'h8220000;
      40049: inst = 32'h10408000;
      40050: inst = 32'hc4053d9;
      40051: inst = 32'h8220000;
      40052: inst = 32'h10408000;
      40053: inst = 32'hc4053da;
      40054: inst = 32'h8220000;
      40055: inst = 32'h10408000;
      40056: inst = 32'hc4053db;
      40057: inst = 32'h8220000;
      40058: inst = 32'h10408000;
      40059: inst = 32'hc4053dc;
      40060: inst = 32'h8220000;
      40061: inst = 32'h10408000;
      40062: inst = 32'hc4053dd;
      40063: inst = 32'h8220000;
      40064: inst = 32'h10408000;
      40065: inst = 32'hc4053de;
      40066: inst = 32'h8220000;
      40067: inst = 32'h10408000;
      40068: inst = 32'hc4053df;
      40069: inst = 32'h8220000;
      40070: inst = 32'h10408000;
      40071: inst = 32'hc4053e0;
      40072: inst = 32'h8220000;
      40073: inst = 32'h10408000;
      40074: inst = 32'hc4053e1;
      40075: inst = 32'h8220000;
      40076: inst = 32'h10408000;
      40077: inst = 32'hc4053e2;
      40078: inst = 32'h8220000;
      40079: inst = 32'h10408000;
      40080: inst = 32'hc4053e3;
      40081: inst = 32'h8220000;
      40082: inst = 32'h10408000;
      40083: inst = 32'hc4053e4;
      40084: inst = 32'h8220000;
      40085: inst = 32'h10408000;
      40086: inst = 32'hc4053e5;
      40087: inst = 32'h8220000;
      40088: inst = 32'h10408000;
      40089: inst = 32'hc4053e6;
      40090: inst = 32'h8220000;
      40091: inst = 32'h10408000;
      40092: inst = 32'hc4053e7;
      40093: inst = 32'h8220000;
      40094: inst = 32'h10408000;
      40095: inst = 32'hc4053e8;
      40096: inst = 32'h8220000;
      40097: inst = 32'h10408000;
      40098: inst = 32'hc4053e9;
      40099: inst = 32'h8220000;
      40100: inst = 32'h10408000;
      40101: inst = 32'hc4053ea;
      40102: inst = 32'h8220000;
      40103: inst = 32'h10408000;
      40104: inst = 32'hc4053eb;
      40105: inst = 32'h8220000;
      40106: inst = 32'h10408000;
      40107: inst = 32'hc4053ec;
      40108: inst = 32'h8220000;
      40109: inst = 32'h10408000;
      40110: inst = 32'hc4053ed;
      40111: inst = 32'h8220000;
      40112: inst = 32'h10408000;
      40113: inst = 32'hc4053ee;
      40114: inst = 32'h8220000;
      40115: inst = 32'h10408000;
      40116: inst = 32'hc4053ef;
      40117: inst = 32'h8220000;
      40118: inst = 32'h10408000;
      40119: inst = 32'hc4053f0;
      40120: inst = 32'h8220000;
      40121: inst = 32'h10408000;
      40122: inst = 32'hc4053f1;
      40123: inst = 32'h8220000;
      40124: inst = 32'h10408000;
      40125: inst = 32'hc4053f2;
      40126: inst = 32'h8220000;
      40127: inst = 32'h10408000;
      40128: inst = 32'hc4053f3;
      40129: inst = 32'h8220000;
      40130: inst = 32'h10408000;
      40131: inst = 32'hc4053f4;
      40132: inst = 32'h8220000;
      40133: inst = 32'h10408000;
      40134: inst = 32'hc4053f5;
      40135: inst = 32'h8220000;
      40136: inst = 32'h10408000;
      40137: inst = 32'hc4053f6;
      40138: inst = 32'h8220000;
      40139: inst = 32'h10408000;
      40140: inst = 32'hc4053f7;
      40141: inst = 32'h8220000;
      40142: inst = 32'h10408000;
      40143: inst = 32'hc4053f8;
      40144: inst = 32'h8220000;
      40145: inst = 32'h10408000;
      40146: inst = 32'hc4053f9;
      40147: inst = 32'h8220000;
      40148: inst = 32'h10408000;
      40149: inst = 32'hc4053fa;
      40150: inst = 32'h8220000;
      40151: inst = 32'h10408000;
      40152: inst = 32'hc4053fb;
      40153: inst = 32'h8220000;
      40154: inst = 32'h10408000;
      40155: inst = 32'hc4053fc;
      40156: inst = 32'h8220000;
      40157: inst = 32'h10408000;
      40158: inst = 32'hc4053fd;
      40159: inst = 32'h8220000;
      40160: inst = 32'h10408000;
      40161: inst = 32'hc4053fe;
      40162: inst = 32'h8220000;
      40163: inst = 32'h10408000;
      40164: inst = 32'hc4053ff;
      40165: inst = 32'h8220000;
      40166: inst = 32'h10408000;
      40167: inst = 32'hc405400;
      40168: inst = 32'h8220000;
      40169: inst = 32'h10408000;
      40170: inst = 32'hc405401;
      40171: inst = 32'h8220000;
      40172: inst = 32'h10408000;
      40173: inst = 32'hc405402;
      40174: inst = 32'h8220000;
      40175: inst = 32'h10408000;
      40176: inst = 32'hc405403;
      40177: inst = 32'h8220000;
      40178: inst = 32'h10408000;
      40179: inst = 32'hc405404;
      40180: inst = 32'h8220000;
      40181: inst = 32'h10408000;
      40182: inst = 32'hc405405;
      40183: inst = 32'h8220000;
      40184: inst = 32'h10408000;
      40185: inst = 32'hc405406;
      40186: inst = 32'h8220000;
      40187: inst = 32'h10408000;
      40188: inst = 32'hc405407;
      40189: inst = 32'h8220000;
      40190: inst = 32'h10408000;
      40191: inst = 32'hc405408;
      40192: inst = 32'h8220000;
      40193: inst = 32'h10408000;
      40194: inst = 32'hc405409;
      40195: inst = 32'h8220000;
      40196: inst = 32'h10408000;
      40197: inst = 32'hc40540a;
      40198: inst = 32'h8220000;
      40199: inst = 32'h10408000;
      40200: inst = 32'hc40540b;
      40201: inst = 32'h8220000;
      40202: inst = 32'h10408000;
      40203: inst = 32'hc40540c;
      40204: inst = 32'h8220000;
      40205: inst = 32'h10408000;
      40206: inst = 32'hc40540d;
      40207: inst = 32'h8220000;
      40208: inst = 32'h10408000;
      40209: inst = 32'hc40540e;
      40210: inst = 32'h8220000;
      40211: inst = 32'h10408000;
      40212: inst = 32'hc40540f;
      40213: inst = 32'h8220000;
      40214: inst = 32'h10408000;
      40215: inst = 32'hc405410;
      40216: inst = 32'h8220000;
      40217: inst = 32'h10408000;
      40218: inst = 32'hc405411;
      40219: inst = 32'h8220000;
      40220: inst = 32'h10408000;
      40221: inst = 32'hc40541c;
      40222: inst = 32'h8220000;
      40223: inst = 32'h10408000;
      40224: inst = 32'hc405423;
      40225: inst = 32'h8220000;
      40226: inst = 32'h10408000;
      40227: inst = 32'hc405424;
      40228: inst = 32'h8220000;
      40229: inst = 32'h10408000;
      40230: inst = 32'hc405425;
      40231: inst = 32'h8220000;
      40232: inst = 32'h10408000;
      40233: inst = 32'hc405426;
      40234: inst = 32'h8220000;
      40235: inst = 32'h10408000;
      40236: inst = 32'hc405430;
      40237: inst = 32'h8220000;
      40238: inst = 32'h10408000;
      40239: inst = 32'hc405431;
      40240: inst = 32'h8220000;
      40241: inst = 32'h10408000;
      40242: inst = 32'hc405432;
      40243: inst = 32'h8220000;
      40244: inst = 32'h10408000;
      40245: inst = 32'hc405433;
      40246: inst = 32'h8220000;
      40247: inst = 32'h10408000;
      40248: inst = 32'hc405434;
      40249: inst = 32'h8220000;
      40250: inst = 32'h10408000;
      40251: inst = 32'hc405435;
      40252: inst = 32'h8220000;
      40253: inst = 32'h10408000;
      40254: inst = 32'hc40544a;
      40255: inst = 32'h8220000;
      40256: inst = 32'h10408000;
      40257: inst = 32'hc40544b;
      40258: inst = 32'h8220000;
      40259: inst = 32'h10408000;
      40260: inst = 32'hc40544c;
      40261: inst = 32'h8220000;
      40262: inst = 32'h10408000;
      40263: inst = 32'hc40544d;
      40264: inst = 32'h8220000;
      40265: inst = 32'h10408000;
      40266: inst = 32'hc40544e;
      40267: inst = 32'h8220000;
      40268: inst = 32'h10408000;
      40269: inst = 32'hc40544f;
      40270: inst = 32'h8220000;
      40271: inst = 32'h10408000;
      40272: inst = 32'hc405450;
      40273: inst = 32'h8220000;
      40274: inst = 32'h10408000;
      40275: inst = 32'hc405451;
      40276: inst = 32'h8220000;
      40277: inst = 32'h10408000;
      40278: inst = 32'hc405452;
      40279: inst = 32'h8220000;
      40280: inst = 32'h10408000;
      40281: inst = 32'hc405453;
      40282: inst = 32'h8220000;
      40283: inst = 32'h10408000;
      40284: inst = 32'hc405454;
      40285: inst = 32'h8220000;
      40286: inst = 32'h10408000;
      40287: inst = 32'hc405455;
      40288: inst = 32'h8220000;
      40289: inst = 32'h10408000;
      40290: inst = 32'hc405456;
      40291: inst = 32'h8220000;
      40292: inst = 32'h10408000;
      40293: inst = 32'hc405457;
      40294: inst = 32'h8220000;
      40295: inst = 32'h10408000;
      40296: inst = 32'hc405458;
      40297: inst = 32'h8220000;
      40298: inst = 32'h10408000;
      40299: inst = 32'hc405459;
      40300: inst = 32'h8220000;
      40301: inst = 32'h10408000;
      40302: inst = 32'hc40545a;
      40303: inst = 32'h8220000;
      40304: inst = 32'h10408000;
      40305: inst = 32'hc40545b;
      40306: inst = 32'h8220000;
      40307: inst = 32'h10408000;
      40308: inst = 32'hc40545c;
      40309: inst = 32'h8220000;
      40310: inst = 32'h10408000;
      40311: inst = 32'hc40545d;
      40312: inst = 32'h8220000;
      40313: inst = 32'h10408000;
      40314: inst = 32'hc40545e;
      40315: inst = 32'h8220000;
      40316: inst = 32'h10408000;
      40317: inst = 32'hc40545f;
      40318: inst = 32'h8220000;
      40319: inst = 32'h10408000;
      40320: inst = 32'hc405460;
      40321: inst = 32'h8220000;
      40322: inst = 32'h10408000;
      40323: inst = 32'hc405461;
      40324: inst = 32'h8220000;
      40325: inst = 32'h10408000;
      40326: inst = 32'hc405462;
      40327: inst = 32'h8220000;
      40328: inst = 32'h10408000;
      40329: inst = 32'hc405463;
      40330: inst = 32'h8220000;
      40331: inst = 32'h10408000;
      40332: inst = 32'hc405464;
      40333: inst = 32'h8220000;
      40334: inst = 32'h10408000;
      40335: inst = 32'hc405465;
      40336: inst = 32'h8220000;
      40337: inst = 32'h10408000;
      40338: inst = 32'hc405466;
      40339: inst = 32'h8220000;
      40340: inst = 32'h10408000;
      40341: inst = 32'hc405467;
      40342: inst = 32'h8220000;
      40343: inst = 32'h10408000;
      40344: inst = 32'hc405468;
      40345: inst = 32'h8220000;
      40346: inst = 32'h10408000;
      40347: inst = 32'hc405469;
      40348: inst = 32'h8220000;
      40349: inst = 32'h10408000;
      40350: inst = 32'hc40546a;
      40351: inst = 32'h8220000;
      40352: inst = 32'h10408000;
      40353: inst = 32'hc40546b;
      40354: inst = 32'h8220000;
      40355: inst = 32'h10408000;
      40356: inst = 32'hc40546c;
      40357: inst = 32'h8220000;
      40358: inst = 32'h10408000;
      40359: inst = 32'hc40546d;
      40360: inst = 32'h8220000;
      40361: inst = 32'h10408000;
      40362: inst = 32'hc40546e;
      40363: inst = 32'h8220000;
      40364: inst = 32'h10408000;
      40365: inst = 32'hc40546f;
      40366: inst = 32'h8220000;
      40367: inst = 32'h10408000;
      40368: inst = 32'hc405470;
      40369: inst = 32'h8220000;
      40370: inst = 32'h10408000;
      40371: inst = 32'hc405471;
      40372: inst = 32'h8220000;
      40373: inst = 32'h10408000;
      40374: inst = 32'hc40547c;
      40375: inst = 32'h8220000;
      40376: inst = 32'h10408000;
      40377: inst = 32'hc405483;
      40378: inst = 32'h8220000;
      40379: inst = 32'h10408000;
      40380: inst = 32'hc405484;
      40381: inst = 32'h8220000;
      40382: inst = 32'h10408000;
      40383: inst = 32'hc405485;
      40384: inst = 32'h8220000;
      40385: inst = 32'h10408000;
      40386: inst = 32'hc405486;
      40387: inst = 32'h8220000;
      40388: inst = 32'h10408000;
      40389: inst = 32'hc405490;
      40390: inst = 32'h8220000;
      40391: inst = 32'h10408000;
      40392: inst = 32'hc405491;
      40393: inst = 32'h8220000;
      40394: inst = 32'h10408000;
      40395: inst = 32'hc405492;
      40396: inst = 32'h8220000;
      40397: inst = 32'h10408000;
      40398: inst = 32'hc405493;
      40399: inst = 32'h8220000;
      40400: inst = 32'h10408000;
      40401: inst = 32'hc405494;
      40402: inst = 32'h8220000;
      40403: inst = 32'h10408000;
      40404: inst = 32'hc405495;
      40405: inst = 32'h8220000;
      40406: inst = 32'h10408000;
      40407: inst = 32'hc4054aa;
      40408: inst = 32'h8220000;
      40409: inst = 32'h10408000;
      40410: inst = 32'hc4054ab;
      40411: inst = 32'h8220000;
      40412: inst = 32'h10408000;
      40413: inst = 32'hc4054ac;
      40414: inst = 32'h8220000;
      40415: inst = 32'h10408000;
      40416: inst = 32'hc4054ad;
      40417: inst = 32'h8220000;
      40418: inst = 32'h10408000;
      40419: inst = 32'hc4054ae;
      40420: inst = 32'h8220000;
      40421: inst = 32'h10408000;
      40422: inst = 32'hc4054af;
      40423: inst = 32'h8220000;
      40424: inst = 32'h10408000;
      40425: inst = 32'hc4054b0;
      40426: inst = 32'h8220000;
      40427: inst = 32'h10408000;
      40428: inst = 32'hc4054b1;
      40429: inst = 32'h8220000;
      40430: inst = 32'h10408000;
      40431: inst = 32'hc4054b2;
      40432: inst = 32'h8220000;
      40433: inst = 32'h10408000;
      40434: inst = 32'hc4054b3;
      40435: inst = 32'h8220000;
      40436: inst = 32'h10408000;
      40437: inst = 32'hc4054b4;
      40438: inst = 32'h8220000;
      40439: inst = 32'h10408000;
      40440: inst = 32'hc4054b5;
      40441: inst = 32'h8220000;
      40442: inst = 32'h10408000;
      40443: inst = 32'hc4054b6;
      40444: inst = 32'h8220000;
      40445: inst = 32'h10408000;
      40446: inst = 32'hc4054b7;
      40447: inst = 32'h8220000;
      40448: inst = 32'h10408000;
      40449: inst = 32'hc4054b8;
      40450: inst = 32'h8220000;
      40451: inst = 32'h10408000;
      40452: inst = 32'hc4054b9;
      40453: inst = 32'h8220000;
      40454: inst = 32'h10408000;
      40455: inst = 32'hc4054ba;
      40456: inst = 32'h8220000;
      40457: inst = 32'h10408000;
      40458: inst = 32'hc4054bb;
      40459: inst = 32'h8220000;
      40460: inst = 32'h10408000;
      40461: inst = 32'hc4054bc;
      40462: inst = 32'h8220000;
      40463: inst = 32'h10408000;
      40464: inst = 32'hc4054bd;
      40465: inst = 32'h8220000;
      40466: inst = 32'h10408000;
      40467: inst = 32'hc4054be;
      40468: inst = 32'h8220000;
      40469: inst = 32'h10408000;
      40470: inst = 32'hc4054bf;
      40471: inst = 32'h8220000;
      40472: inst = 32'h10408000;
      40473: inst = 32'hc4054c0;
      40474: inst = 32'h8220000;
      40475: inst = 32'h10408000;
      40476: inst = 32'hc4054c1;
      40477: inst = 32'h8220000;
      40478: inst = 32'h10408000;
      40479: inst = 32'hc4054c2;
      40480: inst = 32'h8220000;
      40481: inst = 32'h10408000;
      40482: inst = 32'hc4054c3;
      40483: inst = 32'h8220000;
      40484: inst = 32'h10408000;
      40485: inst = 32'hc4054c4;
      40486: inst = 32'h8220000;
      40487: inst = 32'h10408000;
      40488: inst = 32'hc4054c5;
      40489: inst = 32'h8220000;
      40490: inst = 32'h10408000;
      40491: inst = 32'hc4054c6;
      40492: inst = 32'h8220000;
      40493: inst = 32'h10408000;
      40494: inst = 32'hc4054c7;
      40495: inst = 32'h8220000;
      40496: inst = 32'h10408000;
      40497: inst = 32'hc4054c8;
      40498: inst = 32'h8220000;
      40499: inst = 32'h10408000;
      40500: inst = 32'hc4054c9;
      40501: inst = 32'h8220000;
      40502: inst = 32'h10408000;
      40503: inst = 32'hc4054ca;
      40504: inst = 32'h8220000;
      40505: inst = 32'h10408000;
      40506: inst = 32'hc4054cb;
      40507: inst = 32'h8220000;
      40508: inst = 32'h10408000;
      40509: inst = 32'hc4054cc;
      40510: inst = 32'h8220000;
      40511: inst = 32'h10408000;
      40512: inst = 32'hc4054cd;
      40513: inst = 32'h8220000;
      40514: inst = 32'h10408000;
      40515: inst = 32'hc4054ce;
      40516: inst = 32'h8220000;
      40517: inst = 32'h10408000;
      40518: inst = 32'hc4054cf;
      40519: inst = 32'h8220000;
      40520: inst = 32'h10408000;
      40521: inst = 32'hc4054d0;
      40522: inst = 32'h8220000;
      40523: inst = 32'h10408000;
      40524: inst = 32'hc4054d1;
      40525: inst = 32'h8220000;
      40526: inst = 32'h10408000;
      40527: inst = 32'hc4054dc;
      40528: inst = 32'h8220000;
      40529: inst = 32'h10408000;
      40530: inst = 32'hc4054e3;
      40531: inst = 32'h8220000;
      40532: inst = 32'h10408000;
      40533: inst = 32'hc4054e4;
      40534: inst = 32'h8220000;
      40535: inst = 32'h10408000;
      40536: inst = 32'hc4054e5;
      40537: inst = 32'h8220000;
      40538: inst = 32'h10408000;
      40539: inst = 32'hc4054e6;
      40540: inst = 32'h8220000;
      40541: inst = 32'h10408000;
      40542: inst = 32'hc4054f0;
      40543: inst = 32'h8220000;
      40544: inst = 32'h10408000;
      40545: inst = 32'hc4054f1;
      40546: inst = 32'h8220000;
      40547: inst = 32'h10408000;
      40548: inst = 32'hc4054f2;
      40549: inst = 32'h8220000;
      40550: inst = 32'h10408000;
      40551: inst = 32'hc4054f3;
      40552: inst = 32'h8220000;
      40553: inst = 32'h10408000;
      40554: inst = 32'hc4054f4;
      40555: inst = 32'h8220000;
      40556: inst = 32'h10408000;
      40557: inst = 32'hc4054f5;
      40558: inst = 32'h8220000;
      40559: inst = 32'h10408000;
      40560: inst = 32'hc40550a;
      40561: inst = 32'h8220000;
      40562: inst = 32'h10408000;
      40563: inst = 32'hc40550b;
      40564: inst = 32'h8220000;
      40565: inst = 32'h10408000;
      40566: inst = 32'hc40550c;
      40567: inst = 32'h8220000;
      40568: inst = 32'h10408000;
      40569: inst = 32'hc40550d;
      40570: inst = 32'h8220000;
      40571: inst = 32'h10408000;
      40572: inst = 32'hc40550e;
      40573: inst = 32'h8220000;
      40574: inst = 32'h10408000;
      40575: inst = 32'hc40550f;
      40576: inst = 32'h8220000;
      40577: inst = 32'h10408000;
      40578: inst = 32'hc405510;
      40579: inst = 32'h8220000;
      40580: inst = 32'h10408000;
      40581: inst = 32'hc405511;
      40582: inst = 32'h8220000;
      40583: inst = 32'h10408000;
      40584: inst = 32'hc405512;
      40585: inst = 32'h8220000;
      40586: inst = 32'h10408000;
      40587: inst = 32'hc405513;
      40588: inst = 32'h8220000;
      40589: inst = 32'h10408000;
      40590: inst = 32'hc405514;
      40591: inst = 32'h8220000;
      40592: inst = 32'h10408000;
      40593: inst = 32'hc405515;
      40594: inst = 32'h8220000;
      40595: inst = 32'h10408000;
      40596: inst = 32'hc405516;
      40597: inst = 32'h8220000;
      40598: inst = 32'h10408000;
      40599: inst = 32'hc405517;
      40600: inst = 32'h8220000;
      40601: inst = 32'h10408000;
      40602: inst = 32'hc405518;
      40603: inst = 32'h8220000;
      40604: inst = 32'h10408000;
      40605: inst = 32'hc405519;
      40606: inst = 32'h8220000;
      40607: inst = 32'h10408000;
      40608: inst = 32'hc40551a;
      40609: inst = 32'h8220000;
      40610: inst = 32'h10408000;
      40611: inst = 32'hc40551b;
      40612: inst = 32'h8220000;
      40613: inst = 32'h10408000;
      40614: inst = 32'hc40551c;
      40615: inst = 32'h8220000;
      40616: inst = 32'h10408000;
      40617: inst = 32'hc40551d;
      40618: inst = 32'h8220000;
      40619: inst = 32'h10408000;
      40620: inst = 32'hc40551e;
      40621: inst = 32'h8220000;
      40622: inst = 32'h10408000;
      40623: inst = 32'hc40551f;
      40624: inst = 32'h8220000;
      40625: inst = 32'h10408000;
      40626: inst = 32'hc405520;
      40627: inst = 32'h8220000;
      40628: inst = 32'h10408000;
      40629: inst = 32'hc405521;
      40630: inst = 32'h8220000;
      40631: inst = 32'h10408000;
      40632: inst = 32'hc405522;
      40633: inst = 32'h8220000;
      40634: inst = 32'h10408000;
      40635: inst = 32'hc405523;
      40636: inst = 32'h8220000;
      40637: inst = 32'h10408000;
      40638: inst = 32'hc405524;
      40639: inst = 32'h8220000;
      40640: inst = 32'h10408000;
      40641: inst = 32'hc405525;
      40642: inst = 32'h8220000;
      40643: inst = 32'h10408000;
      40644: inst = 32'hc405526;
      40645: inst = 32'h8220000;
      40646: inst = 32'h10408000;
      40647: inst = 32'hc405527;
      40648: inst = 32'h8220000;
      40649: inst = 32'h10408000;
      40650: inst = 32'hc405528;
      40651: inst = 32'h8220000;
      40652: inst = 32'h10408000;
      40653: inst = 32'hc405529;
      40654: inst = 32'h8220000;
      40655: inst = 32'h10408000;
      40656: inst = 32'hc40552a;
      40657: inst = 32'h8220000;
      40658: inst = 32'h10408000;
      40659: inst = 32'hc40552b;
      40660: inst = 32'h8220000;
      40661: inst = 32'h10408000;
      40662: inst = 32'hc40552c;
      40663: inst = 32'h8220000;
      40664: inst = 32'h10408000;
      40665: inst = 32'hc40552d;
      40666: inst = 32'h8220000;
      40667: inst = 32'h10408000;
      40668: inst = 32'hc40552e;
      40669: inst = 32'h8220000;
      40670: inst = 32'h10408000;
      40671: inst = 32'hc40552f;
      40672: inst = 32'h8220000;
      40673: inst = 32'h10408000;
      40674: inst = 32'hc405530;
      40675: inst = 32'h8220000;
      40676: inst = 32'h10408000;
      40677: inst = 32'hc405531;
      40678: inst = 32'h8220000;
      40679: inst = 32'h10408000;
      40680: inst = 32'hc40553c;
      40681: inst = 32'h8220000;
      40682: inst = 32'h10408000;
      40683: inst = 32'hc405543;
      40684: inst = 32'h8220000;
      40685: inst = 32'h10408000;
      40686: inst = 32'hc405544;
      40687: inst = 32'h8220000;
      40688: inst = 32'h10408000;
      40689: inst = 32'hc405545;
      40690: inst = 32'h8220000;
      40691: inst = 32'h10408000;
      40692: inst = 32'hc405546;
      40693: inst = 32'h8220000;
      40694: inst = 32'h10408000;
      40695: inst = 32'hc405550;
      40696: inst = 32'h8220000;
      40697: inst = 32'h10408000;
      40698: inst = 32'hc405551;
      40699: inst = 32'h8220000;
      40700: inst = 32'h10408000;
      40701: inst = 32'hc405552;
      40702: inst = 32'h8220000;
      40703: inst = 32'h10408000;
      40704: inst = 32'hc405553;
      40705: inst = 32'h8220000;
      40706: inst = 32'h10408000;
      40707: inst = 32'hc405554;
      40708: inst = 32'h8220000;
      40709: inst = 32'h10408000;
      40710: inst = 32'hc405555;
      40711: inst = 32'h8220000;
      40712: inst = 32'h10408000;
      40713: inst = 32'hc405559;
      40714: inst = 32'h8220000;
      40715: inst = 32'h10408000;
      40716: inst = 32'hc40555a;
      40717: inst = 32'h8220000;
      40718: inst = 32'h10408000;
      40719: inst = 32'hc40555b;
      40720: inst = 32'h8220000;
      40721: inst = 32'h10408000;
      40722: inst = 32'hc40555c;
      40723: inst = 32'h8220000;
      40724: inst = 32'h10408000;
      40725: inst = 32'hc40555d;
      40726: inst = 32'h8220000;
      40727: inst = 32'h10408000;
      40728: inst = 32'hc40555e;
      40729: inst = 32'h8220000;
      40730: inst = 32'h10408000;
      40731: inst = 32'hc40555f;
      40732: inst = 32'h8220000;
      40733: inst = 32'h10408000;
      40734: inst = 32'hc405560;
      40735: inst = 32'h8220000;
      40736: inst = 32'h10408000;
      40737: inst = 32'hc405561;
      40738: inst = 32'h8220000;
      40739: inst = 32'h10408000;
      40740: inst = 32'hc405562;
      40741: inst = 32'h8220000;
      40742: inst = 32'h10408000;
      40743: inst = 32'hc405563;
      40744: inst = 32'h8220000;
      40745: inst = 32'h10408000;
      40746: inst = 32'hc405564;
      40747: inst = 32'h8220000;
      40748: inst = 32'h10408000;
      40749: inst = 32'hc405565;
      40750: inst = 32'h8220000;
      40751: inst = 32'h10408000;
      40752: inst = 32'hc405566;
      40753: inst = 32'h8220000;
      40754: inst = 32'h10408000;
      40755: inst = 32'hc405567;
      40756: inst = 32'h8220000;
      40757: inst = 32'h10408000;
      40758: inst = 32'hc405568;
      40759: inst = 32'h8220000;
      40760: inst = 32'h10408000;
      40761: inst = 32'hc405569;
      40762: inst = 32'h8220000;
      40763: inst = 32'h10408000;
      40764: inst = 32'hc40556a;
      40765: inst = 32'h8220000;
      40766: inst = 32'h10408000;
      40767: inst = 32'hc40556b;
      40768: inst = 32'h8220000;
      40769: inst = 32'h10408000;
      40770: inst = 32'hc40556c;
      40771: inst = 32'h8220000;
      40772: inst = 32'h10408000;
      40773: inst = 32'hc40556d;
      40774: inst = 32'h8220000;
      40775: inst = 32'h10408000;
      40776: inst = 32'hc40556e;
      40777: inst = 32'h8220000;
      40778: inst = 32'h10408000;
      40779: inst = 32'hc40556f;
      40780: inst = 32'h8220000;
      40781: inst = 32'h10408000;
      40782: inst = 32'hc405570;
      40783: inst = 32'h8220000;
      40784: inst = 32'h10408000;
      40785: inst = 32'hc405571;
      40786: inst = 32'h8220000;
      40787: inst = 32'h10408000;
      40788: inst = 32'hc405572;
      40789: inst = 32'h8220000;
      40790: inst = 32'h10408000;
      40791: inst = 32'hc405573;
      40792: inst = 32'h8220000;
      40793: inst = 32'h10408000;
      40794: inst = 32'hc405574;
      40795: inst = 32'h8220000;
      40796: inst = 32'h10408000;
      40797: inst = 32'hc405575;
      40798: inst = 32'h8220000;
      40799: inst = 32'h10408000;
      40800: inst = 32'hc405576;
      40801: inst = 32'h8220000;
      40802: inst = 32'h10408000;
      40803: inst = 32'hc405577;
      40804: inst = 32'h8220000;
      40805: inst = 32'h10408000;
      40806: inst = 32'hc405578;
      40807: inst = 32'h8220000;
      40808: inst = 32'h10408000;
      40809: inst = 32'hc405579;
      40810: inst = 32'h8220000;
      40811: inst = 32'h10408000;
      40812: inst = 32'hc40557a;
      40813: inst = 32'h8220000;
      40814: inst = 32'h10408000;
      40815: inst = 32'hc40557b;
      40816: inst = 32'h8220000;
      40817: inst = 32'h10408000;
      40818: inst = 32'hc40557c;
      40819: inst = 32'h8220000;
      40820: inst = 32'h10408000;
      40821: inst = 32'hc40557d;
      40822: inst = 32'h8220000;
      40823: inst = 32'h10408000;
      40824: inst = 32'hc40557e;
      40825: inst = 32'h8220000;
      40826: inst = 32'h10408000;
      40827: inst = 32'hc40557f;
      40828: inst = 32'h8220000;
      40829: inst = 32'h10408000;
      40830: inst = 32'hc405580;
      40831: inst = 32'h8220000;
      40832: inst = 32'h10408000;
      40833: inst = 32'hc405581;
      40834: inst = 32'h8220000;
      40835: inst = 32'h10408000;
      40836: inst = 32'hc405582;
      40837: inst = 32'h8220000;
      40838: inst = 32'h10408000;
      40839: inst = 32'hc405583;
      40840: inst = 32'h8220000;
      40841: inst = 32'h10408000;
      40842: inst = 32'hc405584;
      40843: inst = 32'h8220000;
      40844: inst = 32'h10408000;
      40845: inst = 32'hc405585;
      40846: inst = 32'h8220000;
      40847: inst = 32'h10408000;
      40848: inst = 32'hc405586;
      40849: inst = 32'h8220000;
      40850: inst = 32'h10408000;
      40851: inst = 32'hc405587;
      40852: inst = 32'h8220000;
      40853: inst = 32'h10408000;
      40854: inst = 32'hc405588;
      40855: inst = 32'h8220000;
      40856: inst = 32'h10408000;
      40857: inst = 32'hc405589;
      40858: inst = 32'h8220000;
      40859: inst = 32'h10408000;
      40860: inst = 32'hc40558a;
      40861: inst = 32'h8220000;
      40862: inst = 32'h10408000;
      40863: inst = 32'hc40558b;
      40864: inst = 32'h8220000;
      40865: inst = 32'h10408000;
      40866: inst = 32'hc40558c;
      40867: inst = 32'h8220000;
      40868: inst = 32'h10408000;
      40869: inst = 32'hc40558d;
      40870: inst = 32'h8220000;
      40871: inst = 32'h10408000;
      40872: inst = 32'hc40558e;
      40873: inst = 32'h8220000;
      40874: inst = 32'h10408000;
      40875: inst = 32'hc40558f;
      40876: inst = 32'h8220000;
      40877: inst = 32'h10408000;
      40878: inst = 32'hc405590;
      40879: inst = 32'h8220000;
      40880: inst = 32'h10408000;
      40881: inst = 32'hc405591;
      40882: inst = 32'h8220000;
      40883: inst = 32'h10408000;
      40884: inst = 32'hc40559c;
      40885: inst = 32'h8220000;
      40886: inst = 32'h10408000;
      40887: inst = 32'hc4055a3;
      40888: inst = 32'h8220000;
      40889: inst = 32'h10408000;
      40890: inst = 32'hc4055a4;
      40891: inst = 32'h8220000;
      40892: inst = 32'h10408000;
      40893: inst = 32'hc4055a5;
      40894: inst = 32'h8220000;
      40895: inst = 32'h10408000;
      40896: inst = 32'hc4055a6;
      40897: inst = 32'h8220000;
      40898: inst = 32'h10408000;
      40899: inst = 32'hc4055b0;
      40900: inst = 32'h8220000;
      40901: inst = 32'h10408000;
      40902: inst = 32'hc4055b1;
      40903: inst = 32'h8220000;
      40904: inst = 32'h10408000;
      40905: inst = 32'hc4055b2;
      40906: inst = 32'h8220000;
      40907: inst = 32'h10408000;
      40908: inst = 32'hc4055b3;
      40909: inst = 32'h8220000;
      40910: inst = 32'h10408000;
      40911: inst = 32'hc4055b4;
      40912: inst = 32'h8220000;
      40913: inst = 32'h10408000;
      40914: inst = 32'hc4055b5;
      40915: inst = 32'h8220000;
      40916: inst = 32'h10408000;
      40917: inst = 32'hc4055b9;
      40918: inst = 32'h8220000;
      40919: inst = 32'h10408000;
      40920: inst = 32'hc4055ba;
      40921: inst = 32'h8220000;
      40922: inst = 32'h10408000;
      40923: inst = 32'hc4055bb;
      40924: inst = 32'h8220000;
      40925: inst = 32'h10408000;
      40926: inst = 32'hc4055bc;
      40927: inst = 32'h8220000;
      40928: inst = 32'h10408000;
      40929: inst = 32'hc4055bd;
      40930: inst = 32'h8220000;
      40931: inst = 32'h10408000;
      40932: inst = 32'hc4055be;
      40933: inst = 32'h8220000;
      40934: inst = 32'h10408000;
      40935: inst = 32'hc4055bf;
      40936: inst = 32'h8220000;
      40937: inst = 32'h10408000;
      40938: inst = 32'hc4055c0;
      40939: inst = 32'h8220000;
      40940: inst = 32'h10408000;
      40941: inst = 32'hc4055c1;
      40942: inst = 32'h8220000;
      40943: inst = 32'h10408000;
      40944: inst = 32'hc4055c2;
      40945: inst = 32'h8220000;
      40946: inst = 32'h10408000;
      40947: inst = 32'hc4055c3;
      40948: inst = 32'h8220000;
      40949: inst = 32'h10408000;
      40950: inst = 32'hc4055c4;
      40951: inst = 32'h8220000;
      40952: inst = 32'h10408000;
      40953: inst = 32'hc4055c5;
      40954: inst = 32'h8220000;
      40955: inst = 32'h10408000;
      40956: inst = 32'hc4055c6;
      40957: inst = 32'h8220000;
      40958: inst = 32'h10408000;
      40959: inst = 32'hc4055c7;
      40960: inst = 32'h8220000;
      40961: inst = 32'h10408000;
      40962: inst = 32'hc4055c8;
      40963: inst = 32'h8220000;
      40964: inst = 32'h10408000;
      40965: inst = 32'hc4055c9;
      40966: inst = 32'h8220000;
      40967: inst = 32'h10408000;
      40968: inst = 32'hc4055ca;
      40969: inst = 32'h8220000;
      40970: inst = 32'h10408000;
      40971: inst = 32'hc4055cb;
      40972: inst = 32'h8220000;
      40973: inst = 32'h10408000;
      40974: inst = 32'hc4055cc;
      40975: inst = 32'h8220000;
      40976: inst = 32'h10408000;
      40977: inst = 32'hc4055cd;
      40978: inst = 32'h8220000;
      40979: inst = 32'h10408000;
      40980: inst = 32'hc4055ce;
      40981: inst = 32'h8220000;
      40982: inst = 32'h10408000;
      40983: inst = 32'hc4055cf;
      40984: inst = 32'h8220000;
      40985: inst = 32'h10408000;
      40986: inst = 32'hc4055d0;
      40987: inst = 32'h8220000;
      40988: inst = 32'h10408000;
      40989: inst = 32'hc4055d1;
      40990: inst = 32'h8220000;
      40991: inst = 32'h10408000;
      40992: inst = 32'hc4055d2;
      40993: inst = 32'h8220000;
      40994: inst = 32'h10408000;
      40995: inst = 32'hc4055d3;
      40996: inst = 32'h8220000;
      40997: inst = 32'h10408000;
      40998: inst = 32'hc4055d4;
      40999: inst = 32'h8220000;
      41000: inst = 32'h10408000;
      41001: inst = 32'hc4055d5;
      41002: inst = 32'h8220000;
      41003: inst = 32'h10408000;
      41004: inst = 32'hc4055d6;
      41005: inst = 32'h8220000;
      41006: inst = 32'h10408000;
      41007: inst = 32'hc4055d7;
      41008: inst = 32'h8220000;
      41009: inst = 32'h10408000;
      41010: inst = 32'hc4055d8;
      41011: inst = 32'h8220000;
      41012: inst = 32'h10408000;
      41013: inst = 32'hc4055d9;
      41014: inst = 32'h8220000;
      41015: inst = 32'h10408000;
      41016: inst = 32'hc4055da;
      41017: inst = 32'h8220000;
      41018: inst = 32'h10408000;
      41019: inst = 32'hc4055db;
      41020: inst = 32'h8220000;
      41021: inst = 32'h10408000;
      41022: inst = 32'hc4055dc;
      41023: inst = 32'h8220000;
      41024: inst = 32'h10408000;
      41025: inst = 32'hc4055dd;
      41026: inst = 32'h8220000;
      41027: inst = 32'h10408000;
      41028: inst = 32'hc4055de;
      41029: inst = 32'h8220000;
      41030: inst = 32'h10408000;
      41031: inst = 32'hc4055df;
      41032: inst = 32'h8220000;
      41033: inst = 32'h10408000;
      41034: inst = 32'hc4055e0;
      41035: inst = 32'h8220000;
      41036: inst = 32'h10408000;
      41037: inst = 32'hc4055e1;
      41038: inst = 32'h8220000;
      41039: inst = 32'h10408000;
      41040: inst = 32'hc4055e2;
      41041: inst = 32'h8220000;
      41042: inst = 32'h10408000;
      41043: inst = 32'hc4055e3;
      41044: inst = 32'h8220000;
      41045: inst = 32'h10408000;
      41046: inst = 32'hc4055e4;
      41047: inst = 32'h8220000;
      41048: inst = 32'h10408000;
      41049: inst = 32'hc4055e5;
      41050: inst = 32'h8220000;
      41051: inst = 32'h10408000;
      41052: inst = 32'hc4055e6;
      41053: inst = 32'h8220000;
      41054: inst = 32'h10408000;
      41055: inst = 32'hc4055e7;
      41056: inst = 32'h8220000;
      41057: inst = 32'h10408000;
      41058: inst = 32'hc4055e8;
      41059: inst = 32'h8220000;
      41060: inst = 32'h10408000;
      41061: inst = 32'hc4055e9;
      41062: inst = 32'h8220000;
      41063: inst = 32'h10408000;
      41064: inst = 32'hc4055ea;
      41065: inst = 32'h8220000;
      41066: inst = 32'h10408000;
      41067: inst = 32'hc4055eb;
      41068: inst = 32'h8220000;
      41069: inst = 32'h10408000;
      41070: inst = 32'hc4055ec;
      41071: inst = 32'h8220000;
      41072: inst = 32'h10408000;
      41073: inst = 32'hc4055ed;
      41074: inst = 32'h8220000;
      41075: inst = 32'h10408000;
      41076: inst = 32'hc4055ee;
      41077: inst = 32'h8220000;
      41078: inst = 32'h10408000;
      41079: inst = 32'hc4055ef;
      41080: inst = 32'h8220000;
      41081: inst = 32'h10408000;
      41082: inst = 32'hc4055f0;
      41083: inst = 32'h8220000;
      41084: inst = 32'h10408000;
      41085: inst = 32'hc4055f1;
      41086: inst = 32'h8220000;
      41087: inst = 32'h10408000;
      41088: inst = 32'hc4055fc;
      41089: inst = 32'h8220000;
      41090: inst = 32'h10408000;
      41091: inst = 32'hc405603;
      41092: inst = 32'h8220000;
      41093: inst = 32'h10408000;
      41094: inst = 32'hc405604;
      41095: inst = 32'h8220000;
      41096: inst = 32'h10408000;
      41097: inst = 32'hc405605;
      41098: inst = 32'h8220000;
      41099: inst = 32'h10408000;
      41100: inst = 32'hc405606;
      41101: inst = 32'h8220000;
      41102: inst = 32'h10408000;
      41103: inst = 32'hc405613;
      41104: inst = 32'h8220000;
      41105: inst = 32'h10408000;
      41106: inst = 32'hc405614;
      41107: inst = 32'h8220000;
      41108: inst = 32'h10408000;
      41109: inst = 32'hc405615;
      41110: inst = 32'h8220000;
      41111: inst = 32'h10408000;
      41112: inst = 32'hc405619;
      41113: inst = 32'h8220000;
      41114: inst = 32'h10408000;
      41115: inst = 32'hc40561a;
      41116: inst = 32'h8220000;
      41117: inst = 32'h10408000;
      41118: inst = 32'hc40561b;
      41119: inst = 32'h8220000;
      41120: inst = 32'h10408000;
      41121: inst = 32'hc40561c;
      41122: inst = 32'h8220000;
      41123: inst = 32'h10408000;
      41124: inst = 32'hc40561d;
      41125: inst = 32'h8220000;
      41126: inst = 32'h10408000;
      41127: inst = 32'hc40561e;
      41128: inst = 32'h8220000;
      41129: inst = 32'h10408000;
      41130: inst = 32'hc40561f;
      41131: inst = 32'h8220000;
      41132: inst = 32'h10408000;
      41133: inst = 32'hc405620;
      41134: inst = 32'h8220000;
      41135: inst = 32'h10408000;
      41136: inst = 32'hc405621;
      41137: inst = 32'h8220000;
      41138: inst = 32'h10408000;
      41139: inst = 32'hc405622;
      41140: inst = 32'h8220000;
      41141: inst = 32'h10408000;
      41142: inst = 32'hc405623;
      41143: inst = 32'h8220000;
      41144: inst = 32'h10408000;
      41145: inst = 32'hc405624;
      41146: inst = 32'h8220000;
      41147: inst = 32'h10408000;
      41148: inst = 32'hc405625;
      41149: inst = 32'h8220000;
      41150: inst = 32'h10408000;
      41151: inst = 32'hc405626;
      41152: inst = 32'h8220000;
      41153: inst = 32'h10408000;
      41154: inst = 32'hc405627;
      41155: inst = 32'h8220000;
      41156: inst = 32'h10408000;
      41157: inst = 32'hc405628;
      41158: inst = 32'h8220000;
      41159: inst = 32'h10408000;
      41160: inst = 32'hc405629;
      41161: inst = 32'h8220000;
      41162: inst = 32'h10408000;
      41163: inst = 32'hc40562a;
      41164: inst = 32'h8220000;
      41165: inst = 32'h10408000;
      41166: inst = 32'hc40562b;
      41167: inst = 32'h8220000;
      41168: inst = 32'h10408000;
      41169: inst = 32'hc40562c;
      41170: inst = 32'h8220000;
      41171: inst = 32'h10408000;
      41172: inst = 32'hc40562d;
      41173: inst = 32'h8220000;
      41174: inst = 32'h10408000;
      41175: inst = 32'hc40562e;
      41176: inst = 32'h8220000;
      41177: inst = 32'h10408000;
      41178: inst = 32'hc40562f;
      41179: inst = 32'h8220000;
      41180: inst = 32'h10408000;
      41181: inst = 32'hc405630;
      41182: inst = 32'h8220000;
      41183: inst = 32'h10408000;
      41184: inst = 32'hc405631;
      41185: inst = 32'h8220000;
      41186: inst = 32'h10408000;
      41187: inst = 32'hc405632;
      41188: inst = 32'h8220000;
      41189: inst = 32'h10408000;
      41190: inst = 32'hc405633;
      41191: inst = 32'h8220000;
      41192: inst = 32'h10408000;
      41193: inst = 32'hc405634;
      41194: inst = 32'h8220000;
      41195: inst = 32'h10408000;
      41196: inst = 32'hc405635;
      41197: inst = 32'h8220000;
      41198: inst = 32'h10408000;
      41199: inst = 32'hc405636;
      41200: inst = 32'h8220000;
      41201: inst = 32'h10408000;
      41202: inst = 32'hc405637;
      41203: inst = 32'h8220000;
      41204: inst = 32'h10408000;
      41205: inst = 32'hc405638;
      41206: inst = 32'h8220000;
      41207: inst = 32'h10408000;
      41208: inst = 32'hc405639;
      41209: inst = 32'h8220000;
      41210: inst = 32'h10408000;
      41211: inst = 32'hc40563a;
      41212: inst = 32'h8220000;
      41213: inst = 32'h10408000;
      41214: inst = 32'hc40563b;
      41215: inst = 32'h8220000;
      41216: inst = 32'h10408000;
      41217: inst = 32'hc40563c;
      41218: inst = 32'h8220000;
      41219: inst = 32'h10408000;
      41220: inst = 32'hc40563d;
      41221: inst = 32'h8220000;
      41222: inst = 32'h10408000;
      41223: inst = 32'hc40563e;
      41224: inst = 32'h8220000;
      41225: inst = 32'h10408000;
      41226: inst = 32'hc40563f;
      41227: inst = 32'h8220000;
      41228: inst = 32'h10408000;
      41229: inst = 32'hc405640;
      41230: inst = 32'h8220000;
      41231: inst = 32'h10408000;
      41232: inst = 32'hc405641;
      41233: inst = 32'h8220000;
      41234: inst = 32'h10408000;
      41235: inst = 32'hc405642;
      41236: inst = 32'h8220000;
      41237: inst = 32'h10408000;
      41238: inst = 32'hc405643;
      41239: inst = 32'h8220000;
      41240: inst = 32'h10408000;
      41241: inst = 32'hc405644;
      41242: inst = 32'h8220000;
      41243: inst = 32'h10408000;
      41244: inst = 32'hc405645;
      41245: inst = 32'h8220000;
      41246: inst = 32'h10408000;
      41247: inst = 32'hc405646;
      41248: inst = 32'h8220000;
      41249: inst = 32'h10408000;
      41250: inst = 32'hc405647;
      41251: inst = 32'h8220000;
      41252: inst = 32'h10408000;
      41253: inst = 32'hc405648;
      41254: inst = 32'h8220000;
      41255: inst = 32'h10408000;
      41256: inst = 32'hc405649;
      41257: inst = 32'h8220000;
      41258: inst = 32'h10408000;
      41259: inst = 32'hc40564a;
      41260: inst = 32'h8220000;
      41261: inst = 32'h10408000;
      41262: inst = 32'hc40564b;
      41263: inst = 32'h8220000;
      41264: inst = 32'h10408000;
      41265: inst = 32'hc40564c;
      41266: inst = 32'h8220000;
      41267: inst = 32'h10408000;
      41268: inst = 32'hc40564d;
      41269: inst = 32'h8220000;
      41270: inst = 32'h10408000;
      41271: inst = 32'hc40564e;
      41272: inst = 32'h8220000;
      41273: inst = 32'h10408000;
      41274: inst = 32'hc40564f;
      41275: inst = 32'h8220000;
      41276: inst = 32'h10408000;
      41277: inst = 32'hc405650;
      41278: inst = 32'h8220000;
      41279: inst = 32'h10408000;
      41280: inst = 32'hc405651;
      41281: inst = 32'h8220000;
      41282: inst = 32'h10408000;
      41283: inst = 32'hc40565c;
      41284: inst = 32'h8220000;
      41285: inst = 32'h10408000;
      41286: inst = 32'hc405663;
      41287: inst = 32'h8220000;
      41288: inst = 32'h10408000;
      41289: inst = 32'hc405664;
      41290: inst = 32'h8220000;
      41291: inst = 32'h10408000;
      41292: inst = 32'hc405665;
      41293: inst = 32'h8220000;
      41294: inst = 32'h10408000;
      41295: inst = 32'hc405666;
      41296: inst = 32'h8220000;
      41297: inst = 32'h10408000;
      41298: inst = 32'hc405667;
      41299: inst = 32'h8220000;
      41300: inst = 32'h10408000;
      41301: inst = 32'hc405674;
      41302: inst = 32'h8220000;
      41303: inst = 32'h10408000;
      41304: inst = 32'hc405675;
      41305: inst = 32'h8220000;
      41306: inst = 32'h10408000;
      41307: inst = 32'hc405679;
      41308: inst = 32'h8220000;
      41309: inst = 32'h10408000;
      41310: inst = 32'hc40567a;
      41311: inst = 32'h8220000;
      41312: inst = 32'h10408000;
      41313: inst = 32'hc40567b;
      41314: inst = 32'h8220000;
      41315: inst = 32'h10408000;
      41316: inst = 32'hc40567c;
      41317: inst = 32'h8220000;
      41318: inst = 32'h10408000;
      41319: inst = 32'hc40567d;
      41320: inst = 32'h8220000;
      41321: inst = 32'h10408000;
      41322: inst = 32'hc40567e;
      41323: inst = 32'h8220000;
      41324: inst = 32'h10408000;
      41325: inst = 32'hc40567f;
      41326: inst = 32'h8220000;
      41327: inst = 32'h10408000;
      41328: inst = 32'hc405680;
      41329: inst = 32'h8220000;
      41330: inst = 32'h10408000;
      41331: inst = 32'hc405681;
      41332: inst = 32'h8220000;
      41333: inst = 32'h10408000;
      41334: inst = 32'hc405682;
      41335: inst = 32'h8220000;
      41336: inst = 32'h10408000;
      41337: inst = 32'hc405683;
      41338: inst = 32'h8220000;
      41339: inst = 32'h10408000;
      41340: inst = 32'hc405684;
      41341: inst = 32'h8220000;
      41342: inst = 32'h10408000;
      41343: inst = 32'hc405685;
      41344: inst = 32'h8220000;
      41345: inst = 32'h10408000;
      41346: inst = 32'hc405686;
      41347: inst = 32'h8220000;
      41348: inst = 32'h10408000;
      41349: inst = 32'hc405687;
      41350: inst = 32'h8220000;
      41351: inst = 32'h10408000;
      41352: inst = 32'hc405688;
      41353: inst = 32'h8220000;
      41354: inst = 32'h10408000;
      41355: inst = 32'hc405689;
      41356: inst = 32'h8220000;
      41357: inst = 32'h10408000;
      41358: inst = 32'hc40568a;
      41359: inst = 32'h8220000;
      41360: inst = 32'h10408000;
      41361: inst = 32'hc40568b;
      41362: inst = 32'h8220000;
      41363: inst = 32'h10408000;
      41364: inst = 32'hc40568c;
      41365: inst = 32'h8220000;
      41366: inst = 32'h10408000;
      41367: inst = 32'hc40568d;
      41368: inst = 32'h8220000;
      41369: inst = 32'h10408000;
      41370: inst = 32'hc40568e;
      41371: inst = 32'h8220000;
      41372: inst = 32'h10408000;
      41373: inst = 32'hc40568f;
      41374: inst = 32'h8220000;
      41375: inst = 32'h10408000;
      41376: inst = 32'hc405690;
      41377: inst = 32'h8220000;
      41378: inst = 32'h10408000;
      41379: inst = 32'hc405691;
      41380: inst = 32'h8220000;
      41381: inst = 32'h10408000;
      41382: inst = 32'hc405692;
      41383: inst = 32'h8220000;
      41384: inst = 32'h10408000;
      41385: inst = 32'hc405693;
      41386: inst = 32'h8220000;
      41387: inst = 32'h10408000;
      41388: inst = 32'hc405694;
      41389: inst = 32'h8220000;
      41390: inst = 32'h10408000;
      41391: inst = 32'hc405695;
      41392: inst = 32'h8220000;
      41393: inst = 32'h10408000;
      41394: inst = 32'hc405696;
      41395: inst = 32'h8220000;
      41396: inst = 32'h10408000;
      41397: inst = 32'hc405697;
      41398: inst = 32'h8220000;
      41399: inst = 32'h10408000;
      41400: inst = 32'hc405698;
      41401: inst = 32'h8220000;
      41402: inst = 32'h10408000;
      41403: inst = 32'hc405699;
      41404: inst = 32'h8220000;
      41405: inst = 32'h10408000;
      41406: inst = 32'hc40569a;
      41407: inst = 32'h8220000;
      41408: inst = 32'h10408000;
      41409: inst = 32'hc40569b;
      41410: inst = 32'h8220000;
      41411: inst = 32'h10408000;
      41412: inst = 32'hc40569c;
      41413: inst = 32'h8220000;
      41414: inst = 32'h10408000;
      41415: inst = 32'hc40569d;
      41416: inst = 32'h8220000;
      41417: inst = 32'h10408000;
      41418: inst = 32'hc40569e;
      41419: inst = 32'h8220000;
      41420: inst = 32'h10408000;
      41421: inst = 32'hc40569f;
      41422: inst = 32'h8220000;
      41423: inst = 32'h10408000;
      41424: inst = 32'hc4056a0;
      41425: inst = 32'h8220000;
      41426: inst = 32'h10408000;
      41427: inst = 32'hc4056a1;
      41428: inst = 32'h8220000;
      41429: inst = 32'h10408000;
      41430: inst = 32'hc4056a2;
      41431: inst = 32'h8220000;
      41432: inst = 32'h10408000;
      41433: inst = 32'hc4056a3;
      41434: inst = 32'h8220000;
      41435: inst = 32'h10408000;
      41436: inst = 32'hc4056a4;
      41437: inst = 32'h8220000;
      41438: inst = 32'h10408000;
      41439: inst = 32'hc4056a5;
      41440: inst = 32'h8220000;
      41441: inst = 32'h10408000;
      41442: inst = 32'hc4056a6;
      41443: inst = 32'h8220000;
      41444: inst = 32'h10408000;
      41445: inst = 32'hc4056a7;
      41446: inst = 32'h8220000;
      41447: inst = 32'h10408000;
      41448: inst = 32'hc4056a8;
      41449: inst = 32'h8220000;
      41450: inst = 32'h10408000;
      41451: inst = 32'hc4056a9;
      41452: inst = 32'h8220000;
      41453: inst = 32'h10408000;
      41454: inst = 32'hc4056aa;
      41455: inst = 32'h8220000;
      41456: inst = 32'h10408000;
      41457: inst = 32'hc4056ab;
      41458: inst = 32'h8220000;
      41459: inst = 32'h10408000;
      41460: inst = 32'hc4056ac;
      41461: inst = 32'h8220000;
      41462: inst = 32'h10408000;
      41463: inst = 32'hc4056ad;
      41464: inst = 32'h8220000;
      41465: inst = 32'h10408000;
      41466: inst = 32'hc4056ae;
      41467: inst = 32'h8220000;
      41468: inst = 32'h10408000;
      41469: inst = 32'hc4056af;
      41470: inst = 32'h8220000;
      41471: inst = 32'h10408000;
      41472: inst = 32'hc4056b0;
      41473: inst = 32'h8220000;
      41474: inst = 32'h10408000;
      41475: inst = 32'hc4056b1;
      41476: inst = 32'h8220000;
      41477: inst = 32'h10408000;
      41478: inst = 32'hc4056bc;
      41479: inst = 32'h8220000;
      41480: inst = 32'h10408000;
      41481: inst = 32'hc405711;
      41482: inst = 32'h8220000;
      41483: inst = 32'h10408000;
      41484: inst = 32'hc40571c;
      41485: inst = 32'h8220000;
      41486: inst = 32'h10408000;
      41487: inst = 32'hc405771;
      41488: inst = 32'h8220000;
      41489: inst = 32'h10408000;
      41490: inst = 32'hc40577c;
      41491: inst = 32'h8220000;
      41492: inst = 32'h10408000;
      41493: inst = 32'hc4057d1;
      41494: inst = 32'h8220000;
      41495: inst = 32'h10408000;
      41496: inst = 32'hc4057dc;
      41497: inst = 32'h8220000;
      41498: inst = 32'hc20cba6;
      41499: inst = 32'h10408000;
      41500: inst = 32'hc403fe4;
      41501: inst = 32'h8220000;
      41502: inst = 32'h10408000;
      41503: inst = 32'hc403fec;
      41504: inst = 32'h8220000;
      41505: inst = 32'h10408000;
      41506: inst = 32'hc4040ac;
      41507: inst = 32'h8220000;
      41508: inst = 32'h10408000;
      41509: inst = 32'hc40410c;
      41510: inst = 32'h8220000;
      41511: inst = 32'h10408000;
      41512: inst = 32'hc40416c;
      41513: inst = 32'h8220000;
      41514: inst = 32'h10408000;
      41515: inst = 32'hc4041c4;
      41516: inst = 32'h8220000;
      41517: inst = 32'h10408000;
      41518: inst = 32'hc404224;
      41519: inst = 32'h8220000;
      41520: inst = 32'h10408000;
      41521: inst = 32'hc404284;
      41522: inst = 32'h8220000;
      41523: inst = 32'h10408000;
      41524: inst = 32'hc40428c;
      41525: inst = 32'h8220000;
      41526: inst = 32'h10408000;
      41527: inst = 32'hc4042e4;
      41528: inst = 32'h8220000;
      41529: inst = 32'h10408000;
      41530: inst = 32'hc4042ec;
      41531: inst = 32'h8220000;
      41532: inst = 32'h10408000;
      41533: inst = 32'hc404344;
      41534: inst = 32'h8220000;
      41535: inst = 32'h10408000;
      41536: inst = 32'hc40434c;
      41537: inst = 32'h8220000;
      41538: inst = 32'h10408000;
      41539: inst = 32'hc4054d2;
      41540: inst = 32'h8220000;
      41541: inst = 32'hc20cb44;
      41542: inst = 32'h10408000;
      41543: inst = 32'hc403fe5;
      41544: inst = 32'h8220000;
      41545: inst = 32'h10408000;
      41546: inst = 32'hc403fe6;
      41547: inst = 32'h8220000;
      41548: inst = 32'h10408000;
      41549: inst = 32'hc403fe7;
      41550: inst = 32'h8220000;
      41551: inst = 32'h10408000;
      41552: inst = 32'hc403fe8;
      41553: inst = 32'h8220000;
      41554: inst = 32'h10408000;
      41555: inst = 32'hc403fe9;
      41556: inst = 32'h8220000;
      41557: inst = 32'h10408000;
      41558: inst = 32'hc403fea;
      41559: inst = 32'h8220000;
      41560: inst = 32'h10408000;
      41561: inst = 32'hc403feb;
      41562: inst = 32'h8220000;
      41563: inst = 32'h10408000;
      41564: inst = 32'hc404104;
      41565: inst = 32'h8220000;
      41566: inst = 32'h10408000;
      41567: inst = 32'hc4043a6;
      41568: inst = 32'h8220000;
      41569: inst = 32'h10408000;
      41570: inst = 32'hc4043a7;
      41571: inst = 32'h8220000;
      41572: inst = 32'h10408000;
      41573: inst = 32'hc4043a8;
      41574: inst = 32'h8220000;
      41575: inst = 32'h10408000;
      41576: inst = 32'hc4043a9;
      41577: inst = 32'h8220000;
      41578: inst = 32'h10408000;
      41579: inst = 32'hc4043aa;
      41580: inst = 32'h8220000;
      41581: inst = 32'h10408000;
      41582: inst = 32'hc4043ab;
      41583: inst = 32'h8220000;
      41584: inst = 32'h10408000;
      41585: inst = 32'hc405354;
      41586: inst = 32'h8220000;
      41587: inst = 32'h10408000;
      41588: inst = 32'hc4053b2;
      41589: inst = 32'h8220000;
      41590: inst = 32'h10408000;
      41591: inst = 32'hc405532;
      41592: inst = 32'h8220000;
      41593: inst = 32'hc20a5f0;
      41594: inst = 32'h10408000;
      41595: inst = 32'hc403fed;
      41596: inst = 32'h8220000;
      41597: inst = 32'hc203d29;
      41598: inst = 32'h10408000;
      41599: inst = 32'hc403fee;
      41600: inst = 32'h8220000;
      41601: inst = 32'hc203ca9;
      41602: inst = 32'h10408000;
      41603: inst = 32'hc403fef;
      41604: inst = 32'h8220000;
      41605: inst = 32'hc20448a;
      41606: inst = 32'h10408000;
      41607: inst = 32'hc403ff0;
      41608: inst = 32'h8220000;
      41609: inst = 32'hc20636f;
      41610: inst = 32'h10408000;
      41611: inst = 32'hc403ff1;
      41612: inst = 32'h8220000;
      41613: inst = 32'h10408000;
      41614: inst = 32'hc403ff7;
      41615: inst = 32'h8220000;
      41616: inst = 32'h10408000;
      41617: inst = 32'hc404053;
      41618: inst = 32'h8220000;
      41619: inst = 32'h10408000;
      41620: inst = 32'hc404675;
      41621: inst = 32'h8220000;
      41622: inst = 32'h10408000;
      41623: inst = 32'hc404677;
      41624: inst = 32'h8220000;
      41625: inst = 32'h10408000;
      41626: inst = 32'hc4046ca;
      41627: inst = 32'h8220000;
      41628: inst = 32'h10408000;
      41629: inst = 32'hc4046d5;
      41630: inst = 32'h8220000;
      41631: inst = 32'h10408000;
      41632: inst = 32'hc404732;
      41633: inst = 32'h8220000;
      41634: inst = 32'hc2053ac;
      41635: inst = 32'h10408000;
      41636: inst = 32'hc403ff2;
      41637: inst = 32'h8220000;
      41638: inst = 32'hc203427;
      41639: inst = 32'h10408000;
      41640: inst = 32'hc403ff3;
      41641: inst = 32'h8220000;
      41642: inst = 32'hc20638f;
      41643: inst = 32'h10408000;
      41644: inst = 32'hc403ff4;
      41645: inst = 32'h8220000;
      41646: inst = 32'hc204bac;
      41647: inst = 32'h10408000;
      41648: inst = 32'hc403ff6;
      41649: inst = 32'h8220000;
      41650: inst = 32'h10408000;
      41651: inst = 32'hc40404e;
      41652: inst = 32'h8220000;
      41653: inst = 32'hc204549;
      41654: inst = 32'h10408000;
      41655: inst = 32'hc403ffa;
      41656: inst = 32'h8220000;
      41657: inst = 32'hc20546c;
      41658: inst = 32'h10408000;
      41659: inst = 32'hc403ffb;
      41660: inst = 32'h8220000;
      41661: inst = 32'hc20544d;
      41662: inst = 32'h10408000;
      41663: inst = 32'hc403ffc;
      41664: inst = 32'h8220000;
      41665: inst = 32'hc20cb86;
      41666: inst = 32'h10408000;
      41667: inst = 32'hc404044;
      41668: inst = 32'h8220000;
      41669: inst = 32'hc20dba5;
      41670: inst = 32'h10408000;
      41671: inst = 32'hc404045;
      41672: inst = 32'h8220000;
      41673: inst = 32'h10408000;
      41674: inst = 32'hc4041c6;
      41675: inst = 32'h8220000;
      41676: inst = 32'h10408000;
      41677: inst = 32'hc4041c7;
      41678: inst = 32'h8220000;
      41679: inst = 32'h10408000;
      41680: inst = 32'hc40428a;
      41681: inst = 32'h8220000;
      41682: inst = 32'h10408000;
      41683: inst = 32'hc404345;
      41684: inst = 32'h8220000;
      41685: inst = 32'h10408000;
      41686: inst = 32'hc4053b4;
      41687: inst = 32'h8220000;
      41688: inst = 32'h10408000;
      41689: inst = 32'hc405713;
      41690: inst = 32'h8220000;
      41691: inst = 32'hc20dbc5;
      41692: inst = 32'h10408000;
      41693: inst = 32'hc404046;
      41694: inst = 32'h8220000;
      41695: inst = 32'h10408000;
      41696: inst = 32'hc404047;
      41697: inst = 32'h8220000;
      41698: inst = 32'h10408000;
      41699: inst = 32'hc4040a9;
      41700: inst = 32'h8220000;
      41701: inst = 32'h10408000;
      41702: inst = 32'hc4040aa;
      41703: inst = 32'h8220000;
      41704: inst = 32'h10408000;
      41705: inst = 32'hc4040ab;
      41706: inst = 32'h8220000;
      41707: inst = 32'h10408000;
      41708: inst = 32'hc404109;
      41709: inst = 32'h8220000;
      41710: inst = 32'h10408000;
      41711: inst = 32'hc40410a;
      41712: inst = 32'h8220000;
      41713: inst = 32'h10408000;
      41714: inst = 32'hc40410b;
      41715: inst = 32'h8220000;
      41716: inst = 32'h10408000;
      41717: inst = 32'hc404169;
      41718: inst = 32'h8220000;
      41719: inst = 32'h10408000;
      41720: inst = 32'hc4041c8;
      41721: inst = 32'h8220000;
      41722: inst = 32'h10408000;
      41723: inst = 32'hc4041c9;
      41724: inst = 32'h8220000;
      41725: inst = 32'h10408000;
      41726: inst = 32'hc404226;
      41727: inst = 32'h8220000;
      41728: inst = 32'h10408000;
      41729: inst = 32'hc404227;
      41730: inst = 32'h8220000;
      41731: inst = 32'h10408000;
      41732: inst = 32'hc404228;
      41733: inst = 32'h8220000;
      41734: inst = 32'h10408000;
      41735: inst = 32'hc404286;
      41736: inst = 32'h8220000;
      41737: inst = 32'h10408000;
      41738: inst = 32'hc404287;
      41739: inst = 32'h8220000;
      41740: inst = 32'h10408000;
      41741: inst = 32'hc404288;
      41742: inst = 32'h8220000;
      41743: inst = 32'h10408000;
      41744: inst = 32'hc404289;
      41745: inst = 32'h8220000;
      41746: inst = 32'h10408000;
      41747: inst = 32'hc4042e6;
      41748: inst = 32'h8220000;
      41749: inst = 32'h10408000;
      41750: inst = 32'hc4042e7;
      41751: inst = 32'h8220000;
      41752: inst = 32'h10408000;
      41753: inst = 32'hc4042e8;
      41754: inst = 32'h8220000;
      41755: inst = 32'h10408000;
      41756: inst = 32'hc4042e9;
      41757: inst = 32'h8220000;
      41758: inst = 32'h10408000;
      41759: inst = 32'hc4042ea;
      41760: inst = 32'h8220000;
      41761: inst = 32'h10408000;
      41762: inst = 32'hc4042eb;
      41763: inst = 32'h8220000;
      41764: inst = 32'h10408000;
      41765: inst = 32'hc405594;
      41766: inst = 32'h8220000;
      41767: inst = 32'h10408000;
      41768: inst = 32'hc4055f4;
      41769: inst = 32'h8220000;
      41770: inst = 32'h10408000;
      41771: inst = 32'hc405653;
      41772: inst = 32'h8220000;
      41773: inst = 32'hc20dbc6;
      41774: inst = 32'h10408000;
      41775: inst = 32'hc404048;
      41776: inst = 32'h8220000;
      41777: inst = 32'h10408000;
      41778: inst = 32'hc404049;
      41779: inst = 32'h8220000;
      41780: inst = 32'h10408000;
      41781: inst = 32'hc40404a;
      41782: inst = 32'h8220000;
      41783: inst = 32'h10408000;
      41784: inst = 32'hc404229;
      41785: inst = 32'h8220000;
      41786: inst = 32'h10408000;
      41787: inst = 32'hc404347;
      41788: inst = 32'h8220000;
      41789: inst = 32'h10408000;
      41790: inst = 32'hc404348;
      41791: inst = 32'h8220000;
      41792: inst = 32'h10408000;
      41793: inst = 32'hc404349;
      41794: inst = 32'h8220000;
      41795: inst = 32'h10408000;
      41796: inst = 32'hc40434a;
      41797: inst = 32'h8220000;
      41798: inst = 32'h10408000;
      41799: inst = 32'hc4055f3;
      41800: inst = 32'h8220000;
      41801: inst = 32'hc20e3c6;
      41802: inst = 32'h10408000;
      41803: inst = 32'hc40404b;
      41804: inst = 32'h8220000;
      41805: inst = 32'h10408000;
      41806: inst = 32'hc404346;
      41807: inst = 32'h8220000;
      41808: inst = 32'h10408000;
      41809: inst = 32'hc40434b;
      41810: inst = 32'h8220000;
      41811: inst = 32'h10408000;
      41812: inst = 32'hc405654;
      41813: inst = 32'h8220000;
      41814: inst = 32'hc20cb85;
      41815: inst = 32'h10408000;
      41816: inst = 32'hc40404c;
      41817: inst = 32'h8220000;
      41818: inst = 32'hc206d0b;
      41819: inst = 32'h10408000;
      41820: inst = 32'hc40404d;
      41821: inst = 32'h8220000;
      41822: inst = 32'hc205c2d;
      41823: inst = 32'h10408000;
      41824: inst = 32'hc40404f;
      41825: inst = 32'h8220000;
      41826: inst = 32'hc203d88;
      41827: inst = 32'h10408000;
      41828: inst = 32'hc404050;
      41829: inst = 32'h8220000;
      41830: inst = 32'hc206b6f;
      41831: inst = 32'h10408000;
      41832: inst = 32'hc404051;
      41833: inst = 32'h8220000;
      41834: inst = 32'h10408000;
      41835: inst = 32'hc40466d;
      41836: inst = 32'h8220000;
      41837: inst = 32'h10408000;
      41838: inst = 32'hc4046d7;
      41839: inst = 32'h8220000;
      41840: inst = 32'h10408000;
      41841: inst = 32'hc40472e;
      41842: inst = 32'h8220000;
      41843: inst = 32'hc206b4f;
      41844: inst = 32'h10408000;
      41845: inst = 32'hc404052;
      41846: inst = 32'h8220000;
      41847: inst = 32'h10408000;
      41848: inst = 32'hc4056b6;
      41849: inst = 32'h8220000;
      41850: inst = 32'hc20542d;
      41851: inst = 32'h10408000;
      41852: inst = 32'hc404055;
      41853: inst = 32'h8220000;
      41854: inst = 32'h10408000;
      41855: inst = 32'hc4040b1;
      41856: inst = 32'h8220000;
      41857: inst = 32'hc205bee;
      41858: inst = 32'h10408000;
      41859: inst = 32'hc404056;
      41860: inst = 32'h8220000;
      41861: inst = 32'h10408000;
      41862: inst = 32'hc4040b5;
      41863: inst = 32'h8220000;
      41864: inst = 32'hc2063af;
      41865: inst = 32'h10408000;
      41866: inst = 32'hc404059;
      41867: inst = 32'h8220000;
      41868: inst = 32'hc203d49;
      41869: inst = 32'h10408000;
      41870: inst = 32'hc40405a;
      41871: inst = 32'h8220000;
      41872: inst = 32'hc206b70;
      41873: inst = 32'h10408000;
      41874: inst = 32'hc40405b;
      41875: inst = 32'h8220000;
      41876: inst = 32'h10408000;
      41877: inst = 32'hc404679;
      41878: inst = 32'h8220000;
      41879: inst = 32'h10408000;
      41880: inst = 32'hc40472d;
      41881: inst = 32'h8220000;
      41882: inst = 32'h10408000;
      41883: inst = 32'hc404730;
      41884: inst = 32'h8220000;
      41885: inst = 32'hc20cb64;
      41886: inst = 32'h10408000;
      41887: inst = 32'hc4040a4;
      41888: inst = 32'h8220000;
      41889: inst = 32'h10408000;
      41890: inst = 32'hc404164;
      41891: inst = 32'h8220000;
      41892: inst = 32'hc20dc08;
      41893: inst = 32'h10408000;
      41894: inst = 32'hc4040a5;
      41895: inst = 32'h8220000;
      41896: inst = 32'hc20f77b;
      41897: inst = 32'h10408000;
      41898: inst = 32'hc4040a6;
      41899: inst = 32'h8220000;
      41900: inst = 32'h10408000;
      41901: inst = 32'hc404154;
      41902: inst = 32'h8220000;
      41903: inst = 32'h10408000;
      41904: inst = 32'hc404155;
      41905: inst = 32'h8220000;
      41906: inst = 32'h10408000;
      41907: inst = 32'hc4041b0;
      41908: inst = 32'h8220000;
      41909: inst = 32'h10408000;
      41910: inst = 32'hc4041b7;
      41911: inst = 32'h8220000;
      41912: inst = 32'h10408000;
      41913: inst = 32'hc404274;
      41914: inst = 32'h8220000;
      41915: inst = 32'h10408000;
      41916: inst = 32'hc40427a;
      41917: inst = 32'h8220000;
      41918: inst = 32'h10408000;
      41919: inst = 32'hc404339;
      41920: inst = 32'h8220000;
      41921: inst = 32'h10408000;
      41922: inst = 32'hc4043fa;
      41923: inst = 32'h8220000;
      41924: inst = 32'h10408000;
      41925: inst = 32'hc404453;
      41926: inst = 32'h8220000;
      41927: inst = 32'h10408000;
      41928: inst = 32'hc404458;
      41929: inst = 32'h8220000;
      41930: inst = 32'h10408000;
      41931: inst = 32'hc4044b6;
      41932: inst = 32'h8220000;
      41933: inst = 32'h10408000;
      41934: inst = 32'hc4044ba;
      41935: inst = 32'h8220000;
      41936: inst = 32'h10408000;
      41937: inst = 32'hc404519;
      41938: inst = 32'h8220000;
      41939: inst = 32'h10408000;
      41940: inst = 32'hc4045d3;
      41941: inst = 32'h8220000;
      41942: inst = 32'hc20e48a;
      41943: inst = 32'h10408000;
      41944: inst = 32'hc4040a7;
      41945: inst = 32'h8220000;
      41946: inst = 32'hc20db84;
      41947: inst = 32'h10408000;
      41948: inst = 32'hc4040a8;
      41949: inst = 32'h8220000;
      41950: inst = 32'h10408000;
      41951: inst = 32'hc404108;
      41952: inst = 32'h8220000;
      41953: inst = 32'h10408000;
      41954: inst = 32'hc404168;
      41955: inst = 32'h8220000;
      41956: inst = 32'hc20a5d0;
      41957: inst = 32'h10408000;
      41958: inst = 32'hc4040ad;
      41959: inst = 32'h8220000;
      41960: inst = 32'h10408000;
      41961: inst = 32'hc404231;
      41962: inst = 32'h8220000;
      41963: inst = 32'h10408000;
      41964: inst = 32'hc404290;
      41965: inst = 32'h8220000;
      41966: inst = 32'hc205b6e;
      41967: inst = 32'h10408000;
      41968: inst = 32'hc4040ae;
      41969: inst = 32'h8220000;
      41970: inst = 32'hc204ccb;
      41971: inst = 32'h10408000;
      41972: inst = 32'hc4040b0;
      41973: inst = 32'h8220000;
      41974: inst = 32'h10408000;
      41975: inst = 32'hc4040ba;
      41976: inst = 32'h8220000;
      41977: inst = 32'hc2043aa;
      41978: inst = 32'h10408000;
      41979: inst = 32'hc4040b3;
      41980: inst = 32'h8220000;
      41981: inst = 32'h10408000;
      41982: inst = 32'hc4040b4;
      41983: inst = 32'h8220000;
      41984: inst = 32'hc2063ae;
      41985: inst = 32'h10408000;
      41986: inst = 32'hc4040b6;
      41987: inst = 32'h8220000;
      41988: inst = 32'h10408000;
      41989: inst = 32'hc40466a;
      41990: inst = 32'h8220000;
      41991: inst = 32'h10408000;
      41992: inst = 32'hc4046cd;
      41993: inst = 32'h8220000;
      41994: inst = 32'hc20544c;
      41995: inst = 32'h10408000;
      41996: inst = 32'hc4040b9;
      41997: inst = 32'h8220000;
      41998: inst = 32'h10408000;
      41999: inst = 32'hc4046cc;
      42000: inst = 32'h8220000;
      42001: inst = 32'h10408000;
      42002: inst = 32'hc40472b;
      42003: inst = 32'h8220000;
      42004: inst = 32'hc20dc28;
      42005: inst = 32'h10408000;
      42006: inst = 32'hc404105;
      42007: inst = 32'h8220000;
      42008: inst = 32'h10408000;
      42009: inst = 32'hc405533;
      42010: inst = 32'h8220000;
      42011: inst = 32'hc20ffff;
      42012: inst = 32'h10408000;
      42013: inst = 32'hc404106;
      42014: inst = 32'h8220000;
      42015: inst = 32'h10408000;
      42016: inst = 32'hc40439b;
      42017: inst = 32'h8220000;
      42018: inst = 32'h10408000;
      42019: inst = 32'hc404515;
      42020: inst = 32'h8220000;
      42021: inst = 32'hc20e4cc;
      42022: inst = 32'h10408000;
      42023: inst = 32'hc404107;
      42024: inst = 32'h8220000;
      42025: inst = 32'h10408000;
      42026: inst = 32'hc404167;
      42027: inst = 32'h8220000;
      42028: inst = 32'hc20ce94;
      42029: inst = 32'h10408000;
      42030: inst = 32'hc40410d;
      42031: inst = 32'h8220000;
      42032: inst = 32'hc20c632;
      42033: inst = 32'h10408000;
      42034: inst = 32'hc404113;
      42035: inst = 32'h8220000;
      42036: inst = 32'hc204ca9;
      42037: inst = 32'h10408000;
      42038: inst = 32'hc404114;
      42039: inst = 32'h8220000;
      42040: inst = 32'hc207e0d;
      42041: inst = 32'h10408000;
      42042: inst = 32'hc404116;
      42043: inst = 32'h8220000;
      42044: inst = 32'hc20d694;
      42045: inst = 32'h10408000;
      42046: inst = 32'hc404117;
      42047: inst = 32'h8220000;
      42048: inst = 32'h10408000;
      42049: inst = 32'hc4047f3;
      42050: inst = 32'h8220000;
      42051: inst = 32'h10408000;
      42052: inst = 32'hc404919;
      42053: inst = 32'h8220000;
      42054: inst = 32'hc20eed7;
      42055: inst = 32'h10408000;
      42056: inst = 32'hc404151;
      42057: inst = 32'h8220000;
      42058: inst = 32'h10408000;
      42059: inst = 32'hc4041b4;
      42060: inst = 32'h8220000;
      42061: inst = 32'h10408000;
      42062: inst = 32'hc404217;
      42063: inst = 32'h8220000;
      42064: inst = 32'h10408000;
      42065: inst = 32'hc404218;
      42066: inst = 32'h8220000;
      42067: inst = 32'h10408000;
      42068: inst = 32'hc404270;
      42069: inst = 32'h8220000;
      42070: inst = 32'h10408000;
      42071: inst = 32'hc404277;
      42072: inst = 32'h8220000;
      42073: inst = 32'h10408000;
      42074: inst = 32'hc4042d0;
      42075: inst = 32'h8220000;
      42076: inst = 32'h10408000;
      42077: inst = 32'hc4042d4;
      42078: inst = 32'h8220000;
      42079: inst = 32'h10408000;
      42080: inst = 32'hc404391;
      42081: inst = 32'h8220000;
      42082: inst = 32'h10408000;
      42083: inst = 32'hc404450;
      42084: inst = 32'h8220000;
      42085: inst = 32'h10408000;
      42086: inst = 32'hc404451;
      42087: inst = 32'h8220000;
      42088: inst = 32'h10408000;
      42089: inst = 32'hc404454;
      42090: inst = 32'h8220000;
      42091: inst = 32'h10408000;
      42092: inst = 32'hc40445b;
      42093: inst = 32'h8220000;
      42094: inst = 32'h10408000;
      42095: inst = 32'hc40451c;
      42096: inst = 32'h8220000;
      42097: inst = 32'h10408000;
      42098: inst = 32'hc4053c8;
      42099: inst = 32'h8220000;
      42100: inst = 32'h10408000;
      42101: inst = 32'hc4053ce;
      42102: inst = 32'h8220000;
      42103: inst = 32'hc20f73a;
      42104: inst = 32'h10408000;
      42105: inst = 32'hc404152;
      42106: inst = 32'h8220000;
      42107: inst = 32'h10408000;
      42108: inst = 32'hc40415b;
      42109: inst = 32'h8220000;
      42110: inst = 32'h10408000;
      42111: inst = 32'hc40415c;
      42112: inst = 32'h8220000;
      42113: inst = 32'h10408000;
      42114: inst = 32'hc40421a;
      42115: inst = 32'h8220000;
      42116: inst = 32'h10408000;
      42117: inst = 32'hc4042d7;
      42118: inst = 32'h8220000;
      42119: inst = 32'h10408000;
      42120: inst = 32'hc4042d8;
      42121: inst = 32'h8220000;
      42122: inst = 32'h10408000;
      42123: inst = 32'hc4042d9;
      42124: inst = 32'h8220000;
      42125: inst = 32'h10408000;
      42126: inst = 32'hc40433b;
      42127: inst = 32'h8220000;
      42128: inst = 32'h10408000;
      42129: inst = 32'hc40439c;
      42130: inst = 32'h8220000;
      42131: inst = 32'h10408000;
      42132: inst = 32'hc4044b3;
      42133: inst = 32'h8220000;
      42134: inst = 32'h10408000;
      42135: inst = 32'hc4044b5;
      42136: inst = 32'h8220000;
      42137: inst = 32'h10408000;
      42138: inst = 32'hc404577;
      42139: inst = 32'h8220000;
      42140: inst = 32'h10408000;
      42141: inst = 32'hc4045d8;
      42142: inst = 32'h8220000;
      42143: inst = 32'h10408000;
      42144: inst = 32'hc4045d9;
      42145: inst = 32'h8220000;
      42146: inst = 32'hc20f75b;
      42147: inst = 32'h10408000;
      42148: inst = 32'hc404153;
      42149: inst = 32'h8220000;
      42150: inst = 32'h10408000;
      42151: inst = 32'hc404157;
      42152: inst = 32'h8220000;
      42153: inst = 32'h10408000;
      42154: inst = 32'hc4041b2;
      42155: inst = 32'h8220000;
      42156: inst = 32'h10408000;
      42157: inst = 32'hc404271;
      42158: inst = 32'h8220000;
      42159: inst = 32'h10408000;
      42160: inst = 32'hc404276;
      42161: inst = 32'h8220000;
      42162: inst = 32'h10408000;
      42163: inst = 32'hc4042dc;
      42164: inst = 32'h8220000;
      42165: inst = 32'h10408000;
      42166: inst = 32'hc404336;
      42167: inst = 32'h8220000;
      42168: inst = 32'h10408000;
      42169: inst = 32'hc404394;
      42170: inst = 32'h8220000;
      42171: inst = 32'h10408000;
      42172: inst = 32'hc4043f0;
      42173: inst = 32'h8220000;
      42174: inst = 32'h10408000;
      42175: inst = 32'hc4043fb;
      42176: inst = 32'h8220000;
      42177: inst = 32'h10408000;
      42178: inst = 32'hc404510;
      42179: inst = 32'h8220000;
      42180: inst = 32'h10408000;
      42181: inst = 32'hc404516;
      42182: inst = 32'h8220000;
      42183: inst = 32'h10408000;
      42184: inst = 32'hc404574;
      42185: inst = 32'h8220000;
      42186: inst = 32'hc20f739;
      42187: inst = 32'h10408000;
      42188: inst = 32'hc404156;
      42189: inst = 32'h8220000;
      42190: inst = 32'h10408000;
      42191: inst = 32'hc4041b6;
      42192: inst = 32'h8220000;
      42193: inst = 32'h10408000;
      42194: inst = 32'hc404213;
      42195: inst = 32'h8220000;
      42196: inst = 32'h10408000;
      42197: inst = 32'hc404399;
      42198: inst = 32'h8220000;
      42199: inst = 32'h10408000;
      42200: inst = 32'hc404517;
      42201: inst = 32'h8220000;
      42202: inst = 32'h10408000;
      42203: inst = 32'hc404576;
      42204: inst = 32'h8220000;
      42205: inst = 32'h10408000;
      42206: inst = 32'hc4045d1;
      42207: inst = 32'h8220000;
      42208: inst = 32'h10408000;
      42209: inst = 32'hc4045dc;
      42210: inst = 32'h8220000;
      42211: inst = 32'hc20ffde;
      42212: inst = 32'h10408000;
      42213: inst = 32'hc404158;
      42214: inst = 32'h8220000;
      42215: inst = 32'h10408000;
      42216: inst = 32'hc4041b9;
      42217: inst = 32'h8220000;
      42218: inst = 32'h10408000;
      42219: inst = 32'hc404392;
      42220: inst = 32'h8220000;
      42221: inst = 32'h10408000;
      42222: inst = 32'hc4043f2;
      42223: inst = 32'h8220000;
      42224: inst = 32'h10408000;
      42225: inst = 32'hc4043f7;
      42226: inst = 32'h8220000;
      42227: inst = 32'h10408000;
      42228: inst = 32'hc4044b9;
      42229: inst = 32'h8220000;
      42230: inst = 32'hc20f75a;
      42231: inst = 32'h10408000;
      42232: inst = 32'hc404159;
      42233: inst = 32'h8220000;
      42234: inst = 32'h10408000;
      42235: inst = 32'hc40415a;
      42236: inst = 32'h8220000;
      42237: inst = 32'h10408000;
      42238: inst = 32'hc404272;
      42239: inst = 32'h8220000;
      42240: inst = 32'h10408000;
      42241: inst = 32'hc404273;
      42242: inst = 32'h8220000;
      42243: inst = 32'h10408000;
      42244: inst = 32'hc404331;
      42245: inst = 32'h8220000;
      42246: inst = 32'h10408000;
      42247: inst = 32'hc4043f3;
      42248: inst = 32'h8220000;
      42249: inst = 32'h10408000;
      42250: inst = 32'hc4043fc;
      42251: inst = 32'h8220000;
      42252: inst = 32'h10408000;
      42253: inst = 32'hc404452;
      42254: inst = 32'h8220000;
      42255: inst = 32'h10408000;
      42256: inst = 32'hc404456;
      42257: inst = 32'h8220000;
      42258: inst = 32'h10408000;
      42259: inst = 32'hc404459;
      42260: inst = 32'h8220000;
      42261: inst = 32'h10408000;
      42262: inst = 32'hc40445a;
      42263: inst = 32'h8220000;
      42264: inst = 32'h10408000;
      42265: inst = 32'hc4044bb;
      42266: inst = 32'h8220000;
      42267: inst = 32'h10408000;
      42268: inst = 32'hc40451a;
      42269: inst = 32'h8220000;
      42270: inst = 32'h10408000;
      42271: inst = 32'hc404570;
      42272: inst = 32'h8220000;
      42273: inst = 32'h10408000;
      42274: inst = 32'hc404573;
      42275: inst = 32'h8220000;
      42276: inst = 32'hc20dbe7;
      42277: inst = 32'h10408000;
      42278: inst = 32'hc404165;
      42279: inst = 32'h8220000;
      42280: inst = 32'hc20f77c;
      42281: inst = 32'h10408000;
      42282: inst = 32'hc404166;
      42283: inst = 32'h8220000;
      42284: inst = 32'h10408000;
      42285: inst = 32'hc4041b8;
      42286: inst = 32'h8220000;
      42287: inst = 32'hc20e3a4;
      42288: inst = 32'h10408000;
      42289: inst = 32'hc40416a;
      42290: inst = 32'h8220000;
      42291: inst = 32'h10408000;
      42292: inst = 32'hc405415;
      42293: inst = 32'h8220000;
      42294: inst = 32'h10408000;
      42295: inst = 32'hc405534;
      42296: inst = 32'h8220000;
      42297: inst = 32'h10408000;
      42298: inst = 32'hc405655;
      42299: inst = 32'h8220000;
      42300: inst = 32'hc20e3c5;
      42301: inst = 32'h10408000;
      42302: inst = 32'hc40416b;
      42303: inst = 32'h8220000;
      42304: inst = 32'h10408000;
      42305: inst = 32'hc40428b;
      42306: inst = 32'h8220000;
      42307: inst = 32'h10408000;
      42308: inst = 32'hc4053b5;
      42309: inst = 32'h8220000;
      42310: inst = 32'h10408000;
      42311: inst = 32'hc405595;
      42312: inst = 32'h8220000;
      42313: inst = 32'h10408000;
      42314: inst = 32'hc4055f5;
      42315: inst = 32'h8220000;
      42316: inst = 32'hc206e0c;
      42317: inst = 32'h10408000;
      42318: inst = 32'hc40416d;
      42319: inst = 32'h8220000;
      42320: inst = 32'hc209e50;
      42321: inst = 32'h10408000;
      42322: inst = 32'hc404176;
      42323: inst = 32'h8220000;
      42324: inst = 32'hc20860e;
      42325: inst = 32'h10408000;
      42326: inst = 32'hc404177;
      42327: inst = 32'h8220000;
      42328: inst = 32'hc20b5f1;
      42329: inst = 32'h10408000;
      42330: inst = 32'hc40417b;
      42331: inst = 32'h8220000;
      42332: inst = 32'hc20ffbd;
      42333: inst = 32'h10408000;
      42334: inst = 32'hc4041b1;
      42335: inst = 32'h8220000;
      42336: inst = 32'h10408000;
      42337: inst = 32'hc404279;
      42338: inst = 32'h8220000;
      42339: inst = 32'h10408000;
      42340: inst = 32'hc404332;
      42341: inst = 32'h8220000;
      42342: inst = 32'h10408000;
      42343: inst = 32'hc404396;
      42344: inst = 32'h8220000;
      42345: inst = 32'h10408000;
      42346: inst = 32'hc404457;
      42347: inst = 32'h8220000;
      42348: inst = 32'h10408000;
      42349: inst = 32'hc40445c;
      42350: inst = 32'h8220000;
      42351: inst = 32'h10408000;
      42352: inst = 32'hc4044bc;
      42353: inst = 32'h8220000;
      42354: inst = 32'hc20f6f8;
      42355: inst = 32'h10408000;
      42356: inst = 32'hc4041b3;
      42357: inst = 32'h8220000;
      42358: inst = 32'h10408000;
      42359: inst = 32'hc404215;
      42360: inst = 32'h8220000;
      42361: inst = 32'h10408000;
      42362: inst = 32'hc40421b;
      42363: inst = 32'h8220000;
      42364: inst = 32'h10408000;
      42365: inst = 32'hc4043f5;
      42366: inst = 32'h8220000;
      42367: inst = 32'h10408000;
      42368: inst = 32'hc4043f8;
      42369: inst = 32'h8220000;
      42370: inst = 32'h10408000;
      42371: inst = 32'hc404572;
      42372: inst = 32'h8220000;
      42373: inst = 32'hc20f719;
      42374: inst = 32'h10408000;
      42375: inst = 32'hc4041ba;
      42376: inst = 32'h8220000;
      42377: inst = 32'h10408000;
      42378: inst = 32'hc4041bb;
      42379: inst = 32'h8220000;
      42380: inst = 32'h10408000;
      42381: inst = 32'hc404335;
      42382: inst = 32'h8220000;
      42383: inst = 32'h10408000;
      42384: inst = 32'hc404337;
      42385: inst = 32'h8220000;
      42386: inst = 32'h10408000;
      42387: inst = 32'hc40433a;
      42388: inst = 32'h8220000;
      42389: inst = 32'h10408000;
      42390: inst = 32'hc404393;
      42391: inst = 32'h8220000;
      42392: inst = 32'h10408000;
      42393: inst = 32'hc4043f4;
      42394: inst = 32'h8220000;
      42395: inst = 32'h10408000;
      42396: inst = 32'hc4044b8;
      42397: inst = 32'h8220000;
      42398: inst = 32'h10408000;
      42399: inst = 32'hc404511;
      42400: inst = 32'h8220000;
      42401: inst = 32'h10408000;
      42402: inst = 32'hc404518;
      42403: inst = 32'h8220000;
      42404: inst = 32'h10408000;
      42405: inst = 32'hc40451b;
      42406: inst = 32'h8220000;
      42407: inst = 32'h10408000;
      42408: inst = 32'hc404575;
      42409: inst = 32'h8220000;
      42410: inst = 32'hc20ffbe;
      42411: inst = 32'h10408000;
      42412: inst = 32'hc4041bc;
      42413: inst = 32'h8220000;
      42414: inst = 32'h10408000;
      42415: inst = 32'hc404275;
      42416: inst = 32'h8220000;
      42417: inst = 32'hc20db85;
      42418: inst = 32'h10408000;
      42419: inst = 32'hc4041c5;
      42420: inst = 32'h8220000;
      42421: inst = 32'h10408000;
      42422: inst = 32'hc404225;
      42423: inst = 32'h8220000;
      42424: inst = 32'h10408000;
      42425: inst = 32'hc404285;
      42426: inst = 32'h8220000;
      42427: inst = 32'h10408000;
      42428: inst = 32'hc4042e5;
      42429: inst = 32'h8220000;
      42430: inst = 32'hc20c44c;
      42431: inst = 32'h10408000;
      42432: inst = 32'hc4041ca;
      42433: inst = 32'h8220000;
      42434: inst = 32'hc20cbe8;
      42435: inst = 32'h10408000;
      42436: inst = 32'hc4041cb;
      42437: inst = 32'h8220000;
      42438: inst = 32'hc20cba5;
      42439: inst = 32'h10408000;
      42440: inst = 32'hc4041cc;
      42441: inst = 32'h8220000;
      42442: inst = 32'h10408000;
      42443: inst = 32'hc40422c;
      42444: inst = 32'h8220000;
      42445: inst = 32'hc20c633;
      42446: inst = 32'h10408000;
      42447: inst = 32'hc4041d0;
      42448: inst = 32'h8220000;
      42449: inst = 32'hc205cca;
      42450: inst = 32'h10408000;
      42451: inst = 32'hc4041d1;
      42452: inst = 32'h8220000;
      42453: inst = 32'hc20e6b6;
      42454: inst = 32'h10408000;
      42455: inst = 32'hc4041d6;
      42456: inst = 32'h8220000;
      42457: inst = 32'h10408000;
      42458: inst = 32'hc40478f;
      42459: inst = 32'h8220000;
      42460: inst = 32'h10408000;
      42461: inst = 32'hc4047eb;
      42462: inst = 32'h8220000;
      42463: inst = 32'h10408000;
      42464: inst = 32'hc4047f2;
      42465: inst = 32'h8220000;
      42466: inst = 32'h10408000;
      42467: inst = 32'hc4048b6;
      42468: inst = 32'h8220000;
      42469: inst = 32'hc2055ca;
      42470: inst = 32'h10408000;
      42471: inst = 32'hc4041d7;
      42472: inst = 32'h8220000;
      42473: inst = 32'hc20de95;
      42474: inst = 32'h10408000;
      42475: inst = 32'hc4041d8;
      42476: inst = 32'h8220000;
      42477: inst = 32'h10408000;
      42478: inst = 32'hc40429b;
      42479: inst = 32'h8220000;
      42480: inst = 32'h10408000;
      42481: inst = 32'hc404792;
      42482: inst = 32'h8220000;
      42483: inst = 32'h10408000;
      42484: inst = 32'hc404798;
      42485: inst = 32'h8220000;
      42486: inst = 32'h10408000;
      42487: inst = 32'hc4047f5;
      42488: inst = 32'h8220000;
      42489: inst = 32'h10408000;
      42490: inst = 32'hc404857;
      42491: inst = 32'h8220000;
      42492: inst = 32'h10408000;
      42493: inst = 32'hc404915;
      42494: inst = 32'h8220000;
      42495: inst = 32'hc2054c9;
      42496: inst = 32'h10408000;
      42497: inst = 32'hc4041db;
      42498: inst = 32'h8220000;
      42499: inst = 32'h10408000;
      42500: inst = 32'hc404230;
      42501: inst = 32'h8220000;
      42502: inst = 32'hc20de75;
      42503: inst = 32'h10408000;
      42504: inst = 32'hc4041dc;
      42505: inst = 32'h8220000;
      42506: inst = 32'hc20f718;
      42507: inst = 32'h10408000;
      42508: inst = 32'hc404210;
      42509: inst = 32'h8220000;
      42510: inst = 32'h10408000;
      42511: inst = 32'hc404278;
      42512: inst = 32'h8220000;
      42513: inst = 32'hc20ff9d;
      42514: inst = 32'h10408000;
      42515: inst = 32'hc404211;
      42516: inst = 32'h8220000;
      42517: inst = 32'h10408000;
      42518: inst = 32'hc404219;
      42519: inst = 32'h8220000;
      42520: inst = 32'h10408000;
      42521: inst = 32'hc4042d6;
      42522: inst = 32'h8220000;
      42523: inst = 32'hc20ff9c;
      42524: inst = 32'h10408000;
      42525: inst = 32'hc404212;
      42526: inst = 32'h8220000;
      42527: inst = 32'h10408000;
      42528: inst = 32'hc404216;
      42529: inst = 32'h8220000;
      42530: inst = 32'h10408000;
      42531: inst = 32'hc40421c;
      42532: inst = 32'h8220000;
      42533: inst = 32'h10408000;
      42534: inst = 32'hc40427b;
      42535: inst = 32'h8220000;
      42536: inst = 32'h10408000;
      42537: inst = 32'hc4042d1;
      42538: inst = 32'h8220000;
      42539: inst = 32'h10408000;
      42540: inst = 32'hc4042d5;
      42541: inst = 32'h8220000;
      42542: inst = 32'h10408000;
      42543: inst = 32'hc40433c;
      42544: inst = 32'h8220000;
      42545: inst = 32'h10408000;
      42546: inst = 32'hc404395;
      42547: inst = 32'h8220000;
      42548: inst = 32'h10408000;
      42549: inst = 32'hc404397;
      42550: inst = 32'h8220000;
      42551: inst = 32'h10408000;
      42552: inst = 32'hc404398;
      42553: inst = 32'h8220000;
      42554: inst = 32'h10408000;
      42555: inst = 32'hc40439a;
      42556: inst = 32'h8220000;
      42557: inst = 32'h10408000;
      42558: inst = 32'hc4043f1;
      42559: inst = 32'h8220000;
      42560: inst = 32'h10408000;
      42561: inst = 32'hc404514;
      42562: inst = 32'h8220000;
      42563: inst = 32'h10408000;
      42564: inst = 32'hc4045d2;
      42565: inst = 32'h8220000;
      42566: inst = 32'hc20a46f;
      42567: inst = 32'h10408000;
      42568: inst = 32'hc40422a;
      42569: inst = 32'h8220000;
      42570: inst = 32'hc20d3c7;
      42571: inst = 32'h10408000;
      42572: inst = 32'hc40422b;
      42573: inst = 32'h8220000;
      42574: inst = 32'h10408000;
      42575: inst = 32'hc405475;
      42576: inst = 32'h8220000;
      42577: inst = 32'hc20ce53;
      42578: inst = 32'h10408000;
      42579: inst = 32'hc40422f;
      42580: inst = 32'h8220000;
      42581: inst = 32'hc207d4d;
      42582: inst = 32'h10408000;
      42583: inst = 32'hc40423b;
      42584: inst = 32'h8220000;
      42585: inst = 32'h10408000;
      42586: inst = 32'hc40423c;
      42587: inst = 32'h8220000;
      42588: inst = 32'hc20ff7c;
      42589: inst = 32'h10408000;
      42590: inst = 32'hc40427c;
      42591: inst = 32'h8220000;
      42592: inst = 32'h10408000;
      42593: inst = 32'hc4042d2;
      42594: inst = 32'h8220000;
      42595: inst = 32'h10408000;
      42596: inst = 32'hc404338;
      42597: inst = 32'h8220000;
      42598: inst = 32'h10408000;
      42599: inst = 32'hc4043f6;
      42600: inst = 32'h8220000;
      42601: inst = 32'h10408000;
      42602: inst = 32'hc4044b4;
      42603: inst = 32'h8220000;
      42604: inst = 32'h10408000;
      42605: inst = 32'hc404571;
      42606: inst = 32'h8220000;
      42607: inst = 32'h10408000;
      42608: inst = 32'hc404578;
      42609: inst = 32'h8220000;
      42610: inst = 32'h10408000;
      42611: inst = 32'hc404579;
      42612: inst = 32'h8220000;
      42613: inst = 32'hc20be12;
      42614: inst = 32'h10408000;
      42615: inst = 32'hc40428f;
      42616: inst = 32'h8220000;
      42617: inst = 32'hc209db0;
      42618: inst = 32'h10408000;
      42619: inst = 32'hc40429c;
      42620: inst = 32'h8220000;
      42621: inst = 32'hc20cb65;
      42622: inst = 32'h10408000;
      42623: inst = 32'hc4043a4;
      42624: inst = 32'h8220000;
      42625: inst = 32'h10408000;
      42626: inst = 32'hc4043ac;
      42627: inst = 32'h8220000;
      42628: inst = 32'hc20cb43;
      42629: inst = 32'h10408000;
      42630: inst = 32'hc4043a5;
      42631: inst = 32'h8220000;
      42632: inst = 32'h10408000;
      42633: inst = 32'hc405355;
      42634: inst = 32'h8220000;
      42635: inst = 32'h10408000;
      42636: inst = 32'hc405712;
      42637: inst = 32'h8220000;
      42638: inst = 32'hc205bce;
      42639: inst = 32'h10408000;
      42640: inst = 32'hc40466b;
      42641: inst = 32'h8220000;
      42642: inst = 32'h10408000;
      42643: inst = 32'hc404670;
      42644: inst = 32'h8220000;
      42645: inst = 32'h10408000;
      42646: inst = 32'hc404674;
      42647: inst = 32'h8220000;
      42648: inst = 32'h10408000;
      42649: inst = 32'hc4046d2;
      42650: inst = 32'h8220000;
      42651: inst = 32'h10408000;
      42652: inst = 32'hc404735;
      42653: inst = 32'h8220000;
      42654: inst = 32'h10408000;
      42655: inst = 32'hc404739;
      42656: inst = 32'h8220000;
      42657: inst = 32'hc205c2c;
      42658: inst = 32'h10408000;
      42659: inst = 32'hc40466c;
      42660: inst = 32'h8220000;
      42661: inst = 32'hc2063ce;
      42662: inst = 32'h10408000;
      42663: inst = 32'hc404671;
      42664: inst = 32'h8220000;
      42665: inst = 32'hc205bed;
      42666: inst = 32'h10408000;
      42667: inst = 32'hc404672;
      42668: inst = 32'h8220000;
      42669: inst = 32'h10408000;
      42670: inst = 32'hc404678;
      42671: inst = 32'h8220000;
      42672: inst = 32'h10408000;
      42673: inst = 32'hc4046d3;
      42674: inst = 32'h8220000;
      42675: inst = 32'h10408000;
      42676: inst = 32'hc4046d8;
      42677: inst = 32'h8220000;
      42678: inst = 32'h10408000;
      42679: inst = 32'hc404733;
      42680: inst = 32'h8220000;
      42681: inst = 32'hc204c8a;
      42682: inst = 32'h10408000;
      42683: inst = 32'hc4046cb;
      42684: inst = 32'h8220000;
      42685: inst = 32'h10408000;
      42686: inst = 32'hc404734;
      42687: inst = 32'h8220000;
      42688: inst = 32'hc20542c;
      42689: inst = 32'h10408000;
      42690: inst = 32'hc4046d4;
      42691: inst = 32'h8220000;
      42692: inst = 32'h10408000;
      42693: inst = 32'hc40472c;
      42694: inst = 32'h8220000;
      42695: inst = 32'hc205c0d;
      42696: inst = 32'h10408000;
      42697: inst = 32'hc4046d9;
      42698: inst = 32'h8220000;
      42699: inst = 32'h10408000;
      42700: inst = 32'hc404731;
      42701: inst = 32'h8220000;
      42702: inst = 32'hc20e6b5;
      42703: inst = 32'h10408000;
      42704: inst = 32'hc40478b;
      42705: inst = 32'h8220000;
      42706: inst = 32'h10408000;
      42707: inst = 32'hc4048b9;
      42708: inst = 32'h8220000;
      42709: inst = 32'hc20ae51;
      42710: inst = 32'h10408000;
      42711: inst = 32'hc40478c;
      42712: inst = 32'h8220000;
      42713: inst = 32'hc20960e;
      42714: inst = 32'h10408000;
      42715: inst = 32'hc40478d;
      42716: inst = 32'h8220000;
      42717: inst = 32'hc20c673;
      42718: inst = 32'h10408000;
      42719: inst = 32'hc40478e;
      42720: inst = 32'h8220000;
      42721: inst = 32'h10408000;
      42722: inst = 32'hc404793;
      42723: inst = 32'h8220000;
      42724: inst = 32'h10408000;
      42725: inst = 32'hc404854;
      42726: inst = 32'h8220000;
      42727: inst = 32'hc20be52;
      42728: inst = 32'h10408000;
      42729: inst = 32'hc404790;
      42730: inst = 32'h8220000;
      42731: inst = 32'h10408000;
      42732: inst = 32'hc404858;
      42733: inst = 32'h8220000;
      42734: inst = 32'h10408000;
      42735: inst = 32'hc404859;
      42736: inst = 32'h8220000;
      42737: inst = 32'hc209e2f;
      42738: inst = 32'h10408000;
      42739: inst = 32'hc404791;
      42740: inst = 32'h8220000;
      42741: inst = 32'h10408000;
      42742: inst = 32'hc404794;
      42743: inst = 32'h8220000;
      42744: inst = 32'hc20ae30;
      42745: inst = 32'h10408000;
      42746: inst = 32'hc4047ec;
      42747: inst = 32'h8220000;
      42748: inst = 32'h10408000;
      42749: inst = 32'hc4047f1;
      42750: inst = 32'h8220000;
      42751: inst = 32'hc20ce73;
      42752: inst = 32'h10408000;
      42753: inst = 32'hc4047ed;
      42754: inst = 32'h8220000;
      42755: inst = 32'h10408000;
      42756: inst = 32'hc4048b4;
      42757: inst = 32'h8220000;
      42758: inst = 32'hc208e0e;
      42759: inst = 32'h10408000;
      42760: inst = 32'hc4047f0;
      42761: inst = 32'h8220000;
      42762: inst = 32'h10408000;
      42763: inst = 32'hc404855;
      42764: inst = 32'h8220000;
      42765: inst = 32'hc2085ed;
      42766: inst = 32'h10408000;
      42767: inst = 32'hc4047f4;
      42768: inst = 32'h8220000;
      42769: inst = 32'h10408000;
      42770: inst = 32'hc4048b8;
      42771: inst = 32'h8220000;
      42772: inst = 32'hc20b651;
      42773: inst = 32'h10408000;
      42774: inst = 32'hc4047f8;
      42775: inst = 32'h8220000;
      42776: inst = 32'h10408000;
      42777: inst = 32'hc404914;
      42778: inst = 32'h8220000;
      42779: inst = 32'hc20c672;
      42780: inst = 32'h10408000;
      42781: inst = 32'hc4047f9;
      42782: inst = 32'h8220000;
      42783: inst = 32'h10408000;
      42784: inst = 32'hc404856;
      42785: inst = 32'h8220000;
      42786: inst = 32'h10408000;
      42787: inst = 32'hc4048b7;
      42788: inst = 32'h8220000;
      42789: inst = 32'hc209e0f;
      42790: inst = 32'h10408000;
      42791: inst = 32'hc4048b5;
      42792: inst = 32'h8220000;
      42793: inst = 32'h10408000;
      42794: inst = 32'hc404918;
      42795: inst = 32'h8220000;
      42796: inst = 32'hc20de94;
      42797: inst = 32'h10408000;
      42798: inst = 32'hc404917;
      42799: inst = 32'h8220000;
      42800: inst = 32'hc20c2e2;
      42801: inst = 32'h10408000;
      42802: inst = 32'hc405352;
      42803: inst = 32'h8220000;
      42804: inst = 32'hc20cb23;
      42805: inst = 32'h10408000;
      42806: inst = 32'hc405353;
      42807: inst = 32'h8220000;
      42808: inst = 32'h10408000;
      42809: inst = 32'hc405356;
      42810: inst = 32'h8220000;
      42811: inst = 32'h10408000;
      42812: inst = 32'hc405357;
      42813: inst = 32'h8220000;
      42814: inst = 32'h10408000;
      42815: inst = 32'hc405358;
      42816: inst = 32'h8220000;
      42817: inst = 32'h10408000;
      42818: inst = 32'hc405359;
      42819: inst = 32'h8220000;
      42820: inst = 32'h10408000;
      42821: inst = 32'hc40535a;
      42822: inst = 32'h8220000;
      42823: inst = 32'h10408000;
      42824: inst = 32'hc405592;
      42825: inst = 32'h8220000;
      42826: inst = 32'h10408000;
      42827: inst = 32'hc4055f2;
      42828: inst = 32'h8220000;
      42829: inst = 32'h10408000;
      42830: inst = 32'hc405652;
      42831: inst = 32'h8220000;
      42832: inst = 32'h10408000;
      42833: inst = 32'hc4056b2;
      42834: inst = 32'h8220000;
      42835: inst = 32'hc20c323;
      42836: inst = 32'h10408000;
      42837: inst = 32'hc40535b;
      42838: inst = 32'h8220000;
      42839: inst = 32'h10408000;
      42840: inst = 32'hc4057d2;
      42841: inst = 32'h8220000;
      42842: inst = 32'hc20e407;
      42843: inst = 32'h10408000;
      42844: inst = 32'hc4053b3;
      42845: inst = 32'h8220000;
      42846: inst = 32'hc207d9a;
      42847: inst = 32'h10408000;
      42848: inst = 32'hc4053b6;
      42849: inst = 32'h8220000;
      42850: inst = 32'hc2065fe;
      42851: inst = 32'h10408000;
      42852: inst = 32'hc4053b7;
      42853: inst = 32'h8220000;
      42854: inst = 32'hc2065fd;
      42855: inst = 32'h10408000;
      42856: inst = 32'hc4053b8;
      42857: inst = 32'h8220000;
      42858: inst = 32'h10408000;
      42859: inst = 32'hc4053b9;
      42860: inst = 32'h8220000;
      42861: inst = 32'hc20661e;
      42862: inst = 32'h10408000;
      42863: inst = 32'hc4053ba;
      42864: inst = 32'h8220000;
      42865: inst = 32'hc20bb86;
      42866: inst = 32'h10408000;
      42867: inst = 32'hc4053bb;
      42868: inst = 32'h8220000;
      42869: inst = 32'h10408000;
      42870: inst = 32'hc4054db;
      42871: inst = 32'h8220000;
      42872: inst = 32'hc20e6fa;
      42873: inst = 32'h10408000;
      42874: inst = 32'hc4053c9;
      42875: inst = 32'h8220000;
      42876: inst = 32'h10408000;
      42877: inst = 32'hc4053cd;
      42878: inst = 32'h8220000;
      42879: inst = 32'h10408000;
      42880: inst = 32'hc4055a7;
      42881: inst = 32'h8220000;
      42882: inst = 32'hc20e6fb;
      42883: inst = 32'h10408000;
      42884: inst = 32'hc4053ca;
      42885: inst = 32'h8220000;
      42886: inst = 32'h10408000;
      42887: inst = 32'hc4053cc;
      42888: inst = 32'h8220000;
      42889: inst = 32'h10408000;
      42890: inst = 32'hc405487;
      42891: inst = 32'h8220000;
      42892: inst = 32'h10408000;
      42893: inst = 32'hc40548f;
      42894: inst = 32'h8220000;
      42895: inst = 32'h10408000;
      42896: inst = 32'hc405547;
      42897: inst = 32'h8220000;
      42898: inst = 32'h10408000;
      42899: inst = 32'hc40554f;
      42900: inst = 32'h8220000;
      42901: inst = 32'hc20defb;
      42902: inst = 32'h10408000;
      42903: inst = 32'hc4053cb;
      42904: inst = 32'h8220000;
      42905: inst = 32'h10408000;
      42906: inst = 32'hc405428;
      42907: inst = 32'h8220000;
      42908: inst = 32'h10408000;
      42909: inst = 32'hc405429;
      42910: inst = 32'h8220000;
      42911: inst = 32'h10408000;
      42912: inst = 32'hc40542a;
      42913: inst = 32'h8220000;
      42914: inst = 32'h10408000;
      42915: inst = 32'hc40542b;
      42916: inst = 32'h8220000;
      42917: inst = 32'h10408000;
      42918: inst = 32'hc40542c;
      42919: inst = 32'h8220000;
      42920: inst = 32'h10408000;
      42921: inst = 32'hc40542d;
      42922: inst = 32'h8220000;
      42923: inst = 32'h10408000;
      42924: inst = 32'hc40542e;
      42925: inst = 32'h8220000;
      42926: inst = 32'h10408000;
      42927: inst = 32'hc405488;
      42928: inst = 32'h8220000;
      42929: inst = 32'h10408000;
      42930: inst = 32'hc405489;
      42931: inst = 32'h8220000;
      42932: inst = 32'h10408000;
      42933: inst = 32'hc40548a;
      42934: inst = 32'h8220000;
      42935: inst = 32'h10408000;
      42936: inst = 32'hc40548b;
      42937: inst = 32'h8220000;
      42938: inst = 32'h10408000;
      42939: inst = 32'hc40548c;
      42940: inst = 32'h8220000;
      42941: inst = 32'h10408000;
      42942: inst = 32'hc40548d;
      42943: inst = 32'h8220000;
      42944: inst = 32'h10408000;
      42945: inst = 32'hc40548e;
      42946: inst = 32'h8220000;
      42947: inst = 32'h10408000;
      42948: inst = 32'hc4054e7;
      42949: inst = 32'h8220000;
      42950: inst = 32'h10408000;
      42951: inst = 32'hc4054ea;
      42952: inst = 32'h8220000;
      42953: inst = 32'h10408000;
      42954: inst = 32'hc4054ed;
      42955: inst = 32'h8220000;
      42956: inst = 32'h10408000;
      42957: inst = 32'hc4054ee;
      42958: inst = 32'h8220000;
      42959: inst = 32'h10408000;
      42960: inst = 32'hc4054ef;
      42961: inst = 32'h8220000;
      42962: inst = 32'h10408000;
      42963: inst = 32'hc40554a;
      42964: inst = 32'h8220000;
      42965: inst = 32'h10408000;
      42966: inst = 32'hc40554d;
      42967: inst = 32'h8220000;
      42968: inst = 32'h10408000;
      42969: inst = 32'hc40554e;
      42970: inst = 32'h8220000;
      42971: inst = 32'h10408000;
      42972: inst = 32'hc4055a8;
      42973: inst = 32'h8220000;
      42974: inst = 32'h10408000;
      42975: inst = 32'hc4055a9;
      42976: inst = 32'h8220000;
      42977: inst = 32'h10408000;
      42978: inst = 32'hc4055aa;
      42979: inst = 32'h8220000;
      42980: inst = 32'h10408000;
      42981: inst = 32'hc4055ab;
      42982: inst = 32'h8220000;
      42983: inst = 32'h10408000;
      42984: inst = 32'hc4055ac;
      42985: inst = 32'h8220000;
      42986: inst = 32'h10408000;
      42987: inst = 32'hc4055ad;
      42988: inst = 32'h8220000;
      42989: inst = 32'h10408000;
      42990: inst = 32'hc4055ae;
      42991: inst = 32'h8220000;
      42992: inst = 32'h10408000;
      42993: inst = 32'hc405609;
      42994: inst = 32'h8220000;
      42995: inst = 32'h10408000;
      42996: inst = 32'hc40560b;
      42997: inst = 32'h8220000;
      42998: inst = 32'h10408000;
      42999: inst = 32'hc405669;
      43000: inst = 32'h8220000;
      43001: inst = 32'hc20cbc7;
      43002: inst = 32'h10408000;
      43003: inst = 32'hc405412;
      43004: inst = 32'h8220000;
      43005: inst = 32'h10408000;
      43006: inst = 32'hc405472;
      43007: inst = 32'h8220000;
      43008: inst = 32'hc20edb1;
      43009: inst = 32'h10408000;
      43010: inst = 32'hc405413;
      43011: inst = 32'h8220000;
      43012: inst = 32'hc20db43;
      43013: inst = 32'h10408000;
      43014: inst = 32'hc405414;
      43015: inst = 32'h8220000;
      43016: inst = 32'hc207d78;
      43017: inst = 32'h10408000;
      43018: inst = 32'hc405416;
      43019: inst = 32'h8220000;
      43020: inst = 32'hc206dbc;
      43021: inst = 32'h10408000;
      43022: inst = 32'hc405417;
      43023: inst = 32'h8220000;
      43024: inst = 32'h10408000;
      43025: inst = 32'hc405477;
      43026: inst = 32'h8220000;
      43027: inst = 32'hc206dbb;
      43028: inst = 32'h10408000;
      43029: inst = 32'hc405418;
      43030: inst = 32'h8220000;
      43031: inst = 32'h10408000;
      43032: inst = 32'hc405419;
      43033: inst = 32'h8220000;
      43034: inst = 32'h10408000;
      43035: inst = 32'hc405478;
      43036: inst = 32'h8220000;
      43037: inst = 32'h10408000;
      43038: inst = 32'hc405479;
      43039: inst = 32'h8220000;
      43040: inst = 32'hc206ddc;
      43041: inst = 32'h10408000;
      43042: inst = 32'hc40541a;
      43043: inst = 32'h8220000;
      43044: inst = 32'h10408000;
      43045: inst = 32'hc40547a;
      43046: inst = 32'h8220000;
      43047: inst = 32'hc20bb66;
      43048: inst = 32'h10408000;
      43049: inst = 32'hc40541b;
      43050: inst = 32'h8220000;
      43051: inst = 32'h10408000;
      43052: inst = 32'hc40547b;
      43053: inst = 32'h8220000;
      43054: inst = 32'h10408000;
      43055: inst = 32'hc40559b;
      43056: inst = 32'h8220000;
      43057: inst = 32'hc20eed8;
      43058: inst = 32'h10408000;
      43059: inst = 32'hc405427;
      43060: inst = 32'h8220000;
      43061: inst = 32'h10408000;
      43062: inst = 32'hc40542f;
      43063: inst = 32'h8220000;
      43064: inst = 32'hc20edd2;
      43065: inst = 32'h10408000;
      43066: inst = 32'hc405473;
      43067: inst = 32'h8220000;
      43068: inst = 32'hc20db42;
      43069: inst = 32'h10408000;
      43070: inst = 32'hc405474;
      43071: inst = 32'h8220000;
      43072: inst = 32'hc207d79;
      43073: inst = 32'h10408000;
      43074: inst = 32'hc405476;
      43075: inst = 32'h8220000;
      43076: inst = 32'hc20e590;
      43077: inst = 32'h10408000;
      43078: inst = 32'hc4054d3;
      43079: inst = 32'h8220000;
      43080: inst = 32'hc20e363;
      43081: inst = 32'h10408000;
      43082: inst = 32'hc4054d4;
      43083: inst = 32'h8220000;
      43084: inst = 32'hc20d3a6;
      43085: inst = 32'h10408000;
      43086: inst = 32'hc4054d5;
      43087: inst = 32'h8220000;
      43088: inst = 32'hc207dba;
      43089: inst = 32'h10408000;
      43090: inst = 32'hc4054d6;
      43091: inst = 32'h8220000;
      43092: inst = 32'hc2075fd;
      43093: inst = 32'h10408000;
      43094: inst = 32'hc4054d7;
      43095: inst = 32'h8220000;
      43096: inst = 32'h10408000;
      43097: inst = 32'hc4054d8;
      43098: inst = 32'h8220000;
      43099: inst = 32'h10408000;
      43100: inst = 32'hc4054d9;
      43101: inst = 32'h8220000;
      43102: inst = 32'hc206e1e;
      43103: inst = 32'h10408000;
      43104: inst = 32'hc4054da;
      43105: inst = 32'h8220000;
      43106: inst = 32'hc204a69;
      43107: inst = 32'h10408000;
      43108: inst = 32'hc4054e8;
      43109: inst = 32'h8220000;
      43110: inst = 32'h10408000;
      43111: inst = 32'hc4054e9;
      43112: inst = 32'h8220000;
      43113: inst = 32'h10408000;
      43114: inst = 32'hc4054eb;
      43115: inst = 32'h8220000;
      43116: inst = 32'h10408000;
      43117: inst = 32'hc4054ec;
      43118: inst = 32'h8220000;
      43119: inst = 32'h10408000;
      43120: inst = 32'hc405548;
      43121: inst = 32'h8220000;
      43122: inst = 32'h10408000;
      43123: inst = 32'hc405549;
      43124: inst = 32'h8220000;
      43125: inst = 32'h10408000;
      43126: inst = 32'hc40554b;
      43127: inst = 32'h8220000;
      43128: inst = 32'h10408000;
      43129: inst = 32'hc40554c;
      43130: inst = 32'h8220000;
      43131: inst = 32'h10408000;
      43132: inst = 32'hc405608;
      43133: inst = 32'h8220000;
      43134: inst = 32'h10408000;
      43135: inst = 32'hc40560a;
      43136: inst = 32'h8220000;
      43137: inst = 32'h10408000;
      43138: inst = 32'hc40560c;
      43139: inst = 32'h8220000;
      43140: inst = 32'h10408000;
      43141: inst = 32'hc405668;
      43142: inst = 32'h8220000;
      43143: inst = 32'h10408000;
      43144: inst = 32'hc40566a;
      43145: inst = 32'h8220000;
      43146: inst = 32'hc20eba3;
      43147: inst = 32'h10408000;
      43148: inst = 32'hc405535;
      43149: inst = 32'h8220000;
      43150: inst = 32'hc207411;
      43151: inst = 32'h10408000;
      43152: inst = 32'hc405536;
      43153: inst = 32'h8220000;
      43154: inst = 32'hc205bf2;
      43155: inst = 32'h10408000;
      43156: inst = 32'hc405537;
      43157: inst = 32'h8220000;
      43158: inst = 32'h10408000;
      43159: inst = 32'hc40553a;
      43160: inst = 32'h8220000;
      43161: inst = 32'hc205c12;
      43162: inst = 32'h10408000;
      43163: inst = 32'hc405538;
      43164: inst = 32'h8220000;
      43165: inst = 32'h10408000;
      43166: inst = 32'hc405539;
      43167: inst = 32'h8220000;
      43168: inst = 32'h10408000;
      43169: inst = 32'hc4055f9;
      43170: inst = 32'h8220000;
      43171: inst = 32'hc20bb25;
      43172: inst = 32'h10408000;
      43173: inst = 32'hc40553b;
      43174: inst = 32'h8220000;
      43175: inst = 32'h10408000;
      43176: inst = 32'hc4056bb;
      43177: inst = 32'h8220000;
      43178: inst = 32'h10408000;
      43179: inst = 32'hc40571b;
      43180: inst = 32'h8220000;
      43181: inst = 32'h10408000;
      43182: inst = 32'hc40577b;
      43183: inst = 32'h8220000;
      43184: inst = 32'hc20dba4;
      43185: inst = 32'h10408000;
      43186: inst = 32'hc405593;
      43187: inst = 32'h8220000;
      43188: inst = 32'h10408000;
      43189: inst = 32'hc4056b4;
      43190: inst = 32'h8220000;
      43191: inst = 32'hc206288;
      43192: inst = 32'h10408000;
      43193: inst = 32'hc405596;
      43194: inst = 32'h8220000;
      43195: inst = 32'hc205bb1;
      43196: inst = 32'h10408000;
      43197: inst = 32'hc405597;
      43198: inst = 32'h8220000;
      43199: inst = 32'hc2052ec;
      43200: inst = 32'h10408000;
      43201: inst = 32'hc405598;
      43202: inst = 32'h8220000;
      43203: inst = 32'hc20532d;
      43204: inst = 32'h10408000;
      43205: inst = 32'hc405599;
      43206: inst = 32'h8220000;
      43207: inst = 32'hc205390;
      43208: inst = 32'h10408000;
      43209: inst = 32'hc40559a;
      43210: inst = 32'h8220000;
      43211: inst = 32'hc20e6d9;
      43212: inst = 32'h10408000;
      43213: inst = 32'hc4055af;
      43214: inst = 32'h8220000;
      43215: inst = 32'hc2062ea;
      43216: inst = 32'h10408000;
      43217: inst = 32'hc4055f6;
      43218: inst = 32'h8220000;
      43219: inst = 32'hc2064f8;
      43220: inst = 32'h10408000;
      43221: inst = 32'hc4055f7;
      43222: inst = 32'h8220000;
      43223: inst = 32'hc205bd1;
      43224: inst = 32'h10408000;
      43225: inst = 32'hc4055f8;
      43226: inst = 32'h8220000;
      43227: inst = 32'hc2064d6;
      43228: inst = 32'h10408000;
      43229: inst = 32'hc4055fa;
      43230: inst = 32'h8220000;
      43231: inst = 32'hc20bba7;
      43232: inst = 32'h10408000;
      43233: inst = 32'hc4055fb;
      43234: inst = 32'h8220000;
      43235: inst = 32'hc20eeb7;
      43236: inst = 32'h10408000;
      43237: inst = 32'hc405607;
      43238: inst = 32'h8220000;
      43239: inst = 32'hc20d699;
      43240: inst = 32'h10408000;
      43241: inst = 32'hc40560d;
      43242: inst = 32'h8220000;
      43243: inst = 32'hc20b553;
      43244: inst = 32'h10408000;
      43245: inst = 32'hc40560e;
      43246: inst = 32'h8220000;
      43247: inst = 32'hc2083cd;
      43248: inst = 32'h10408000;
      43249: inst = 32'hc40560f;
      43250: inst = 32'h8220000;
      43251: inst = 32'hc20736c;
      43252: inst = 32'h10408000;
      43253: inst = 32'hc405610;
      43254: inst = 32'h8220000;
      43255: inst = 32'hc20a4d0;
      43256: inst = 32'h10408000;
      43257: inst = 32'hc405611;
      43258: inst = 32'h8220000;
      43259: inst = 32'hc20de55;
      43260: inst = 32'h10408000;
      43261: inst = 32'hc405612;
      43262: inst = 32'h8220000;
      43263: inst = 32'hc2062eb;
      43264: inst = 32'h10408000;
      43265: inst = 32'hc405656;
      43266: inst = 32'h8220000;
      43267: inst = 32'hc206496;
      43268: inst = 32'h10408000;
      43269: inst = 32'hc405657;
      43270: inst = 32'h8220000;
      43271: inst = 32'hc205bb0;
      43272: inst = 32'h10408000;
      43273: inst = 32'hc405658;
      43274: inst = 32'h8220000;
      43275: inst = 32'hc2063f2;
      43276: inst = 32'h10408000;
      43277: inst = 32'hc405659;
      43278: inst = 32'h8220000;
      43279: inst = 32'hc206475;
      43280: inst = 32'h10408000;
      43281: inst = 32'hc40565a;
      43282: inst = 32'h8220000;
      43283: inst = 32'hc20bb87;
      43284: inst = 32'h10408000;
      43285: inst = 32'hc40565b;
      43286: inst = 32'h8220000;
      43287: inst = 32'hc209492;
      43288: inst = 32'h10408000;
      43289: inst = 32'hc40566b;
      43290: inst = 32'h8220000;
      43291: inst = 32'hc204228;
      43292: inst = 32'h10408000;
      43293: inst = 32'hc40566c;
      43294: inst = 32'h8220000;
      43295: inst = 32'h10408000;
      43296: inst = 32'hc405760;
      43297: inst = 32'h8220000;
      43298: inst = 32'hc20632c;
      43299: inst = 32'h10408000;
      43300: inst = 32'hc40566d;
      43301: inst = 32'h8220000;
      43302: inst = 32'hc20a4d1;
      43303: inst = 32'h10408000;
      43304: inst = 32'hc40566e;
      43305: inst = 32'h8220000;
      43306: inst = 32'hc20cdf4;
      43307: inst = 32'h10408000;
      43308: inst = 32'hc40566f;
      43309: inst = 32'h8220000;
      43310: inst = 32'hc20c593;
      43311: inst = 32'h10408000;
      43312: inst = 32'hc405670;
      43313: inst = 32'h8220000;
      43314: inst = 32'hc20944f;
      43315: inst = 32'h10408000;
      43316: inst = 32'hc405671;
      43317: inst = 32'h8220000;
      43318: inst = 32'hc20734c;
      43319: inst = 32'h10408000;
      43320: inst = 32'hc405672;
      43321: inst = 32'h8220000;
      43322: inst = 32'hc20a4b0;
      43323: inst = 32'h10408000;
      43324: inst = 32'hc405673;
      43325: inst = 32'h8220000;
      43326: inst = 32'hc20e3e6;
      43327: inst = 32'h10408000;
      43328: inst = 32'hc4056b3;
      43329: inst = 32'h8220000;
      43330: inst = 32'hc209ac5;
      43331: inst = 32'h10408000;
      43332: inst = 32'hc4056b5;
      43333: inst = 32'h8220000;
      43334: inst = 32'hc206350;
      43335: inst = 32'h10408000;
      43336: inst = 32'hc4056ba;
      43337: inst = 32'h8220000;
      43338: inst = 32'h10408000;
      43339: inst = 32'hc40571a;
      43340: inst = 32'h8220000;
      43341: inst = 32'h10408000;
      43342: inst = 32'hc405776;
      43343: inst = 32'h8220000;
      43344: inst = 32'hc2052ac;
      43345: inst = 32'h10408000;
      43346: inst = 32'hc4056ca;
      43347: inst = 32'h8220000;
      43348: inst = 32'h10408000;
      43349: inst = 32'hc4056d0;
      43350: inst = 32'h8220000;
      43351: inst = 32'h10408000;
      43352: inst = 32'hc4057bf;
      43353: inst = 32'h8220000;
      43354: inst = 32'hc204a6a;
      43355: inst = 32'h10408000;
      43356: inst = 32'hc4056cb;
      43357: inst = 32'h8220000;
      43358: inst = 32'h10408000;
      43359: inst = 32'hc4056cc;
      43360: inst = 32'h8220000;
      43361: inst = 32'h10408000;
      43362: inst = 32'hc4056cd;
      43363: inst = 32'h8220000;
      43364: inst = 32'h10408000;
      43365: inst = 32'hc4056ce;
      43366: inst = 32'h8220000;
      43367: inst = 32'h10408000;
      43368: inst = 32'hc4057c0;
      43369: inst = 32'h8220000;
      43370: inst = 32'hc20528b;
      43371: inst = 32'h10408000;
      43372: inst = 32'hc4056cf;
      43373: inst = 32'h8220000;
      43374: inst = 32'hc205acd;
      43375: inst = 32'h10408000;
      43376: inst = 32'hc4056d1;
      43377: inst = 32'h8220000;
      43378: inst = 32'hc205aed;
      43379: inst = 32'h10408000;
      43380: inst = 32'hc4056d2;
      43381: inst = 32'h8220000;
      43382: inst = 32'h10408000;
      43383: inst = 32'hc40575f;
      43384: inst = 32'h8220000;
      43385: inst = 32'hc20632f;
      43386: inst = 32'h10408000;
      43387: inst = 32'hc4056d3;
      43388: inst = 32'h8220000;
      43389: inst = 32'h10408000;
      43390: inst = 32'hc405715;
      43391: inst = 32'h8220000;
      43392: inst = 32'hc20634f;
      43393: inst = 32'h10408000;
      43394: inst = 32'hc4056fe;
      43395: inst = 32'h8220000;
      43396: inst = 32'hc204208;
      43397: inst = 32'h10408000;
      43398: inst = 32'hc4056ff;
      43399: inst = 32'h8220000;
      43400: inst = 32'h10408000;
      43401: inst = 32'hc405700;
      43402: inst = 32'h8220000;
      43403: inst = 32'hc209ae6;
      43404: inst = 32'h10408000;
      43405: inst = 32'hc405714;
      43406: inst = 32'h8220000;
      43407: inst = 32'hc206370;
      43408: inst = 32'h10408000;
      43409: inst = 32'hc405716;
      43410: inst = 32'h8220000;
      43411: inst = 32'h10408000;
      43412: inst = 32'hc405777;
      43413: inst = 32'h8220000;
      43414: inst = 32'h10408000;
      43415: inst = 32'hc405778;
      43416: inst = 32'h8220000;
      43417: inst = 32'h10408000;
      43418: inst = 32'hc405779;
      43419: inst = 32'h8220000;
      43420: inst = 32'hc20c303;
      43421: inst = 32'h10408000;
      43422: inst = 32'hc405772;
      43423: inst = 32'h8220000;
      43424: inst = 32'hc20aaa2;
      43425: inst = 32'h10408000;
      43426: inst = 32'hc405773;
      43427: inst = 32'h8220000;
      43428: inst = 32'hc2072ea;
      43429: inst = 32'h10408000;
      43430: inst = 32'hc405774;
      43431: inst = 32'h8220000;
      43432: inst = 32'hc205b72;
      43433: inst = 32'h10408000;
      43434: inst = 32'hc405775;
      43435: inst = 32'h8220000;
      43436: inst = 32'hc206371;
      43437: inst = 32'h10408000;
      43438: inst = 32'hc40577a;
      43439: inst = 32'h8220000;
      43440: inst = 32'hc20bae3;
      43441: inst = 32'h10408000;
      43442: inst = 32'hc4057d3;
      43443: inst = 32'h8220000;
      43444: inst = 32'hc20bb04;
      43445: inst = 32'h10408000;
      43446: inst = 32'hc4057d4;
      43447: inst = 32'h8220000;
      43448: inst = 32'hc20b325;
      43449: inst = 32'h10408000;
      43450: inst = 32'hc4057d5;
      43451: inst = 32'h8220000;
      43452: inst = 32'h10408000;
      43453: inst = 32'hc4057d6;
      43454: inst = 32'h8220000;
      43455: inst = 32'h10408000;
      43456: inst = 32'hc4057d7;
      43457: inst = 32'h8220000;
      43458: inst = 32'h10408000;
      43459: inst = 32'hc4057d8;
      43460: inst = 32'h8220000;
      43461: inst = 32'h10408000;
      43462: inst = 32'hc4057d9;
      43463: inst = 32'h8220000;
      43464: inst = 32'h10408000;
      43465: inst = 32'hc4057da;
      43466: inst = 32'h8220000;
      43467: inst = 32'hc20c344;
      43468: inst = 32'h10408000;
      43469: inst = 32'hc4057db;
      43470: inst = 32'h8220000;
      43471: inst = 32'h58000000;
      43472: inst = 32'h11800000;
      43473: inst = 32'hd800000;
      43474: inst = 32'h11a00000;
      43475: inst = 32'hda00000;
      43476: inst = 32'h25ad5800;
      43477: inst = 32'h15ca6800;
      43478: inst = 32'h21c00001;
      43479: inst = 32'h59200000;
      43480: inst = 32'h298c0001;
      43481: inst = 32'h13e00000;
      43482: inst = 32'hfe0a9d4;
      43483: inst = 32'h5be00000;
      43484: inst = 32'h11800000;
      43485: inst = 32'hd800000;
      43486: inst = 32'h258c5800;
      43487: inst = 32'h15aa6000;
      43488: inst = 32'h13e00000;
      43489: inst = 32'hfe0a9e7;
      43490: inst = 32'h21a00001;
      43491: inst = 32'h5be00000;
      43492: inst = 32'h13e00000;
      43493: inst = 32'hfe0a9de;
      43494: inst = 32'h5be00000;
      43495: inst = 32'h2d8c5800;
      43496: inst = 32'h2d8a6000;
      43497: inst = 32'h59200000;
      43498: inst = 32'h11800000;
      43499: inst = 32'hd800000;
      43500: inst = 32'h29ab0000;
      43501: inst = 32'h31ad0001;
      43502: inst = 32'h258c5000;
      43503: inst = 32'h21a00000;
      43504: inst = 32'h59200000;
      43505: inst = 32'h13e00000;
      43506: inst = 32'hfe0a9ed;
      43507: inst = 32'h5be00000;
      43508: inst = 32'h10608000;
      43509: inst = 32'hc600000;
      43510: inst = 32'hc20aaaa;
      43511: inst = 32'h4c210000;
      43512: inst = 32'h8230000;
      43513: inst = 32'h104000fe;
      43514: inst = 32'hc40502a;
      43515: inst = 32'h30420001;
      43516: inst = 32'h13e00000;
      43517: inst = 32'hfe0a9fb;
      43518: inst = 32'h1c400000;
      43519: inst = 32'h5be00000;
      43520: inst = 32'h13e00000;
      43521: inst = 32'hfe0a9f7;
      43522: inst = 32'h5be00000;
    endcase
  end
endmodule
