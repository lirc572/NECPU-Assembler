`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Company: lirc572
// Engineer: lirc572
// 
// Create Date: 
// Design Name: NECPU
// Module Name: InstMem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module instMem (
    input  [31:0]  address,
    output reg [31:0] inst
  );
  always @ (address) begin
    inst = 32'd0;
    case (address)
      0: inst = 32'h10000000;
      1: inst = 32'hc000005;
      2: inst = 32'h13e00000;
      3: inst = 32'hfe000b6;
      4: inst = 32'h5be00000;
      5: inst = 32'h1020007f;
      6: inst = 32'hc202815;
      7: inst = 32'h30210001;
      8: inst = 32'h13e00000;
      9: inst = 32'hfe00007;
      10: inst = 32'h1c200000;
      11: inst = 32'h5be00000;
      12: inst = 32'h10000000;
      13: inst = 32'hc000011;
      14: inst = 32'h13e00000;
      15: inst = 32'hfe0490e;
      16: inst = 32'h5be00000;
      17: inst = 32'h1020007f;
      18: inst = 32'hc202815;
      19: inst = 32'h30210001;
      20: inst = 32'h13e00000;
      21: inst = 32'hfe00013;
      22: inst = 32'h1c200000;
      23: inst = 32'h5be00000;
      24: inst = 32'h10000000;
      25: inst = 32'hc000000;
      26: inst = 32'h10200000;
      27: inst = 32'hc20001f;
      28: inst = 32'h13e00000;
      29: inst = 32'hfe06127;
      30: inst = 32'h5be00000;
      31: inst = 32'h10000000;
      32: inst = 32'hc000024;
      33: inst = 32'h13a00000;
      34: inst = 32'hfa00000;
      35: inst = 32'h13600000;
      36: inst = 32'hf600000;
      37: inst = 32'h13800000;
      38: inst = 32'hf800000;
      39: inst = 32'h12800000;
      40: inst = 32'he800045;
      41: inst = 32'h12a00000;
      42: inst = 32'hea0002b;
      43: inst = 32'h1734d800;
      44: inst = 32'h1755e000;
      45: inst = 32'h13e00000;
      46: inst = 32'hfe00038;
      47: inst = 32'h1f200001;
      48: inst = 32'h5be00000;
      49: inst = 32'h13e00000;
      50: inst = 32'hfe00038;
      51: inst = 32'h1f400001;
      52: inst = 32'h5be00000;
      53: inst = 32'h13e00000;
      54: inst = 32'hfe000a6;
      55: inst = 32'h5be00000;
      56: inst = 32'h12800000;
      57: inst = 32'he80000e;
      58: inst = 32'h12a00000;
      59: inst = 32'hea0002b;
      60: inst = 32'h173ba000;
      61: inst = 32'h1755e000;
      62: inst = 32'h13e00000;
      63: inst = 32'hfe00049;
      64: inst = 32'h1f200001;
      65: inst = 32'h5be00000;
      66: inst = 32'h13e00000;
      67: inst = 32'hfe00049;
      68: inst = 32'h1f400001;
      69: inst = 32'h5be00000;
      70: inst = 32'h13e00000;
      71: inst = 32'hfe000ae;
      72: inst = 32'h5be00000;
      73: inst = 32'h10208000;
      74: inst = 32'hc200001;
      75: inst = 32'h4210000;
      76: inst = 32'h10400000;
      77: inst = 32'hc40001b;
      78: inst = 32'h34211000;
      79: inst = 32'h38211000;
      80: inst = 32'h13e00000;
      81: inst = 32'hfe00063;
      82: inst = 32'h20200010;
      83: inst = 32'h5be00000;
      84: inst = 32'h13e00000;
      85: inst = 32'hfe0006d;
      86: inst = 32'h20200008;
      87: inst = 32'h5be00000;
      88: inst = 32'h13e00000;
      89: inst = 32'hfe00077;
      90: inst = 32'h20200004;
      91: inst = 32'h5be00000;
      92: inst = 32'h13e00000;
      93: inst = 32'hfe00081;
      94: inst = 32'h20200002;
      95: inst = 32'h5be00000;
      96: inst = 32'h13e00000;
      97: inst = 32'hfe0008b;
      98: inst = 32'h5be00000;
      99: inst = 32'h2b9c0001;
      100: inst = 32'h13a00000;
      101: inst = 32'hfa00000;
      102: inst = 32'hca00001;
      103: inst = 32'h10c08000;
      104: inst = 32'hcc00000;
      105: inst = 32'h8a60000;
      106: inst = 32'h13e00000;
      107: inst = 32'hfe0008f;
      108: inst = 32'h5be00000;
      109: inst = 32'h2b7b0001;
      110: inst = 32'h13a00000;
      111: inst = 32'hfa00003;
      112: inst = 32'hca00002;
      113: inst = 32'h10c08000;
      114: inst = 32'hcc00000;
      115: inst = 32'h8a60000;
      116: inst = 32'h13e00000;
      117: inst = 32'hfe0008f;
      118: inst = 32'h5be00000;
      119: inst = 32'h337b0001;
      120: inst = 32'h13a00000;
      121: inst = 32'hfa00001;
      122: inst = 32'hca00004;
      123: inst = 32'h10c08000;
      124: inst = 32'hcc00000;
      125: inst = 32'h8a60000;
      126: inst = 32'h13e00000;
      127: inst = 32'hfe0008f;
      128: inst = 32'h5be00000;
      129: inst = 32'h339c0001;
      130: inst = 32'h13a00000;
      131: inst = 32'hfa00005;
      132: inst = 32'hca00008;
      133: inst = 32'h10c08000;
      134: inst = 32'hcc00000;
      135: inst = 32'h8a60000;
      136: inst = 32'h13e00000;
      137: inst = 32'hfe0008f;
      138: inst = 32'h5be00000;
      139: inst = 32'hca00010;
      140: inst = 32'h10c08000;
      141: inst = 32'hcc00000;
      142: inst = 32'h8a60000;
      143: inst = 32'h10000000;
      144: inst = 32'hc000094;
      145: inst = 32'h13e00000;
      146: inst = 32'hfe06131;
      147: inst = 32'h5be00000;
      148: inst = 32'h283d0000;
      149: inst = 32'h285b0000;
      150: inst = 32'h287c0000;
      151: inst = 32'h10000000;
      152: inst = 32'hc00009c;
      153: inst = 32'h13e00000;
      154: inst = 32'hfe0515f;
      155: inst = 32'h5be00000;
      156: inst = 32'h10200007;
      157: inst = 32'hc20a120;
      158: inst = 32'h30210001;
      159: inst = 32'h13e00000;
      160: inst = 32'hfe0009e;
      161: inst = 32'h1c200000;
      162: inst = 32'h5be00000;
      163: inst = 32'h13e00000;
      164: inst = 32'hfe00027;
      165: inst = 32'h5be00000;
      166: inst = 32'h10000000;
      167: inst = 32'hc0000ab;
      168: inst = 32'h13e00000;
      169: inst = 32'hfe0aa23;
      170: inst = 32'h5be00000;
      171: inst = 32'h13e00000;
      172: inst = 32'hfe0b093;
      173: inst = 32'h5be00000;
      174: inst = 32'h10000000;
      175: inst = 32'hc0000b3;
      176: inst = 32'h13e00000;
      177: inst = 32'hfe0aecc;
      178: inst = 32'h5be00000;
      179: inst = 32'h13e00000;
      180: inst = 32'hfe0b093;
      181: inst = 32'h5be00000;
      182: inst = 32'hc20eeb6;
      183: inst = 32'h10408000;
      184: inst = 32'hc403fe0;
      185: inst = 32'h8220000;
      186: inst = 32'h10408000;
      187: inst = 32'hc403fe1;
      188: inst = 32'h8220000;
      189: inst = 32'h10408000;
      190: inst = 32'hc403fe2;
      191: inst = 32'h8220000;
      192: inst = 32'h10408000;
      193: inst = 32'hc403fe3;
      194: inst = 32'h8220000;
      195: inst = 32'h10408000;
      196: inst = 32'hc403fe4;
      197: inst = 32'h8220000;
      198: inst = 32'h10408000;
      199: inst = 32'hc403fe5;
      200: inst = 32'h8220000;
      201: inst = 32'h10408000;
      202: inst = 32'hc403fe6;
      203: inst = 32'h8220000;
      204: inst = 32'h10408000;
      205: inst = 32'hc403fe7;
      206: inst = 32'h8220000;
      207: inst = 32'h10408000;
      208: inst = 32'hc403fe8;
      209: inst = 32'h8220000;
      210: inst = 32'h10408000;
      211: inst = 32'hc403fe9;
      212: inst = 32'h8220000;
      213: inst = 32'h10408000;
      214: inst = 32'hc403fea;
      215: inst = 32'h8220000;
      216: inst = 32'h10408000;
      217: inst = 32'hc403fec;
      218: inst = 32'h8220000;
      219: inst = 32'h10408000;
      220: inst = 32'hc403fed;
      221: inst = 32'h8220000;
      222: inst = 32'h10408000;
      223: inst = 32'hc403fee;
      224: inst = 32'h8220000;
      225: inst = 32'h10408000;
      226: inst = 32'hc403fef;
      227: inst = 32'h8220000;
      228: inst = 32'h10408000;
      229: inst = 32'hc403ff0;
      230: inst = 32'h8220000;
      231: inst = 32'h10408000;
      232: inst = 32'hc403ff1;
      233: inst = 32'h8220000;
      234: inst = 32'h10408000;
      235: inst = 32'hc403ff2;
      236: inst = 32'h8220000;
      237: inst = 32'h10408000;
      238: inst = 32'hc403ff3;
      239: inst = 32'h8220000;
      240: inst = 32'h10408000;
      241: inst = 32'hc403ff4;
      242: inst = 32'h8220000;
      243: inst = 32'h10408000;
      244: inst = 32'hc403ff5;
      245: inst = 32'h8220000;
      246: inst = 32'h10408000;
      247: inst = 32'hc403ff6;
      248: inst = 32'h8220000;
      249: inst = 32'h10408000;
      250: inst = 32'hc403ff7;
      251: inst = 32'h8220000;
      252: inst = 32'h10408000;
      253: inst = 32'hc403ff8;
      254: inst = 32'h8220000;
      255: inst = 32'h10408000;
      256: inst = 32'hc403ff9;
      257: inst = 32'h8220000;
      258: inst = 32'h10408000;
      259: inst = 32'hc403ffa;
      260: inst = 32'h8220000;
      261: inst = 32'h10408000;
      262: inst = 32'hc403ffb;
      263: inst = 32'h8220000;
      264: inst = 32'h10408000;
      265: inst = 32'hc403ffc;
      266: inst = 32'h8220000;
      267: inst = 32'h10408000;
      268: inst = 32'hc403ffd;
      269: inst = 32'h8220000;
      270: inst = 32'h10408000;
      271: inst = 32'hc403ffe;
      272: inst = 32'h8220000;
      273: inst = 32'h10408000;
      274: inst = 32'hc403fff;
      275: inst = 32'h8220000;
      276: inst = 32'h10408000;
      277: inst = 32'hc404000;
      278: inst = 32'h8220000;
      279: inst = 32'h10408000;
      280: inst = 32'hc404001;
      281: inst = 32'h8220000;
      282: inst = 32'h10408000;
      283: inst = 32'hc404002;
      284: inst = 32'h8220000;
      285: inst = 32'h10408000;
      286: inst = 32'hc404003;
      287: inst = 32'h8220000;
      288: inst = 32'h10408000;
      289: inst = 32'hc404004;
      290: inst = 32'h8220000;
      291: inst = 32'h10408000;
      292: inst = 32'hc404005;
      293: inst = 32'h8220000;
      294: inst = 32'h10408000;
      295: inst = 32'hc404006;
      296: inst = 32'h8220000;
      297: inst = 32'h10408000;
      298: inst = 32'hc404007;
      299: inst = 32'h8220000;
      300: inst = 32'h10408000;
      301: inst = 32'hc404008;
      302: inst = 32'h8220000;
      303: inst = 32'h10408000;
      304: inst = 32'hc404009;
      305: inst = 32'h8220000;
      306: inst = 32'h10408000;
      307: inst = 32'hc40400a;
      308: inst = 32'h8220000;
      309: inst = 32'h10408000;
      310: inst = 32'hc40400b;
      311: inst = 32'h8220000;
      312: inst = 32'h10408000;
      313: inst = 32'hc40400c;
      314: inst = 32'h8220000;
      315: inst = 32'h10408000;
      316: inst = 32'hc40400d;
      317: inst = 32'h8220000;
      318: inst = 32'h10408000;
      319: inst = 32'hc40400e;
      320: inst = 32'h8220000;
      321: inst = 32'h10408000;
      322: inst = 32'hc40400f;
      323: inst = 32'h8220000;
      324: inst = 32'h10408000;
      325: inst = 32'hc404010;
      326: inst = 32'h8220000;
      327: inst = 32'h10408000;
      328: inst = 32'hc404011;
      329: inst = 32'h8220000;
      330: inst = 32'h10408000;
      331: inst = 32'hc404012;
      332: inst = 32'h8220000;
      333: inst = 32'h10408000;
      334: inst = 32'hc404013;
      335: inst = 32'h8220000;
      336: inst = 32'h10408000;
      337: inst = 32'hc404014;
      338: inst = 32'h8220000;
      339: inst = 32'h10408000;
      340: inst = 32'hc404015;
      341: inst = 32'h8220000;
      342: inst = 32'h10408000;
      343: inst = 32'hc404016;
      344: inst = 32'h8220000;
      345: inst = 32'h10408000;
      346: inst = 32'hc404017;
      347: inst = 32'h8220000;
      348: inst = 32'h10408000;
      349: inst = 32'hc404018;
      350: inst = 32'h8220000;
      351: inst = 32'h10408000;
      352: inst = 32'hc404019;
      353: inst = 32'h8220000;
      354: inst = 32'h10408000;
      355: inst = 32'hc40401a;
      356: inst = 32'h8220000;
      357: inst = 32'h10408000;
      358: inst = 32'hc40401b;
      359: inst = 32'h8220000;
      360: inst = 32'h10408000;
      361: inst = 32'hc40401c;
      362: inst = 32'h8220000;
      363: inst = 32'h10408000;
      364: inst = 32'hc40401d;
      365: inst = 32'h8220000;
      366: inst = 32'h10408000;
      367: inst = 32'hc40401e;
      368: inst = 32'h8220000;
      369: inst = 32'h10408000;
      370: inst = 32'hc40401f;
      371: inst = 32'h8220000;
      372: inst = 32'h10408000;
      373: inst = 32'hc404020;
      374: inst = 32'h8220000;
      375: inst = 32'h10408000;
      376: inst = 32'hc404021;
      377: inst = 32'h8220000;
      378: inst = 32'h10408000;
      379: inst = 32'hc404022;
      380: inst = 32'h8220000;
      381: inst = 32'h10408000;
      382: inst = 32'hc404023;
      383: inst = 32'h8220000;
      384: inst = 32'h10408000;
      385: inst = 32'hc404024;
      386: inst = 32'h8220000;
      387: inst = 32'h10408000;
      388: inst = 32'hc404025;
      389: inst = 32'h8220000;
      390: inst = 32'h10408000;
      391: inst = 32'hc404026;
      392: inst = 32'h8220000;
      393: inst = 32'h10408000;
      394: inst = 32'hc404027;
      395: inst = 32'h8220000;
      396: inst = 32'h10408000;
      397: inst = 32'hc404028;
      398: inst = 32'h8220000;
      399: inst = 32'h10408000;
      400: inst = 32'hc404029;
      401: inst = 32'h8220000;
      402: inst = 32'h10408000;
      403: inst = 32'hc40402a;
      404: inst = 32'h8220000;
      405: inst = 32'h10408000;
      406: inst = 32'hc40402b;
      407: inst = 32'h8220000;
      408: inst = 32'h10408000;
      409: inst = 32'hc40402c;
      410: inst = 32'h8220000;
      411: inst = 32'h10408000;
      412: inst = 32'hc40402d;
      413: inst = 32'h8220000;
      414: inst = 32'h10408000;
      415: inst = 32'hc40402e;
      416: inst = 32'h8220000;
      417: inst = 32'h10408000;
      418: inst = 32'hc40402f;
      419: inst = 32'h8220000;
      420: inst = 32'h10408000;
      421: inst = 32'hc404030;
      422: inst = 32'h8220000;
      423: inst = 32'h10408000;
      424: inst = 32'hc404031;
      425: inst = 32'h8220000;
      426: inst = 32'h10408000;
      427: inst = 32'hc404032;
      428: inst = 32'h8220000;
      429: inst = 32'h10408000;
      430: inst = 32'hc404033;
      431: inst = 32'h8220000;
      432: inst = 32'h10408000;
      433: inst = 32'hc404034;
      434: inst = 32'h8220000;
      435: inst = 32'h10408000;
      436: inst = 32'hc404035;
      437: inst = 32'h8220000;
      438: inst = 32'h10408000;
      439: inst = 32'hc404036;
      440: inst = 32'h8220000;
      441: inst = 32'h10408000;
      442: inst = 32'hc404037;
      443: inst = 32'h8220000;
      444: inst = 32'h10408000;
      445: inst = 32'hc404038;
      446: inst = 32'h8220000;
      447: inst = 32'h10408000;
      448: inst = 32'hc404039;
      449: inst = 32'h8220000;
      450: inst = 32'h10408000;
      451: inst = 32'hc40403a;
      452: inst = 32'h8220000;
      453: inst = 32'h10408000;
      454: inst = 32'hc40403b;
      455: inst = 32'h8220000;
      456: inst = 32'h10408000;
      457: inst = 32'hc40403c;
      458: inst = 32'h8220000;
      459: inst = 32'h10408000;
      460: inst = 32'hc40403d;
      461: inst = 32'h8220000;
      462: inst = 32'h10408000;
      463: inst = 32'hc40403e;
      464: inst = 32'h8220000;
      465: inst = 32'h10408000;
      466: inst = 32'hc40403f;
      467: inst = 32'h8220000;
      468: inst = 32'h10408000;
      469: inst = 32'hc404040;
      470: inst = 32'h8220000;
      471: inst = 32'h10408000;
      472: inst = 32'hc404041;
      473: inst = 32'h8220000;
      474: inst = 32'h10408000;
      475: inst = 32'hc404042;
      476: inst = 32'h8220000;
      477: inst = 32'h10408000;
      478: inst = 32'hc404043;
      479: inst = 32'h8220000;
      480: inst = 32'h10408000;
      481: inst = 32'hc404044;
      482: inst = 32'h8220000;
      483: inst = 32'h10408000;
      484: inst = 32'hc404045;
      485: inst = 32'h8220000;
      486: inst = 32'h10408000;
      487: inst = 32'hc404046;
      488: inst = 32'h8220000;
      489: inst = 32'h10408000;
      490: inst = 32'hc404047;
      491: inst = 32'h8220000;
      492: inst = 32'h10408000;
      493: inst = 32'hc404048;
      494: inst = 32'h8220000;
      495: inst = 32'h10408000;
      496: inst = 32'hc404049;
      497: inst = 32'h8220000;
      498: inst = 32'h10408000;
      499: inst = 32'hc40404a;
      500: inst = 32'h8220000;
      501: inst = 32'h10408000;
      502: inst = 32'hc40404c;
      503: inst = 32'h8220000;
      504: inst = 32'h10408000;
      505: inst = 32'hc40404d;
      506: inst = 32'h8220000;
      507: inst = 32'h10408000;
      508: inst = 32'hc40404e;
      509: inst = 32'h8220000;
      510: inst = 32'h10408000;
      511: inst = 32'hc40404f;
      512: inst = 32'h8220000;
      513: inst = 32'h10408000;
      514: inst = 32'hc404050;
      515: inst = 32'h8220000;
      516: inst = 32'h10408000;
      517: inst = 32'hc404051;
      518: inst = 32'h8220000;
      519: inst = 32'h10408000;
      520: inst = 32'hc404052;
      521: inst = 32'h8220000;
      522: inst = 32'h10408000;
      523: inst = 32'hc404053;
      524: inst = 32'h8220000;
      525: inst = 32'h10408000;
      526: inst = 32'hc404054;
      527: inst = 32'h8220000;
      528: inst = 32'h10408000;
      529: inst = 32'hc404055;
      530: inst = 32'h8220000;
      531: inst = 32'h10408000;
      532: inst = 32'hc404056;
      533: inst = 32'h8220000;
      534: inst = 32'h10408000;
      535: inst = 32'hc404057;
      536: inst = 32'h8220000;
      537: inst = 32'h10408000;
      538: inst = 32'hc404058;
      539: inst = 32'h8220000;
      540: inst = 32'h10408000;
      541: inst = 32'hc404059;
      542: inst = 32'h8220000;
      543: inst = 32'h10408000;
      544: inst = 32'hc40405a;
      545: inst = 32'h8220000;
      546: inst = 32'h10408000;
      547: inst = 32'hc40405b;
      548: inst = 32'h8220000;
      549: inst = 32'h10408000;
      550: inst = 32'hc40405c;
      551: inst = 32'h8220000;
      552: inst = 32'h10408000;
      553: inst = 32'hc40405d;
      554: inst = 32'h8220000;
      555: inst = 32'h10408000;
      556: inst = 32'hc40405e;
      557: inst = 32'h8220000;
      558: inst = 32'h10408000;
      559: inst = 32'hc40405f;
      560: inst = 32'h8220000;
      561: inst = 32'h10408000;
      562: inst = 32'hc404060;
      563: inst = 32'h8220000;
      564: inst = 32'h10408000;
      565: inst = 32'hc404061;
      566: inst = 32'h8220000;
      567: inst = 32'h10408000;
      568: inst = 32'hc404062;
      569: inst = 32'h8220000;
      570: inst = 32'h10408000;
      571: inst = 32'hc404063;
      572: inst = 32'h8220000;
      573: inst = 32'h10408000;
      574: inst = 32'hc404064;
      575: inst = 32'h8220000;
      576: inst = 32'h10408000;
      577: inst = 32'hc404065;
      578: inst = 32'h8220000;
      579: inst = 32'h10408000;
      580: inst = 32'hc404066;
      581: inst = 32'h8220000;
      582: inst = 32'h10408000;
      583: inst = 32'hc404067;
      584: inst = 32'h8220000;
      585: inst = 32'h10408000;
      586: inst = 32'hc404068;
      587: inst = 32'h8220000;
      588: inst = 32'h10408000;
      589: inst = 32'hc404069;
      590: inst = 32'h8220000;
      591: inst = 32'h10408000;
      592: inst = 32'hc40406a;
      593: inst = 32'h8220000;
      594: inst = 32'h10408000;
      595: inst = 32'hc40406b;
      596: inst = 32'h8220000;
      597: inst = 32'h10408000;
      598: inst = 32'hc40406c;
      599: inst = 32'h8220000;
      600: inst = 32'h10408000;
      601: inst = 32'hc40406d;
      602: inst = 32'h8220000;
      603: inst = 32'h10408000;
      604: inst = 32'hc40406e;
      605: inst = 32'h8220000;
      606: inst = 32'h10408000;
      607: inst = 32'hc40406f;
      608: inst = 32'h8220000;
      609: inst = 32'h10408000;
      610: inst = 32'hc404070;
      611: inst = 32'h8220000;
      612: inst = 32'h10408000;
      613: inst = 32'hc404071;
      614: inst = 32'h8220000;
      615: inst = 32'h10408000;
      616: inst = 32'hc404072;
      617: inst = 32'h8220000;
      618: inst = 32'h10408000;
      619: inst = 32'hc404073;
      620: inst = 32'h8220000;
      621: inst = 32'h10408000;
      622: inst = 32'hc404074;
      623: inst = 32'h8220000;
      624: inst = 32'h10408000;
      625: inst = 32'hc404075;
      626: inst = 32'h8220000;
      627: inst = 32'h10408000;
      628: inst = 32'hc404076;
      629: inst = 32'h8220000;
      630: inst = 32'h10408000;
      631: inst = 32'hc404077;
      632: inst = 32'h8220000;
      633: inst = 32'h10408000;
      634: inst = 32'hc404078;
      635: inst = 32'h8220000;
      636: inst = 32'h10408000;
      637: inst = 32'hc404079;
      638: inst = 32'h8220000;
      639: inst = 32'h10408000;
      640: inst = 32'hc40407a;
      641: inst = 32'h8220000;
      642: inst = 32'h10408000;
      643: inst = 32'hc40407b;
      644: inst = 32'h8220000;
      645: inst = 32'h10408000;
      646: inst = 32'hc40407c;
      647: inst = 32'h8220000;
      648: inst = 32'h10408000;
      649: inst = 32'hc40407d;
      650: inst = 32'h8220000;
      651: inst = 32'h10408000;
      652: inst = 32'hc40407e;
      653: inst = 32'h8220000;
      654: inst = 32'h10408000;
      655: inst = 32'hc40407f;
      656: inst = 32'h8220000;
      657: inst = 32'h10408000;
      658: inst = 32'hc404080;
      659: inst = 32'h8220000;
      660: inst = 32'h10408000;
      661: inst = 32'hc404081;
      662: inst = 32'h8220000;
      663: inst = 32'h10408000;
      664: inst = 32'hc404082;
      665: inst = 32'h8220000;
      666: inst = 32'h10408000;
      667: inst = 32'hc404083;
      668: inst = 32'h8220000;
      669: inst = 32'h10408000;
      670: inst = 32'hc404084;
      671: inst = 32'h8220000;
      672: inst = 32'h10408000;
      673: inst = 32'hc404085;
      674: inst = 32'h8220000;
      675: inst = 32'h10408000;
      676: inst = 32'hc404086;
      677: inst = 32'h8220000;
      678: inst = 32'h10408000;
      679: inst = 32'hc404087;
      680: inst = 32'h8220000;
      681: inst = 32'h10408000;
      682: inst = 32'hc404088;
      683: inst = 32'h8220000;
      684: inst = 32'h10408000;
      685: inst = 32'hc404089;
      686: inst = 32'h8220000;
      687: inst = 32'h10408000;
      688: inst = 32'hc40408a;
      689: inst = 32'h8220000;
      690: inst = 32'h10408000;
      691: inst = 32'hc40408b;
      692: inst = 32'h8220000;
      693: inst = 32'h10408000;
      694: inst = 32'hc40408c;
      695: inst = 32'h8220000;
      696: inst = 32'h10408000;
      697: inst = 32'hc40408d;
      698: inst = 32'h8220000;
      699: inst = 32'h10408000;
      700: inst = 32'hc40408e;
      701: inst = 32'h8220000;
      702: inst = 32'h10408000;
      703: inst = 32'hc40408f;
      704: inst = 32'h8220000;
      705: inst = 32'h10408000;
      706: inst = 32'hc404090;
      707: inst = 32'h8220000;
      708: inst = 32'h10408000;
      709: inst = 32'hc404091;
      710: inst = 32'h8220000;
      711: inst = 32'h10408000;
      712: inst = 32'hc404092;
      713: inst = 32'h8220000;
      714: inst = 32'h10408000;
      715: inst = 32'hc404093;
      716: inst = 32'h8220000;
      717: inst = 32'h10408000;
      718: inst = 32'hc404094;
      719: inst = 32'h8220000;
      720: inst = 32'h10408000;
      721: inst = 32'hc404095;
      722: inst = 32'h8220000;
      723: inst = 32'h10408000;
      724: inst = 32'hc404096;
      725: inst = 32'h8220000;
      726: inst = 32'h10408000;
      727: inst = 32'hc404097;
      728: inst = 32'h8220000;
      729: inst = 32'h10408000;
      730: inst = 32'hc404098;
      731: inst = 32'h8220000;
      732: inst = 32'h10408000;
      733: inst = 32'hc404099;
      734: inst = 32'h8220000;
      735: inst = 32'h10408000;
      736: inst = 32'hc40409a;
      737: inst = 32'h8220000;
      738: inst = 32'h10408000;
      739: inst = 32'hc40409b;
      740: inst = 32'h8220000;
      741: inst = 32'h10408000;
      742: inst = 32'hc40409c;
      743: inst = 32'h8220000;
      744: inst = 32'h10408000;
      745: inst = 32'hc40409d;
      746: inst = 32'h8220000;
      747: inst = 32'h10408000;
      748: inst = 32'hc40409e;
      749: inst = 32'h8220000;
      750: inst = 32'h10408000;
      751: inst = 32'hc40409f;
      752: inst = 32'h8220000;
      753: inst = 32'h10408000;
      754: inst = 32'hc4040a0;
      755: inst = 32'h8220000;
      756: inst = 32'h10408000;
      757: inst = 32'hc4040a1;
      758: inst = 32'h8220000;
      759: inst = 32'h10408000;
      760: inst = 32'hc4040a2;
      761: inst = 32'h8220000;
      762: inst = 32'h10408000;
      763: inst = 32'hc4040a3;
      764: inst = 32'h8220000;
      765: inst = 32'h10408000;
      766: inst = 32'hc4040a4;
      767: inst = 32'h8220000;
      768: inst = 32'h10408000;
      769: inst = 32'hc4040a5;
      770: inst = 32'h8220000;
      771: inst = 32'h10408000;
      772: inst = 32'hc4040a6;
      773: inst = 32'h8220000;
      774: inst = 32'h10408000;
      775: inst = 32'hc4040a7;
      776: inst = 32'h8220000;
      777: inst = 32'h10408000;
      778: inst = 32'hc4040a8;
      779: inst = 32'h8220000;
      780: inst = 32'h10408000;
      781: inst = 32'hc4040a9;
      782: inst = 32'h8220000;
      783: inst = 32'h10408000;
      784: inst = 32'hc4040aa;
      785: inst = 32'h8220000;
      786: inst = 32'h10408000;
      787: inst = 32'hc4040ac;
      788: inst = 32'h8220000;
      789: inst = 32'h10408000;
      790: inst = 32'hc4040ad;
      791: inst = 32'h8220000;
      792: inst = 32'h10408000;
      793: inst = 32'hc4040ae;
      794: inst = 32'h8220000;
      795: inst = 32'h10408000;
      796: inst = 32'hc4040af;
      797: inst = 32'h8220000;
      798: inst = 32'h10408000;
      799: inst = 32'hc4040b0;
      800: inst = 32'h8220000;
      801: inst = 32'h10408000;
      802: inst = 32'hc4040b1;
      803: inst = 32'h8220000;
      804: inst = 32'h10408000;
      805: inst = 32'hc4040b2;
      806: inst = 32'h8220000;
      807: inst = 32'h10408000;
      808: inst = 32'hc4040b3;
      809: inst = 32'h8220000;
      810: inst = 32'h10408000;
      811: inst = 32'hc4040b4;
      812: inst = 32'h8220000;
      813: inst = 32'h10408000;
      814: inst = 32'hc4040b5;
      815: inst = 32'h8220000;
      816: inst = 32'h10408000;
      817: inst = 32'hc4040b6;
      818: inst = 32'h8220000;
      819: inst = 32'h10408000;
      820: inst = 32'hc4040b7;
      821: inst = 32'h8220000;
      822: inst = 32'h10408000;
      823: inst = 32'hc4040b8;
      824: inst = 32'h8220000;
      825: inst = 32'h10408000;
      826: inst = 32'hc4040b9;
      827: inst = 32'h8220000;
      828: inst = 32'h10408000;
      829: inst = 32'hc4040ba;
      830: inst = 32'h8220000;
      831: inst = 32'h10408000;
      832: inst = 32'hc4040bb;
      833: inst = 32'h8220000;
      834: inst = 32'h10408000;
      835: inst = 32'hc4040bc;
      836: inst = 32'h8220000;
      837: inst = 32'h10408000;
      838: inst = 32'hc4040bd;
      839: inst = 32'h8220000;
      840: inst = 32'h10408000;
      841: inst = 32'hc4040be;
      842: inst = 32'h8220000;
      843: inst = 32'h10408000;
      844: inst = 32'hc4040bf;
      845: inst = 32'h8220000;
      846: inst = 32'h10408000;
      847: inst = 32'hc4040c0;
      848: inst = 32'h8220000;
      849: inst = 32'h10408000;
      850: inst = 32'hc4040c1;
      851: inst = 32'h8220000;
      852: inst = 32'h10408000;
      853: inst = 32'hc4040c2;
      854: inst = 32'h8220000;
      855: inst = 32'h10408000;
      856: inst = 32'hc4040c3;
      857: inst = 32'h8220000;
      858: inst = 32'h10408000;
      859: inst = 32'hc4040c4;
      860: inst = 32'h8220000;
      861: inst = 32'h10408000;
      862: inst = 32'hc4040c5;
      863: inst = 32'h8220000;
      864: inst = 32'h10408000;
      865: inst = 32'hc4040c6;
      866: inst = 32'h8220000;
      867: inst = 32'h10408000;
      868: inst = 32'hc4040c7;
      869: inst = 32'h8220000;
      870: inst = 32'h10408000;
      871: inst = 32'hc4040c8;
      872: inst = 32'h8220000;
      873: inst = 32'h10408000;
      874: inst = 32'hc4040c9;
      875: inst = 32'h8220000;
      876: inst = 32'h10408000;
      877: inst = 32'hc4040ca;
      878: inst = 32'h8220000;
      879: inst = 32'h10408000;
      880: inst = 32'hc4040cb;
      881: inst = 32'h8220000;
      882: inst = 32'h10408000;
      883: inst = 32'hc4040cc;
      884: inst = 32'h8220000;
      885: inst = 32'h10408000;
      886: inst = 32'hc4040cd;
      887: inst = 32'h8220000;
      888: inst = 32'h10408000;
      889: inst = 32'hc4040ce;
      890: inst = 32'h8220000;
      891: inst = 32'h10408000;
      892: inst = 32'hc4040cf;
      893: inst = 32'h8220000;
      894: inst = 32'h10408000;
      895: inst = 32'hc4040d0;
      896: inst = 32'h8220000;
      897: inst = 32'h10408000;
      898: inst = 32'hc4040d1;
      899: inst = 32'h8220000;
      900: inst = 32'h10408000;
      901: inst = 32'hc4040d2;
      902: inst = 32'h8220000;
      903: inst = 32'h10408000;
      904: inst = 32'hc4040d3;
      905: inst = 32'h8220000;
      906: inst = 32'h10408000;
      907: inst = 32'hc4040d4;
      908: inst = 32'h8220000;
      909: inst = 32'h10408000;
      910: inst = 32'hc4040d5;
      911: inst = 32'h8220000;
      912: inst = 32'h10408000;
      913: inst = 32'hc4040d6;
      914: inst = 32'h8220000;
      915: inst = 32'h10408000;
      916: inst = 32'hc4040d7;
      917: inst = 32'h8220000;
      918: inst = 32'h10408000;
      919: inst = 32'hc4040d8;
      920: inst = 32'h8220000;
      921: inst = 32'h10408000;
      922: inst = 32'hc4040d9;
      923: inst = 32'h8220000;
      924: inst = 32'h10408000;
      925: inst = 32'hc4040da;
      926: inst = 32'h8220000;
      927: inst = 32'h10408000;
      928: inst = 32'hc4040db;
      929: inst = 32'h8220000;
      930: inst = 32'h10408000;
      931: inst = 32'hc4040dc;
      932: inst = 32'h8220000;
      933: inst = 32'h10408000;
      934: inst = 32'hc4040dd;
      935: inst = 32'h8220000;
      936: inst = 32'h10408000;
      937: inst = 32'hc4040de;
      938: inst = 32'h8220000;
      939: inst = 32'h10408000;
      940: inst = 32'hc4040df;
      941: inst = 32'h8220000;
      942: inst = 32'h10408000;
      943: inst = 32'hc4040e0;
      944: inst = 32'h8220000;
      945: inst = 32'h10408000;
      946: inst = 32'hc4040e1;
      947: inst = 32'h8220000;
      948: inst = 32'h10408000;
      949: inst = 32'hc4040e2;
      950: inst = 32'h8220000;
      951: inst = 32'h10408000;
      952: inst = 32'hc4040e3;
      953: inst = 32'h8220000;
      954: inst = 32'h10408000;
      955: inst = 32'hc4040e4;
      956: inst = 32'h8220000;
      957: inst = 32'h10408000;
      958: inst = 32'hc4040e5;
      959: inst = 32'h8220000;
      960: inst = 32'h10408000;
      961: inst = 32'hc4040e6;
      962: inst = 32'h8220000;
      963: inst = 32'h10408000;
      964: inst = 32'hc4040e7;
      965: inst = 32'h8220000;
      966: inst = 32'h10408000;
      967: inst = 32'hc4040e8;
      968: inst = 32'h8220000;
      969: inst = 32'h10408000;
      970: inst = 32'hc4040e9;
      971: inst = 32'h8220000;
      972: inst = 32'h10408000;
      973: inst = 32'hc4040ea;
      974: inst = 32'h8220000;
      975: inst = 32'h10408000;
      976: inst = 32'hc4040eb;
      977: inst = 32'h8220000;
      978: inst = 32'h10408000;
      979: inst = 32'hc4040ec;
      980: inst = 32'h8220000;
      981: inst = 32'h10408000;
      982: inst = 32'hc4040ed;
      983: inst = 32'h8220000;
      984: inst = 32'h10408000;
      985: inst = 32'hc4040ee;
      986: inst = 32'h8220000;
      987: inst = 32'h10408000;
      988: inst = 32'hc4040ef;
      989: inst = 32'h8220000;
      990: inst = 32'h10408000;
      991: inst = 32'hc4040f0;
      992: inst = 32'h8220000;
      993: inst = 32'h10408000;
      994: inst = 32'hc4040f1;
      995: inst = 32'h8220000;
      996: inst = 32'h10408000;
      997: inst = 32'hc4040f2;
      998: inst = 32'h8220000;
      999: inst = 32'h10408000;
      1000: inst = 32'hc4040f3;
      1001: inst = 32'h8220000;
      1002: inst = 32'h10408000;
      1003: inst = 32'hc4040f4;
      1004: inst = 32'h8220000;
      1005: inst = 32'h10408000;
      1006: inst = 32'hc4040f5;
      1007: inst = 32'h8220000;
      1008: inst = 32'h10408000;
      1009: inst = 32'hc4040f6;
      1010: inst = 32'h8220000;
      1011: inst = 32'h10408000;
      1012: inst = 32'hc4040f7;
      1013: inst = 32'h8220000;
      1014: inst = 32'h10408000;
      1015: inst = 32'hc4040f8;
      1016: inst = 32'h8220000;
      1017: inst = 32'h10408000;
      1018: inst = 32'hc4040f9;
      1019: inst = 32'h8220000;
      1020: inst = 32'h10408000;
      1021: inst = 32'hc4040fa;
      1022: inst = 32'h8220000;
      1023: inst = 32'h10408000;
      1024: inst = 32'hc4040fb;
      1025: inst = 32'h8220000;
      1026: inst = 32'h10408000;
      1027: inst = 32'hc4040fc;
      1028: inst = 32'h8220000;
      1029: inst = 32'h10408000;
      1030: inst = 32'hc4040fd;
      1031: inst = 32'h8220000;
      1032: inst = 32'h10408000;
      1033: inst = 32'hc4040fe;
      1034: inst = 32'h8220000;
      1035: inst = 32'h10408000;
      1036: inst = 32'hc4040ff;
      1037: inst = 32'h8220000;
      1038: inst = 32'h10408000;
      1039: inst = 32'hc404100;
      1040: inst = 32'h8220000;
      1041: inst = 32'h10408000;
      1042: inst = 32'hc404101;
      1043: inst = 32'h8220000;
      1044: inst = 32'h10408000;
      1045: inst = 32'hc404102;
      1046: inst = 32'h8220000;
      1047: inst = 32'h10408000;
      1048: inst = 32'hc404103;
      1049: inst = 32'h8220000;
      1050: inst = 32'h10408000;
      1051: inst = 32'hc404104;
      1052: inst = 32'h8220000;
      1053: inst = 32'h10408000;
      1054: inst = 32'hc404105;
      1055: inst = 32'h8220000;
      1056: inst = 32'h10408000;
      1057: inst = 32'hc404106;
      1058: inst = 32'h8220000;
      1059: inst = 32'h10408000;
      1060: inst = 32'hc404107;
      1061: inst = 32'h8220000;
      1062: inst = 32'h10408000;
      1063: inst = 32'hc404108;
      1064: inst = 32'h8220000;
      1065: inst = 32'h10408000;
      1066: inst = 32'hc404109;
      1067: inst = 32'h8220000;
      1068: inst = 32'h10408000;
      1069: inst = 32'hc40410a;
      1070: inst = 32'h8220000;
      1071: inst = 32'h10408000;
      1072: inst = 32'hc40410c;
      1073: inst = 32'h8220000;
      1074: inst = 32'h10408000;
      1075: inst = 32'hc40410d;
      1076: inst = 32'h8220000;
      1077: inst = 32'h10408000;
      1078: inst = 32'hc40410e;
      1079: inst = 32'h8220000;
      1080: inst = 32'h10408000;
      1081: inst = 32'hc40410f;
      1082: inst = 32'h8220000;
      1083: inst = 32'h10408000;
      1084: inst = 32'hc404110;
      1085: inst = 32'h8220000;
      1086: inst = 32'h10408000;
      1087: inst = 32'hc404111;
      1088: inst = 32'h8220000;
      1089: inst = 32'h10408000;
      1090: inst = 32'hc404112;
      1091: inst = 32'h8220000;
      1092: inst = 32'h10408000;
      1093: inst = 32'hc404113;
      1094: inst = 32'h8220000;
      1095: inst = 32'h10408000;
      1096: inst = 32'hc404114;
      1097: inst = 32'h8220000;
      1098: inst = 32'h10408000;
      1099: inst = 32'hc404115;
      1100: inst = 32'h8220000;
      1101: inst = 32'h10408000;
      1102: inst = 32'hc404116;
      1103: inst = 32'h8220000;
      1104: inst = 32'h10408000;
      1105: inst = 32'hc404117;
      1106: inst = 32'h8220000;
      1107: inst = 32'h10408000;
      1108: inst = 32'hc404118;
      1109: inst = 32'h8220000;
      1110: inst = 32'h10408000;
      1111: inst = 32'hc404119;
      1112: inst = 32'h8220000;
      1113: inst = 32'h10408000;
      1114: inst = 32'hc40411a;
      1115: inst = 32'h8220000;
      1116: inst = 32'h10408000;
      1117: inst = 32'hc40411b;
      1118: inst = 32'h8220000;
      1119: inst = 32'h10408000;
      1120: inst = 32'hc40411c;
      1121: inst = 32'h8220000;
      1122: inst = 32'h10408000;
      1123: inst = 32'hc40411d;
      1124: inst = 32'h8220000;
      1125: inst = 32'h10408000;
      1126: inst = 32'hc40411e;
      1127: inst = 32'h8220000;
      1128: inst = 32'h10408000;
      1129: inst = 32'hc40411f;
      1130: inst = 32'h8220000;
      1131: inst = 32'h10408000;
      1132: inst = 32'hc404120;
      1133: inst = 32'h8220000;
      1134: inst = 32'h10408000;
      1135: inst = 32'hc404121;
      1136: inst = 32'h8220000;
      1137: inst = 32'h10408000;
      1138: inst = 32'hc404122;
      1139: inst = 32'h8220000;
      1140: inst = 32'h10408000;
      1141: inst = 32'hc404123;
      1142: inst = 32'h8220000;
      1143: inst = 32'h10408000;
      1144: inst = 32'hc404124;
      1145: inst = 32'h8220000;
      1146: inst = 32'h10408000;
      1147: inst = 32'hc404125;
      1148: inst = 32'h8220000;
      1149: inst = 32'h10408000;
      1150: inst = 32'hc404126;
      1151: inst = 32'h8220000;
      1152: inst = 32'h10408000;
      1153: inst = 32'hc404127;
      1154: inst = 32'h8220000;
      1155: inst = 32'h10408000;
      1156: inst = 32'hc404128;
      1157: inst = 32'h8220000;
      1158: inst = 32'h10408000;
      1159: inst = 32'hc404129;
      1160: inst = 32'h8220000;
      1161: inst = 32'h10408000;
      1162: inst = 32'hc40412a;
      1163: inst = 32'h8220000;
      1164: inst = 32'h10408000;
      1165: inst = 32'hc40412b;
      1166: inst = 32'h8220000;
      1167: inst = 32'h10408000;
      1168: inst = 32'hc40412c;
      1169: inst = 32'h8220000;
      1170: inst = 32'h10408000;
      1171: inst = 32'hc40412d;
      1172: inst = 32'h8220000;
      1173: inst = 32'h10408000;
      1174: inst = 32'hc40412e;
      1175: inst = 32'h8220000;
      1176: inst = 32'h10408000;
      1177: inst = 32'hc40412f;
      1178: inst = 32'h8220000;
      1179: inst = 32'h10408000;
      1180: inst = 32'hc404130;
      1181: inst = 32'h8220000;
      1182: inst = 32'h10408000;
      1183: inst = 32'hc404131;
      1184: inst = 32'h8220000;
      1185: inst = 32'h10408000;
      1186: inst = 32'hc404132;
      1187: inst = 32'h8220000;
      1188: inst = 32'h10408000;
      1189: inst = 32'hc404133;
      1190: inst = 32'h8220000;
      1191: inst = 32'h10408000;
      1192: inst = 32'hc404134;
      1193: inst = 32'h8220000;
      1194: inst = 32'h10408000;
      1195: inst = 32'hc404135;
      1196: inst = 32'h8220000;
      1197: inst = 32'h10408000;
      1198: inst = 32'hc404136;
      1199: inst = 32'h8220000;
      1200: inst = 32'h10408000;
      1201: inst = 32'hc404137;
      1202: inst = 32'h8220000;
      1203: inst = 32'h10408000;
      1204: inst = 32'hc404138;
      1205: inst = 32'h8220000;
      1206: inst = 32'h10408000;
      1207: inst = 32'hc404139;
      1208: inst = 32'h8220000;
      1209: inst = 32'h10408000;
      1210: inst = 32'hc40413a;
      1211: inst = 32'h8220000;
      1212: inst = 32'h10408000;
      1213: inst = 32'hc40413b;
      1214: inst = 32'h8220000;
      1215: inst = 32'h10408000;
      1216: inst = 32'hc40413c;
      1217: inst = 32'h8220000;
      1218: inst = 32'h10408000;
      1219: inst = 32'hc40413d;
      1220: inst = 32'h8220000;
      1221: inst = 32'h10408000;
      1222: inst = 32'hc40413e;
      1223: inst = 32'h8220000;
      1224: inst = 32'h10408000;
      1225: inst = 32'hc40413f;
      1226: inst = 32'h8220000;
      1227: inst = 32'h10408000;
      1228: inst = 32'hc404140;
      1229: inst = 32'h8220000;
      1230: inst = 32'h10408000;
      1231: inst = 32'hc404141;
      1232: inst = 32'h8220000;
      1233: inst = 32'h10408000;
      1234: inst = 32'hc404142;
      1235: inst = 32'h8220000;
      1236: inst = 32'h10408000;
      1237: inst = 32'hc404143;
      1238: inst = 32'h8220000;
      1239: inst = 32'h10408000;
      1240: inst = 32'hc404144;
      1241: inst = 32'h8220000;
      1242: inst = 32'h10408000;
      1243: inst = 32'hc404145;
      1244: inst = 32'h8220000;
      1245: inst = 32'h10408000;
      1246: inst = 32'hc404146;
      1247: inst = 32'h8220000;
      1248: inst = 32'h10408000;
      1249: inst = 32'hc404147;
      1250: inst = 32'h8220000;
      1251: inst = 32'h10408000;
      1252: inst = 32'hc404148;
      1253: inst = 32'h8220000;
      1254: inst = 32'h10408000;
      1255: inst = 32'hc404149;
      1256: inst = 32'h8220000;
      1257: inst = 32'h10408000;
      1258: inst = 32'hc40414a;
      1259: inst = 32'h8220000;
      1260: inst = 32'h10408000;
      1261: inst = 32'hc40414b;
      1262: inst = 32'h8220000;
      1263: inst = 32'h10408000;
      1264: inst = 32'hc40414c;
      1265: inst = 32'h8220000;
      1266: inst = 32'h10408000;
      1267: inst = 32'hc40414d;
      1268: inst = 32'h8220000;
      1269: inst = 32'h10408000;
      1270: inst = 32'hc40414e;
      1271: inst = 32'h8220000;
      1272: inst = 32'h10408000;
      1273: inst = 32'hc40414f;
      1274: inst = 32'h8220000;
      1275: inst = 32'h10408000;
      1276: inst = 32'hc404150;
      1277: inst = 32'h8220000;
      1278: inst = 32'h10408000;
      1279: inst = 32'hc404151;
      1280: inst = 32'h8220000;
      1281: inst = 32'h10408000;
      1282: inst = 32'hc404152;
      1283: inst = 32'h8220000;
      1284: inst = 32'h10408000;
      1285: inst = 32'hc404153;
      1286: inst = 32'h8220000;
      1287: inst = 32'h10408000;
      1288: inst = 32'hc404154;
      1289: inst = 32'h8220000;
      1290: inst = 32'h10408000;
      1291: inst = 32'hc404155;
      1292: inst = 32'h8220000;
      1293: inst = 32'h10408000;
      1294: inst = 32'hc404156;
      1295: inst = 32'h8220000;
      1296: inst = 32'h10408000;
      1297: inst = 32'hc404157;
      1298: inst = 32'h8220000;
      1299: inst = 32'h10408000;
      1300: inst = 32'hc404158;
      1301: inst = 32'h8220000;
      1302: inst = 32'h10408000;
      1303: inst = 32'hc404159;
      1304: inst = 32'h8220000;
      1305: inst = 32'h10408000;
      1306: inst = 32'hc40415a;
      1307: inst = 32'h8220000;
      1308: inst = 32'h10408000;
      1309: inst = 32'hc40415b;
      1310: inst = 32'h8220000;
      1311: inst = 32'h10408000;
      1312: inst = 32'hc40415c;
      1313: inst = 32'h8220000;
      1314: inst = 32'h10408000;
      1315: inst = 32'hc40415d;
      1316: inst = 32'h8220000;
      1317: inst = 32'h10408000;
      1318: inst = 32'hc40415e;
      1319: inst = 32'h8220000;
      1320: inst = 32'h10408000;
      1321: inst = 32'hc40415f;
      1322: inst = 32'h8220000;
      1323: inst = 32'h10408000;
      1324: inst = 32'hc404160;
      1325: inst = 32'h8220000;
      1326: inst = 32'h10408000;
      1327: inst = 32'hc404161;
      1328: inst = 32'h8220000;
      1329: inst = 32'h10408000;
      1330: inst = 32'hc404162;
      1331: inst = 32'h8220000;
      1332: inst = 32'h10408000;
      1333: inst = 32'hc404163;
      1334: inst = 32'h8220000;
      1335: inst = 32'h10408000;
      1336: inst = 32'hc404164;
      1337: inst = 32'h8220000;
      1338: inst = 32'h10408000;
      1339: inst = 32'hc404165;
      1340: inst = 32'h8220000;
      1341: inst = 32'h10408000;
      1342: inst = 32'hc404166;
      1343: inst = 32'h8220000;
      1344: inst = 32'h10408000;
      1345: inst = 32'hc404167;
      1346: inst = 32'h8220000;
      1347: inst = 32'h10408000;
      1348: inst = 32'hc404168;
      1349: inst = 32'h8220000;
      1350: inst = 32'h10408000;
      1351: inst = 32'hc404169;
      1352: inst = 32'h8220000;
      1353: inst = 32'h10408000;
      1354: inst = 32'hc40416a;
      1355: inst = 32'h8220000;
      1356: inst = 32'h10408000;
      1357: inst = 32'hc40416c;
      1358: inst = 32'h8220000;
      1359: inst = 32'h10408000;
      1360: inst = 32'hc40416d;
      1361: inst = 32'h8220000;
      1362: inst = 32'h10408000;
      1363: inst = 32'hc40416e;
      1364: inst = 32'h8220000;
      1365: inst = 32'h10408000;
      1366: inst = 32'hc40416f;
      1367: inst = 32'h8220000;
      1368: inst = 32'h10408000;
      1369: inst = 32'hc404170;
      1370: inst = 32'h8220000;
      1371: inst = 32'h10408000;
      1372: inst = 32'hc404171;
      1373: inst = 32'h8220000;
      1374: inst = 32'h10408000;
      1375: inst = 32'hc404172;
      1376: inst = 32'h8220000;
      1377: inst = 32'h10408000;
      1378: inst = 32'hc404173;
      1379: inst = 32'h8220000;
      1380: inst = 32'h10408000;
      1381: inst = 32'hc404174;
      1382: inst = 32'h8220000;
      1383: inst = 32'h10408000;
      1384: inst = 32'hc404175;
      1385: inst = 32'h8220000;
      1386: inst = 32'h10408000;
      1387: inst = 32'hc404176;
      1388: inst = 32'h8220000;
      1389: inst = 32'h10408000;
      1390: inst = 32'hc404177;
      1391: inst = 32'h8220000;
      1392: inst = 32'h10408000;
      1393: inst = 32'hc404178;
      1394: inst = 32'h8220000;
      1395: inst = 32'h10408000;
      1396: inst = 32'hc404179;
      1397: inst = 32'h8220000;
      1398: inst = 32'h10408000;
      1399: inst = 32'hc40417a;
      1400: inst = 32'h8220000;
      1401: inst = 32'h10408000;
      1402: inst = 32'hc40417b;
      1403: inst = 32'h8220000;
      1404: inst = 32'h10408000;
      1405: inst = 32'hc40417c;
      1406: inst = 32'h8220000;
      1407: inst = 32'h10408000;
      1408: inst = 32'hc40417d;
      1409: inst = 32'h8220000;
      1410: inst = 32'h10408000;
      1411: inst = 32'hc40417e;
      1412: inst = 32'h8220000;
      1413: inst = 32'h10408000;
      1414: inst = 32'hc40417f;
      1415: inst = 32'h8220000;
      1416: inst = 32'h10408000;
      1417: inst = 32'hc404180;
      1418: inst = 32'h8220000;
      1419: inst = 32'h10408000;
      1420: inst = 32'hc404181;
      1421: inst = 32'h8220000;
      1422: inst = 32'h10408000;
      1423: inst = 32'hc404182;
      1424: inst = 32'h8220000;
      1425: inst = 32'h10408000;
      1426: inst = 32'hc404183;
      1427: inst = 32'h8220000;
      1428: inst = 32'h10408000;
      1429: inst = 32'hc404184;
      1430: inst = 32'h8220000;
      1431: inst = 32'h10408000;
      1432: inst = 32'hc404185;
      1433: inst = 32'h8220000;
      1434: inst = 32'h10408000;
      1435: inst = 32'hc404186;
      1436: inst = 32'h8220000;
      1437: inst = 32'h10408000;
      1438: inst = 32'hc404187;
      1439: inst = 32'h8220000;
      1440: inst = 32'h10408000;
      1441: inst = 32'hc404188;
      1442: inst = 32'h8220000;
      1443: inst = 32'h10408000;
      1444: inst = 32'hc404189;
      1445: inst = 32'h8220000;
      1446: inst = 32'h10408000;
      1447: inst = 32'hc40418a;
      1448: inst = 32'h8220000;
      1449: inst = 32'h10408000;
      1450: inst = 32'hc40418b;
      1451: inst = 32'h8220000;
      1452: inst = 32'h10408000;
      1453: inst = 32'hc40418c;
      1454: inst = 32'h8220000;
      1455: inst = 32'h10408000;
      1456: inst = 32'hc40418d;
      1457: inst = 32'h8220000;
      1458: inst = 32'h10408000;
      1459: inst = 32'hc40418e;
      1460: inst = 32'h8220000;
      1461: inst = 32'h10408000;
      1462: inst = 32'hc40418f;
      1463: inst = 32'h8220000;
      1464: inst = 32'h10408000;
      1465: inst = 32'hc404190;
      1466: inst = 32'h8220000;
      1467: inst = 32'h10408000;
      1468: inst = 32'hc404191;
      1469: inst = 32'h8220000;
      1470: inst = 32'h10408000;
      1471: inst = 32'hc404192;
      1472: inst = 32'h8220000;
      1473: inst = 32'h10408000;
      1474: inst = 32'hc404193;
      1475: inst = 32'h8220000;
      1476: inst = 32'h10408000;
      1477: inst = 32'hc404194;
      1478: inst = 32'h8220000;
      1479: inst = 32'h10408000;
      1480: inst = 32'hc404195;
      1481: inst = 32'h8220000;
      1482: inst = 32'h10408000;
      1483: inst = 32'hc404196;
      1484: inst = 32'h8220000;
      1485: inst = 32'h10408000;
      1486: inst = 32'hc404197;
      1487: inst = 32'h8220000;
      1488: inst = 32'h10408000;
      1489: inst = 32'hc404198;
      1490: inst = 32'h8220000;
      1491: inst = 32'h10408000;
      1492: inst = 32'hc404199;
      1493: inst = 32'h8220000;
      1494: inst = 32'h10408000;
      1495: inst = 32'hc40419a;
      1496: inst = 32'h8220000;
      1497: inst = 32'h10408000;
      1498: inst = 32'hc40419b;
      1499: inst = 32'h8220000;
      1500: inst = 32'h10408000;
      1501: inst = 32'hc40419c;
      1502: inst = 32'h8220000;
      1503: inst = 32'h10408000;
      1504: inst = 32'hc40419d;
      1505: inst = 32'h8220000;
      1506: inst = 32'h10408000;
      1507: inst = 32'hc40419e;
      1508: inst = 32'h8220000;
      1509: inst = 32'h10408000;
      1510: inst = 32'hc40419f;
      1511: inst = 32'h8220000;
      1512: inst = 32'h10408000;
      1513: inst = 32'hc4041a0;
      1514: inst = 32'h8220000;
      1515: inst = 32'h10408000;
      1516: inst = 32'hc4041a1;
      1517: inst = 32'h8220000;
      1518: inst = 32'h10408000;
      1519: inst = 32'hc4041a2;
      1520: inst = 32'h8220000;
      1521: inst = 32'h10408000;
      1522: inst = 32'hc4041a3;
      1523: inst = 32'h8220000;
      1524: inst = 32'h10408000;
      1525: inst = 32'hc4041a4;
      1526: inst = 32'h8220000;
      1527: inst = 32'h10408000;
      1528: inst = 32'hc4041a5;
      1529: inst = 32'h8220000;
      1530: inst = 32'h10408000;
      1531: inst = 32'hc4041a6;
      1532: inst = 32'h8220000;
      1533: inst = 32'h10408000;
      1534: inst = 32'hc4041a7;
      1535: inst = 32'h8220000;
      1536: inst = 32'h10408000;
      1537: inst = 32'hc4041a8;
      1538: inst = 32'h8220000;
      1539: inst = 32'h10408000;
      1540: inst = 32'hc4041a9;
      1541: inst = 32'h8220000;
      1542: inst = 32'h10408000;
      1543: inst = 32'hc4041aa;
      1544: inst = 32'h8220000;
      1545: inst = 32'h10408000;
      1546: inst = 32'hc4041ab;
      1547: inst = 32'h8220000;
      1548: inst = 32'h10408000;
      1549: inst = 32'hc4041ac;
      1550: inst = 32'h8220000;
      1551: inst = 32'h10408000;
      1552: inst = 32'hc4041ad;
      1553: inst = 32'h8220000;
      1554: inst = 32'h10408000;
      1555: inst = 32'hc4041ae;
      1556: inst = 32'h8220000;
      1557: inst = 32'h10408000;
      1558: inst = 32'hc4041af;
      1559: inst = 32'h8220000;
      1560: inst = 32'h10408000;
      1561: inst = 32'hc4041b0;
      1562: inst = 32'h8220000;
      1563: inst = 32'h10408000;
      1564: inst = 32'hc4041b1;
      1565: inst = 32'h8220000;
      1566: inst = 32'h10408000;
      1567: inst = 32'hc4041b2;
      1568: inst = 32'h8220000;
      1569: inst = 32'h10408000;
      1570: inst = 32'hc4041b3;
      1571: inst = 32'h8220000;
      1572: inst = 32'h10408000;
      1573: inst = 32'hc4041b4;
      1574: inst = 32'h8220000;
      1575: inst = 32'h10408000;
      1576: inst = 32'hc4041b5;
      1577: inst = 32'h8220000;
      1578: inst = 32'h10408000;
      1579: inst = 32'hc4041b6;
      1580: inst = 32'h8220000;
      1581: inst = 32'h10408000;
      1582: inst = 32'hc4041b7;
      1583: inst = 32'h8220000;
      1584: inst = 32'h10408000;
      1585: inst = 32'hc4041b8;
      1586: inst = 32'h8220000;
      1587: inst = 32'h10408000;
      1588: inst = 32'hc4041b9;
      1589: inst = 32'h8220000;
      1590: inst = 32'h10408000;
      1591: inst = 32'hc4041ba;
      1592: inst = 32'h8220000;
      1593: inst = 32'h10408000;
      1594: inst = 32'hc4041bb;
      1595: inst = 32'h8220000;
      1596: inst = 32'h10408000;
      1597: inst = 32'hc4041bc;
      1598: inst = 32'h8220000;
      1599: inst = 32'h10408000;
      1600: inst = 32'hc4041bd;
      1601: inst = 32'h8220000;
      1602: inst = 32'h10408000;
      1603: inst = 32'hc4041be;
      1604: inst = 32'h8220000;
      1605: inst = 32'h10408000;
      1606: inst = 32'hc4041bf;
      1607: inst = 32'h8220000;
      1608: inst = 32'h10408000;
      1609: inst = 32'hc4041c0;
      1610: inst = 32'h8220000;
      1611: inst = 32'h10408000;
      1612: inst = 32'hc4041c1;
      1613: inst = 32'h8220000;
      1614: inst = 32'h10408000;
      1615: inst = 32'hc4041c2;
      1616: inst = 32'h8220000;
      1617: inst = 32'h10408000;
      1618: inst = 32'hc4041c3;
      1619: inst = 32'h8220000;
      1620: inst = 32'h10408000;
      1621: inst = 32'hc4041c4;
      1622: inst = 32'h8220000;
      1623: inst = 32'h10408000;
      1624: inst = 32'hc4041c5;
      1625: inst = 32'h8220000;
      1626: inst = 32'h10408000;
      1627: inst = 32'hc4041c6;
      1628: inst = 32'h8220000;
      1629: inst = 32'h10408000;
      1630: inst = 32'hc4041c7;
      1631: inst = 32'h8220000;
      1632: inst = 32'h10408000;
      1633: inst = 32'hc4041c8;
      1634: inst = 32'h8220000;
      1635: inst = 32'h10408000;
      1636: inst = 32'hc4041c9;
      1637: inst = 32'h8220000;
      1638: inst = 32'h10408000;
      1639: inst = 32'hc4041ca;
      1640: inst = 32'h8220000;
      1641: inst = 32'h10408000;
      1642: inst = 32'hc4041cc;
      1643: inst = 32'h8220000;
      1644: inst = 32'h10408000;
      1645: inst = 32'hc4041cd;
      1646: inst = 32'h8220000;
      1647: inst = 32'h10408000;
      1648: inst = 32'hc4041ce;
      1649: inst = 32'h8220000;
      1650: inst = 32'h10408000;
      1651: inst = 32'hc4041cf;
      1652: inst = 32'h8220000;
      1653: inst = 32'h10408000;
      1654: inst = 32'hc4041d0;
      1655: inst = 32'h8220000;
      1656: inst = 32'h10408000;
      1657: inst = 32'hc4041d1;
      1658: inst = 32'h8220000;
      1659: inst = 32'h10408000;
      1660: inst = 32'hc4041d2;
      1661: inst = 32'h8220000;
      1662: inst = 32'h10408000;
      1663: inst = 32'hc4041d3;
      1664: inst = 32'h8220000;
      1665: inst = 32'h10408000;
      1666: inst = 32'hc4041d4;
      1667: inst = 32'h8220000;
      1668: inst = 32'h10408000;
      1669: inst = 32'hc4041d5;
      1670: inst = 32'h8220000;
      1671: inst = 32'h10408000;
      1672: inst = 32'hc4041d6;
      1673: inst = 32'h8220000;
      1674: inst = 32'h10408000;
      1675: inst = 32'hc4041d7;
      1676: inst = 32'h8220000;
      1677: inst = 32'h10408000;
      1678: inst = 32'hc4041d8;
      1679: inst = 32'h8220000;
      1680: inst = 32'h10408000;
      1681: inst = 32'hc4041d9;
      1682: inst = 32'h8220000;
      1683: inst = 32'h10408000;
      1684: inst = 32'hc404206;
      1685: inst = 32'h8220000;
      1686: inst = 32'h10408000;
      1687: inst = 32'hc404207;
      1688: inst = 32'h8220000;
      1689: inst = 32'h10408000;
      1690: inst = 32'hc404208;
      1691: inst = 32'h8220000;
      1692: inst = 32'h10408000;
      1693: inst = 32'hc404209;
      1694: inst = 32'h8220000;
      1695: inst = 32'h10408000;
      1696: inst = 32'hc40420a;
      1697: inst = 32'h8220000;
      1698: inst = 32'h10408000;
      1699: inst = 32'hc40420b;
      1700: inst = 32'h8220000;
      1701: inst = 32'h10408000;
      1702: inst = 32'hc40420c;
      1703: inst = 32'h8220000;
      1704: inst = 32'h10408000;
      1705: inst = 32'hc40420d;
      1706: inst = 32'h8220000;
      1707: inst = 32'h10408000;
      1708: inst = 32'hc40420e;
      1709: inst = 32'h8220000;
      1710: inst = 32'h10408000;
      1711: inst = 32'hc40420f;
      1712: inst = 32'h8220000;
      1713: inst = 32'h10408000;
      1714: inst = 32'hc404210;
      1715: inst = 32'h8220000;
      1716: inst = 32'h10408000;
      1717: inst = 32'hc404211;
      1718: inst = 32'h8220000;
      1719: inst = 32'h10408000;
      1720: inst = 32'hc404212;
      1721: inst = 32'h8220000;
      1722: inst = 32'h10408000;
      1723: inst = 32'hc404213;
      1724: inst = 32'h8220000;
      1725: inst = 32'h10408000;
      1726: inst = 32'hc404214;
      1727: inst = 32'h8220000;
      1728: inst = 32'h10408000;
      1729: inst = 32'hc404215;
      1730: inst = 32'h8220000;
      1731: inst = 32'h10408000;
      1732: inst = 32'hc404216;
      1733: inst = 32'h8220000;
      1734: inst = 32'h10408000;
      1735: inst = 32'hc404217;
      1736: inst = 32'h8220000;
      1737: inst = 32'h10408000;
      1738: inst = 32'hc404218;
      1739: inst = 32'h8220000;
      1740: inst = 32'h10408000;
      1741: inst = 32'hc404219;
      1742: inst = 32'h8220000;
      1743: inst = 32'h10408000;
      1744: inst = 32'hc40421a;
      1745: inst = 32'h8220000;
      1746: inst = 32'h10408000;
      1747: inst = 32'hc40421b;
      1748: inst = 32'h8220000;
      1749: inst = 32'h10408000;
      1750: inst = 32'hc40421c;
      1751: inst = 32'h8220000;
      1752: inst = 32'h10408000;
      1753: inst = 32'hc40421d;
      1754: inst = 32'h8220000;
      1755: inst = 32'h10408000;
      1756: inst = 32'hc40421e;
      1757: inst = 32'h8220000;
      1758: inst = 32'h10408000;
      1759: inst = 32'hc40421f;
      1760: inst = 32'h8220000;
      1761: inst = 32'h10408000;
      1762: inst = 32'hc404220;
      1763: inst = 32'h8220000;
      1764: inst = 32'h10408000;
      1765: inst = 32'hc404221;
      1766: inst = 32'h8220000;
      1767: inst = 32'h10408000;
      1768: inst = 32'hc404222;
      1769: inst = 32'h8220000;
      1770: inst = 32'h10408000;
      1771: inst = 32'hc404223;
      1772: inst = 32'h8220000;
      1773: inst = 32'h10408000;
      1774: inst = 32'hc404224;
      1775: inst = 32'h8220000;
      1776: inst = 32'h10408000;
      1777: inst = 32'hc404225;
      1778: inst = 32'h8220000;
      1779: inst = 32'h10408000;
      1780: inst = 32'hc404226;
      1781: inst = 32'h8220000;
      1782: inst = 32'h10408000;
      1783: inst = 32'hc404227;
      1784: inst = 32'h8220000;
      1785: inst = 32'h10408000;
      1786: inst = 32'hc404228;
      1787: inst = 32'h8220000;
      1788: inst = 32'h10408000;
      1789: inst = 32'hc404229;
      1790: inst = 32'h8220000;
      1791: inst = 32'h10408000;
      1792: inst = 32'hc40422a;
      1793: inst = 32'h8220000;
      1794: inst = 32'h10408000;
      1795: inst = 32'hc40422c;
      1796: inst = 32'h8220000;
      1797: inst = 32'h10408000;
      1798: inst = 32'hc40422d;
      1799: inst = 32'h8220000;
      1800: inst = 32'h10408000;
      1801: inst = 32'hc40422e;
      1802: inst = 32'h8220000;
      1803: inst = 32'h10408000;
      1804: inst = 32'hc40422f;
      1805: inst = 32'h8220000;
      1806: inst = 32'h10408000;
      1807: inst = 32'hc404230;
      1808: inst = 32'h8220000;
      1809: inst = 32'h10408000;
      1810: inst = 32'hc404231;
      1811: inst = 32'h8220000;
      1812: inst = 32'h10408000;
      1813: inst = 32'hc404232;
      1814: inst = 32'h8220000;
      1815: inst = 32'h10408000;
      1816: inst = 32'hc404233;
      1817: inst = 32'h8220000;
      1818: inst = 32'h10408000;
      1819: inst = 32'hc404234;
      1820: inst = 32'h8220000;
      1821: inst = 32'h10408000;
      1822: inst = 32'hc404235;
      1823: inst = 32'h8220000;
      1824: inst = 32'h10408000;
      1825: inst = 32'hc404236;
      1826: inst = 32'h8220000;
      1827: inst = 32'h10408000;
      1828: inst = 32'hc404237;
      1829: inst = 32'h8220000;
      1830: inst = 32'h10408000;
      1831: inst = 32'hc404238;
      1832: inst = 32'h8220000;
      1833: inst = 32'h10408000;
      1834: inst = 32'hc404239;
      1835: inst = 32'h8220000;
      1836: inst = 32'h10408000;
      1837: inst = 32'hc40423a;
      1838: inst = 32'h8220000;
      1839: inst = 32'h10408000;
      1840: inst = 32'hc40423b;
      1841: inst = 32'h8220000;
      1842: inst = 32'h10408000;
      1843: inst = 32'hc404264;
      1844: inst = 32'h8220000;
      1845: inst = 32'h10408000;
      1846: inst = 32'hc404265;
      1847: inst = 32'h8220000;
      1848: inst = 32'h10408000;
      1849: inst = 32'hc404266;
      1850: inst = 32'h8220000;
      1851: inst = 32'h10408000;
      1852: inst = 32'hc404267;
      1853: inst = 32'h8220000;
      1854: inst = 32'h10408000;
      1855: inst = 32'hc404268;
      1856: inst = 32'h8220000;
      1857: inst = 32'h10408000;
      1858: inst = 32'hc404269;
      1859: inst = 32'h8220000;
      1860: inst = 32'h10408000;
      1861: inst = 32'hc40426a;
      1862: inst = 32'h8220000;
      1863: inst = 32'h10408000;
      1864: inst = 32'hc40426b;
      1865: inst = 32'h8220000;
      1866: inst = 32'h10408000;
      1867: inst = 32'hc40426c;
      1868: inst = 32'h8220000;
      1869: inst = 32'h10408000;
      1870: inst = 32'hc40426d;
      1871: inst = 32'h8220000;
      1872: inst = 32'h10408000;
      1873: inst = 32'hc40426e;
      1874: inst = 32'h8220000;
      1875: inst = 32'h10408000;
      1876: inst = 32'hc40426f;
      1877: inst = 32'h8220000;
      1878: inst = 32'h10408000;
      1879: inst = 32'hc404270;
      1880: inst = 32'h8220000;
      1881: inst = 32'h10408000;
      1882: inst = 32'hc404271;
      1883: inst = 32'h8220000;
      1884: inst = 32'h10408000;
      1885: inst = 32'hc404272;
      1886: inst = 32'h8220000;
      1887: inst = 32'h10408000;
      1888: inst = 32'hc404273;
      1889: inst = 32'h8220000;
      1890: inst = 32'h10408000;
      1891: inst = 32'hc404274;
      1892: inst = 32'h8220000;
      1893: inst = 32'h10408000;
      1894: inst = 32'hc404275;
      1895: inst = 32'h8220000;
      1896: inst = 32'h10408000;
      1897: inst = 32'hc404276;
      1898: inst = 32'h8220000;
      1899: inst = 32'h10408000;
      1900: inst = 32'hc404277;
      1901: inst = 32'h8220000;
      1902: inst = 32'h10408000;
      1903: inst = 32'hc404278;
      1904: inst = 32'h8220000;
      1905: inst = 32'h10408000;
      1906: inst = 32'hc404279;
      1907: inst = 32'h8220000;
      1908: inst = 32'h10408000;
      1909: inst = 32'hc40427a;
      1910: inst = 32'h8220000;
      1911: inst = 32'h10408000;
      1912: inst = 32'hc40427b;
      1913: inst = 32'h8220000;
      1914: inst = 32'h10408000;
      1915: inst = 32'hc40427c;
      1916: inst = 32'h8220000;
      1917: inst = 32'h10408000;
      1918: inst = 32'hc40427d;
      1919: inst = 32'h8220000;
      1920: inst = 32'h10408000;
      1921: inst = 32'hc40427e;
      1922: inst = 32'h8220000;
      1923: inst = 32'h10408000;
      1924: inst = 32'hc40427f;
      1925: inst = 32'h8220000;
      1926: inst = 32'h10408000;
      1927: inst = 32'hc404280;
      1928: inst = 32'h8220000;
      1929: inst = 32'h10408000;
      1930: inst = 32'hc404281;
      1931: inst = 32'h8220000;
      1932: inst = 32'h10408000;
      1933: inst = 32'hc404282;
      1934: inst = 32'h8220000;
      1935: inst = 32'h10408000;
      1936: inst = 32'hc404283;
      1937: inst = 32'h8220000;
      1938: inst = 32'h10408000;
      1939: inst = 32'hc404284;
      1940: inst = 32'h8220000;
      1941: inst = 32'h10408000;
      1942: inst = 32'hc404285;
      1943: inst = 32'h8220000;
      1944: inst = 32'h10408000;
      1945: inst = 32'hc404286;
      1946: inst = 32'h8220000;
      1947: inst = 32'h10408000;
      1948: inst = 32'hc404287;
      1949: inst = 32'h8220000;
      1950: inst = 32'h10408000;
      1951: inst = 32'hc404288;
      1952: inst = 32'h8220000;
      1953: inst = 32'h10408000;
      1954: inst = 32'hc404289;
      1955: inst = 32'h8220000;
      1956: inst = 32'h10408000;
      1957: inst = 32'hc40428a;
      1958: inst = 32'h8220000;
      1959: inst = 32'h10408000;
      1960: inst = 32'hc40428c;
      1961: inst = 32'h8220000;
      1962: inst = 32'h10408000;
      1963: inst = 32'hc40428d;
      1964: inst = 32'h8220000;
      1965: inst = 32'h10408000;
      1966: inst = 32'hc40428e;
      1967: inst = 32'h8220000;
      1968: inst = 32'h10408000;
      1969: inst = 32'hc40428f;
      1970: inst = 32'h8220000;
      1971: inst = 32'h10408000;
      1972: inst = 32'hc404290;
      1973: inst = 32'h8220000;
      1974: inst = 32'h10408000;
      1975: inst = 32'hc404291;
      1976: inst = 32'h8220000;
      1977: inst = 32'h10408000;
      1978: inst = 32'hc404292;
      1979: inst = 32'h8220000;
      1980: inst = 32'h10408000;
      1981: inst = 32'hc404293;
      1982: inst = 32'h8220000;
      1983: inst = 32'h10408000;
      1984: inst = 32'hc404294;
      1985: inst = 32'h8220000;
      1986: inst = 32'h10408000;
      1987: inst = 32'hc404295;
      1988: inst = 32'h8220000;
      1989: inst = 32'h10408000;
      1990: inst = 32'hc404296;
      1991: inst = 32'h8220000;
      1992: inst = 32'h10408000;
      1993: inst = 32'hc404297;
      1994: inst = 32'h8220000;
      1995: inst = 32'h10408000;
      1996: inst = 32'hc404298;
      1997: inst = 32'h8220000;
      1998: inst = 32'h10408000;
      1999: inst = 32'hc404299;
      2000: inst = 32'h8220000;
      2001: inst = 32'h10408000;
      2002: inst = 32'hc40429a;
      2003: inst = 32'h8220000;
      2004: inst = 32'h10408000;
      2005: inst = 32'hc40429b;
      2006: inst = 32'h8220000;
      2007: inst = 32'h10408000;
      2008: inst = 32'hc4042c4;
      2009: inst = 32'h8220000;
      2010: inst = 32'h10408000;
      2011: inst = 32'hc4042c5;
      2012: inst = 32'h8220000;
      2013: inst = 32'h10408000;
      2014: inst = 32'hc4042c6;
      2015: inst = 32'h8220000;
      2016: inst = 32'h10408000;
      2017: inst = 32'hc4042c7;
      2018: inst = 32'h8220000;
      2019: inst = 32'h10408000;
      2020: inst = 32'hc4042c8;
      2021: inst = 32'h8220000;
      2022: inst = 32'h10408000;
      2023: inst = 32'hc4042c9;
      2024: inst = 32'h8220000;
      2025: inst = 32'h10408000;
      2026: inst = 32'hc4042ca;
      2027: inst = 32'h8220000;
      2028: inst = 32'h10408000;
      2029: inst = 32'hc4042cb;
      2030: inst = 32'h8220000;
      2031: inst = 32'h10408000;
      2032: inst = 32'hc4042cc;
      2033: inst = 32'h8220000;
      2034: inst = 32'h10408000;
      2035: inst = 32'hc4042cd;
      2036: inst = 32'h8220000;
      2037: inst = 32'h10408000;
      2038: inst = 32'hc4042ce;
      2039: inst = 32'h8220000;
      2040: inst = 32'h10408000;
      2041: inst = 32'hc4042cf;
      2042: inst = 32'h8220000;
      2043: inst = 32'h10408000;
      2044: inst = 32'hc4042d0;
      2045: inst = 32'h8220000;
      2046: inst = 32'h10408000;
      2047: inst = 32'hc4042d1;
      2048: inst = 32'h8220000;
      2049: inst = 32'h10408000;
      2050: inst = 32'hc4042d2;
      2051: inst = 32'h8220000;
      2052: inst = 32'h10408000;
      2053: inst = 32'hc4042d3;
      2054: inst = 32'h8220000;
      2055: inst = 32'h10408000;
      2056: inst = 32'hc4042d4;
      2057: inst = 32'h8220000;
      2058: inst = 32'h10408000;
      2059: inst = 32'hc4042d5;
      2060: inst = 32'h8220000;
      2061: inst = 32'h10408000;
      2062: inst = 32'hc4042d6;
      2063: inst = 32'h8220000;
      2064: inst = 32'h10408000;
      2065: inst = 32'hc4042d7;
      2066: inst = 32'h8220000;
      2067: inst = 32'h10408000;
      2068: inst = 32'hc4042d8;
      2069: inst = 32'h8220000;
      2070: inst = 32'h10408000;
      2071: inst = 32'hc4042d9;
      2072: inst = 32'h8220000;
      2073: inst = 32'h10408000;
      2074: inst = 32'hc4042da;
      2075: inst = 32'h8220000;
      2076: inst = 32'h10408000;
      2077: inst = 32'hc4042db;
      2078: inst = 32'h8220000;
      2079: inst = 32'h10408000;
      2080: inst = 32'hc4042dc;
      2081: inst = 32'h8220000;
      2082: inst = 32'h10408000;
      2083: inst = 32'hc4042dd;
      2084: inst = 32'h8220000;
      2085: inst = 32'h10408000;
      2086: inst = 32'hc4042de;
      2087: inst = 32'h8220000;
      2088: inst = 32'h10408000;
      2089: inst = 32'hc4042df;
      2090: inst = 32'h8220000;
      2091: inst = 32'h10408000;
      2092: inst = 32'hc4042e0;
      2093: inst = 32'h8220000;
      2094: inst = 32'h10408000;
      2095: inst = 32'hc4042e1;
      2096: inst = 32'h8220000;
      2097: inst = 32'h10408000;
      2098: inst = 32'hc4042e2;
      2099: inst = 32'h8220000;
      2100: inst = 32'h10408000;
      2101: inst = 32'hc4042e3;
      2102: inst = 32'h8220000;
      2103: inst = 32'h10408000;
      2104: inst = 32'hc4042e4;
      2105: inst = 32'h8220000;
      2106: inst = 32'h10408000;
      2107: inst = 32'hc4042e5;
      2108: inst = 32'h8220000;
      2109: inst = 32'h10408000;
      2110: inst = 32'hc4042e6;
      2111: inst = 32'h8220000;
      2112: inst = 32'h10408000;
      2113: inst = 32'hc4042e7;
      2114: inst = 32'h8220000;
      2115: inst = 32'h10408000;
      2116: inst = 32'hc4042e8;
      2117: inst = 32'h8220000;
      2118: inst = 32'h10408000;
      2119: inst = 32'hc4042e9;
      2120: inst = 32'h8220000;
      2121: inst = 32'h10408000;
      2122: inst = 32'hc4042ee;
      2123: inst = 32'h8220000;
      2124: inst = 32'h10408000;
      2125: inst = 32'hc4042ef;
      2126: inst = 32'h8220000;
      2127: inst = 32'h10408000;
      2128: inst = 32'hc4042f0;
      2129: inst = 32'h8220000;
      2130: inst = 32'h10408000;
      2131: inst = 32'hc4042f1;
      2132: inst = 32'h8220000;
      2133: inst = 32'h10408000;
      2134: inst = 32'hc4042f2;
      2135: inst = 32'h8220000;
      2136: inst = 32'h10408000;
      2137: inst = 32'hc4042f3;
      2138: inst = 32'h8220000;
      2139: inst = 32'h10408000;
      2140: inst = 32'hc4042f4;
      2141: inst = 32'h8220000;
      2142: inst = 32'h10408000;
      2143: inst = 32'hc4042f5;
      2144: inst = 32'h8220000;
      2145: inst = 32'h10408000;
      2146: inst = 32'hc4042f6;
      2147: inst = 32'h8220000;
      2148: inst = 32'h10408000;
      2149: inst = 32'hc4042f7;
      2150: inst = 32'h8220000;
      2151: inst = 32'h10408000;
      2152: inst = 32'hc4042f8;
      2153: inst = 32'h8220000;
      2154: inst = 32'h10408000;
      2155: inst = 32'hc4042f9;
      2156: inst = 32'h8220000;
      2157: inst = 32'h10408000;
      2158: inst = 32'hc4042fa;
      2159: inst = 32'h8220000;
      2160: inst = 32'h10408000;
      2161: inst = 32'hc4042fb;
      2162: inst = 32'h8220000;
      2163: inst = 32'h10408000;
      2164: inst = 32'hc404324;
      2165: inst = 32'h8220000;
      2166: inst = 32'h10408000;
      2167: inst = 32'hc404325;
      2168: inst = 32'h8220000;
      2169: inst = 32'h10408000;
      2170: inst = 32'hc404326;
      2171: inst = 32'h8220000;
      2172: inst = 32'h10408000;
      2173: inst = 32'hc404327;
      2174: inst = 32'h8220000;
      2175: inst = 32'h10408000;
      2176: inst = 32'hc404328;
      2177: inst = 32'h8220000;
      2178: inst = 32'h10408000;
      2179: inst = 32'hc404329;
      2180: inst = 32'h8220000;
      2181: inst = 32'h10408000;
      2182: inst = 32'hc40432a;
      2183: inst = 32'h8220000;
      2184: inst = 32'h10408000;
      2185: inst = 32'hc40432b;
      2186: inst = 32'h8220000;
      2187: inst = 32'h10408000;
      2188: inst = 32'hc40432c;
      2189: inst = 32'h8220000;
      2190: inst = 32'h10408000;
      2191: inst = 32'hc40432d;
      2192: inst = 32'h8220000;
      2193: inst = 32'h10408000;
      2194: inst = 32'hc40432e;
      2195: inst = 32'h8220000;
      2196: inst = 32'h10408000;
      2197: inst = 32'hc40432f;
      2198: inst = 32'h8220000;
      2199: inst = 32'h10408000;
      2200: inst = 32'hc404330;
      2201: inst = 32'h8220000;
      2202: inst = 32'h10408000;
      2203: inst = 32'hc404331;
      2204: inst = 32'h8220000;
      2205: inst = 32'h10408000;
      2206: inst = 32'hc404332;
      2207: inst = 32'h8220000;
      2208: inst = 32'h10408000;
      2209: inst = 32'hc404333;
      2210: inst = 32'h8220000;
      2211: inst = 32'h10408000;
      2212: inst = 32'hc404334;
      2213: inst = 32'h8220000;
      2214: inst = 32'h10408000;
      2215: inst = 32'hc404335;
      2216: inst = 32'h8220000;
      2217: inst = 32'h10408000;
      2218: inst = 32'hc404336;
      2219: inst = 32'h8220000;
      2220: inst = 32'h10408000;
      2221: inst = 32'hc404337;
      2222: inst = 32'h8220000;
      2223: inst = 32'h10408000;
      2224: inst = 32'hc404338;
      2225: inst = 32'h8220000;
      2226: inst = 32'h10408000;
      2227: inst = 32'hc404339;
      2228: inst = 32'h8220000;
      2229: inst = 32'h10408000;
      2230: inst = 32'hc40433a;
      2231: inst = 32'h8220000;
      2232: inst = 32'h10408000;
      2233: inst = 32'hc40433b;
      2234: inst = 32'h8220000;
      2235: inst = 32'h10408000;
      2236: inst = 32'hc40433c;
      2237: inst = 32'h8220000;
      2238: inst = 32'h10408000;
      2239: inst = 32'hc40433d;
      2240: inst = 32'h8220000;
      2241: inst = 32'h10408000;
      2242: inst = 32'hc40433e;
      2243: inst = 32'h8220000;
      2244: inst = 32'h10408000;
      2245: inst = 32'hc40433f;
      2246: inst = 32'h8220000;
      2247: inst = 32'h10408000;
      2248: inst = 32'hc404340;
      2249: inst = 32'h8220000;
      2250: inst = 32'h10408000;
      2251: inst = 32'hc404341;
      2252: inst = 32'h8220000;
      2253: inst = 32'h10408000;
      2254: inst = 32'hc404342;
      2255: inst = 32'h8220000;
      2256: inst = 32'h10408000;
      2257: inst = 32'hc404343;
      2258: inst = 32'h8220000;
      2259: inst = 32'h10408000;
      2260: inst = 32'hc404344;
      2261: inst = 32'h8220000;
      2262: inst = 32'h10408000;
      2263: inst = 32'hc404345;
      2264: inst = 32'h8220000;
      2265: inst = 32'h10408000;
      2266: inst = 32'hc404346;
      2267: inst = 32'h8220000;
      2268: inst = 32'h10408000;
      2269: inst = 32'hc404347;
      2270: inst = 32'h8220000;
      2271: inst = 32'h10408000;
      2272: inst = 32'hc404348;
      2273: inst = 32'h8220000;
      2274: inst = 32'h10408000;
      2275: inst = 32'hc40434f;
      2276: inst = 32'h8220000;
      2277: inst = 32'h10408000;
      2278: inst = 32'hc404350;
      2279: inst = 32'h8220000;
      2280: inst = 32'h10408000;
      2281: inst = 32'hc404351;
      2282: inst = 32'h8220000;
      2283: inst = 32'h10408000;
      2284: inst = 32'hc404352;
      2285: inst = 32'h8220000;
      2286: inst = 32'h10408000;
      2287: inst = 32'hc404353;
      2288: inst = 32'h8220000;
      2289: inst = 32'h10408000;
      2290: inst = 32'hc404354;
      2291: inst = 32'h8220000;
      2292: inst = 32'h10408000;
      2293: inst = 32'hc404355;
      2294: inst = 32'h8220000;
      2295: inst = 32'h10408000;
      2296: inst = 32'hc404356;
      2297: inst = 32'h8220000;
      2298: inst = 32'h10408000;
      2299: inst = 32'hc404357;
      2300: inst = 32'h8220000;
      2301: inst = 32'h10408000;
      2302: inst = 32'hc404358;
      2303: inst = 32'h8220000;
      2304: inst = 32'h10408000;
      2305: inst = 32'hc404359;
      2306: inst = 32'h8220000;
      2307: inst = 32'h10408000;
      2308: inst = 32'hc40435a;
      2309: inst = 32'h8220000;
      2310: inst = 32'h10408000;
      2311: inst = 32'hc40435b;
      2312: inst = 32'h8220000;
      2313: inst = 32'h10408000;
      2314: inst = 32'hc404384;
      2315: inst = 32'h8220000;
      2316: inst = 32'h10408000;
      2317: inst = 32'hc404385;
      2318: inst = 32'h8220000;
      2319: inst = 32'h10408000;
      2320: inst = 32'hc404386;
      2321: inst = 32'h8220000;
      2322: inst = 32'h10408000;
      2323: inst = 32'hc404387;
      2324: inst = 32'h8220000;
      2325: inst = 32'h10408000;
      2326: inst = 32'hc404388;
      2327: inst = 32'h8220000;
      2328: inst = 32'h10408000;
      2329: inst = 32'hc404389;
      2330: inst = 32'h8220000;
      2331: inst = 32'h10408000;
      2332: inst = 32'hc40438a;
      2333: inst = 32'h8220000;
      2334: inst = 32'h10408000;
      2335: inst = 32'hc40438b;
      2336: inst = 32'h8220000;
      2337: inst = 32'h10408000;
      2338: inst = 32'hc40438c;
      2339: inst = 32'h8220000;
      2340: inst = 32'h10408000;
      2341: inst = 32'hc40438d;
      2342: inst = 32'h8220000;
      2343: inst = 32'h10408000;
      2344: inst = 32'hc40438e;
      2345: inst = 32'h8220000;
      2346: inst = 32'h10408000;
      2347: inst = 32'hc40438f;
      2348: inst = 32'h8220000;
      2349: inst = 32'h10408000;
      2350: inst = 32'hc404390;
      2351: inst = 32'h8220000;
      2352: inst = 32'h10408000;
      2353: inst = 32'hc404391;
      2354: inst = 32'h8220000;
      2355: inst = 32'h10408000;
      2356: inst = 32'hc404392;
      2357: inst = 32'h8220000;
      2358: inst = 32'h10408000;
      2359: inst = 32'hc404393;
      2360: inst = 32'h8220000;
      2361: inst = 32'h10408000;
      2362: inst = 32'hc404394;
      2363: inst = 32'h8220000;
      2364: inst = 32'h10408000;
      2365: inst = 32'hc404395;
      2366: inst = 32'h8220000;
      2367: inst = 32'h10408000;
      2368: inst = 32'hc404396;
      2369: inst = 32'h8220000;
      2370: inst = 32'h10408000;
      2371: inst = 32'hc404397;
      2372: inst = 32'h8220000;
      2373: inst = 32'h10408000;
      2374: inst = 32'hc404398;
      2375: inst = 32'h8220000;
      2376: inst = 32'h10408000;
      2377: inst = 32'hc404399;
      2378: inst = 32'h8220000;
      2379: inst = 32'h10408000;
      2380: inst = 32'hc40439a;
      2381: inst = 32'h8220000;
      2382: inst = 32'h10408000;
      2383: inst = 32'hc40439b;
      2384: inst = 32'h8220000;
      2385: inst = 32'h10408000;
      2386: inst = 32'hc40439c;
      2387: inst = 32'h8220000;
      2388: inst = 32'h10408000;
      2389: inst = 32'hc40439d;
      2390: inst = 32'h8220000;
      2391: inst = 32'h10408000;
      2392: inst = 32'hc40439e;
      2393: inst = 32'h8220000;
      2394: inst = 32'h10408000;
      2395: inst = 32'hc40439f;
      2396: inst = 32'h8220000;
      2397: inst = 32'h10408000;
      2398: inst = 32'hc4043a0;
      2399: inst = 32'h8220000;
      2400: inst = 32'h10408000;
      2401: inst = 32'hc4043a1;
      2402: inst = 32'h8220000;
      2403: inst = 32'h10408000;
      2404: inst = 32'hc4043a2;
      2405: inst = 32'h8220000;
      2406: inst = 32'h10408000;
      2407: inst = 32'hc4043a3;
      2408: inst = 32'h8220000;
      2409: inst = 32'h10408000;
      2410: inst = 32'hc4043a4;
      2411: inst = 32'h8220000;
      2412: inst = 32'h10408000;
      2413: inst = 32'hc4043a5;
      2414: inst = 32'h8220000;
      2415: inst = 32'h10408000;
      2416: inst = 32'hc4043a6;
      2417: inst = 32'h8220000;
      2418: inst = 32'h10408000;
      2419: inst = 32'hc4043b1;
      2420: inst = 32'h8220000;
      2421: inst = 32'h10408000;
      2422: inst = 32'hc4043b2;
      2423: inst = 32'h8220000;
      2424: inst = 32'h10408000;
      2425: inst = 32'hc4043b3;
      2426: inst = 32'h8220000;
      2427: inst = 32'h10408000;
      2428: inst = 32'hc4043b4;
      2429: inst = 32'h8220000;
      2430: inst = 32'h10408000;
      2431: inst = 32'hc4043b5;
      2432: inst = 32'h8220000;
      2433: inst = 32'h10408000;
      2434: inst = 32'hc4043b6;
      2435: inst = 32'h8220000;
      2436: inst = 32'h10408000;
      2437: inst = 32'hc4043b7;
      2438: inst = 32'h8220000;
      2439: inst = 32'h10408000;
      2440: inst = 32'hc4043b8;
      2441: inst = 32'h8220000;
      2442: inst = 32'h10408000;
      2443: inst = 32'hc4043b9;
      2444: inst = 32'h8220000;
      2445: inst = 32'h10408000;
      2446: inst = 32'hc4043ba;
      2447: inst = 32'h8220000;
      2448: inst = 32'h10408000;
      2449: inst = 32'hc4043bb;
      2450: inst = 32'h8220000;
      2451: inst = 32'h10408000;
      2452: inst = 32'hc4043e4;
      2453: inst = 32'h8220000;
      2454: inst = 32'h10408000;
      2455: inst = 32'hc4043e5;
      2456: inst = 32'h8220000;
      2457: inst = 32'h10408000;
      2458: inst = 32'hc4043e6;
      2459: inst = 32'h8220000;
      2460: inst = 32'h10408000;
      2461: inst = 32'hc4043e7;
      2462: inst = 32'h8220000;
      2463: inst = 32'h10408000;
      2464: inst = 32'hc4043e8;
      2465: inst = 32'h8220000;
      2466: inst = 32'h10408000;
      2467: inst = 32'hc4043e9;
      2468: inst = 32'h8220000;
      2469: inst = 32'h10408000;
      2470: inst = 32'hc4043ea;
      2471: inst = 32'h8220000;
      2472: inst = 32'h10408000;
      2473: inst = 32'hc4043eb;
      2474: inst = 32'h8220000;
      2475: inst = 32'h10408000;
      2476: inst = 32'hc4043ec;
      2477: inst = 32'h8220000;
      2478: inst = 32'h10408000;
      2479: inst = 32'hc4043ed;
      2480: inst = 32'h8220000;
      2481: inst = 32'h10408000;
      2482: inst = 32'hc4043ee;
      2483: inst = 32'h8220000;
      2484: inst = 32'h10408000;
      2485: inst = 32'hc4043ef;
      2486: inst = 32'h8220000;
      2487: inst = 32'h10408000;
      2488: inst = 32'hc4043f0;
      2489: inst = 32'h8220000;
      2490: inst = 32'h10408000;
      2491: inst = 32'hc4043f1;
      2492: inst = 32'h8220000;
      2493: inst = 32'h10408000;
      2494: inst = 32'hc4043f2;
      2495: inst = 32'h8220000;
      2496: inst = 32'h10408000;
      2497: inst = 32'hc4043f3;
      2498: inst = 32'h8220000;
      2499: inst = 32'h10408000;
      2500: inst = 32'hc4043f4;
      2501: inst = 32'h8220000;
      2502: inst = 32'h10408000;
      2503: inst = 32'hc4043f5;
      2504: inst = 32'h8220000;
      2505: inst = 32'h10408000;
      2506: inst = 32'hc4043f6;
      2507: inst = 32'h8220000;
      2508: inst = 32'h10408000;
      2509: inst = 32'hc4043f7;
      2510: inst = 32'h8220000;
      2511: inst = 32'h10408000;
      2512: inst = 32'hc4043f8;
      2513: inst = 32'h8220000;
      2514: inst = 32'h10408000;
      2515: inst = 32'hc4043f9;
      2516: inst = 32'h8220000;
      2517: inst = 32'h10408000;
      2518: inst = 32'hc4043fa;
      2519: inst = 32'h8220000;
      2520: inst = 32'h10408000;
      2521: inst = 32'hc4043fb;
      2522: inst = 32'h8220000;
      2523: inst = 32'h10408000;
      2524: inst = 32'hc4043fc;
      2525: inst = 32'h8220000;
      2526: inst = 32'h10408000;
      2527: inst = 32'hc4043fd;
      2528: inst = 32'h8220000;
      2529: inst = 32'h10408000;
      2530: inst = 32'hc4043fe;
      2531: inst = 32'h8220000;
      2532: inst = 32'h10408000;
      2533: inst = 32'hc4043ff;
      2534: inst = 32'h8220000;
      2535: inst = 32'h10408000;
      2536: inst = 32'hc404400;
      2537: inst = 32'h8220000;
      2538: inst = 32'h10408000;
      2539: inst = 32'hc404401;
      2540: inst = 32'h8220000;
      2541: inst = 32'h10408000;
      2542: inst = 32'hc404402;
      2543: inst = 32'h8220000;
      2544: inst = 32'h10408000;
      2545: inst = 32'hc404403;
      2546: inst = 32'h8220000;
      2547: inst = 32'h10408000;
      2548: inst = 32'hc404404;
      2549: inst = 32'h8220000;
      2550: inst = 32'h10408000;
      2551: inst = 32'hc404405;
      2552: inst = 32'h8220000;
      2553: inst = 32'h10408000;
      2554: inst = 32'hc404412;
      2555: inst = 32'h8220000;
      2556: inst = 32'h10408000;
      2557: inst = 32'hc404413;
      2558: inst = 32'h8220000;
      2559: inst = 32'h10408000;
      2560: inst = 32'hc404414;
      2561: inst = 32'h8220000;
      2562: inst = 32'h10408000;
      2563: inst = 32'hc404415;
      2564: inst = 32'h8220000;
      2565: inst = 32'h10408000;
      2566: inst = 32'hc404416;
      2567: inst = 32'h8220000;
      2568: inst = 32'h10408000;
      2569: inst = 32'hc404417;
      2570: inst = 32'h8220000;
      2571: inst = 32'h10408000;
      2572: inst = 32'hc404418;
      2573: inst = 32'h8220000;
      2574: inst = 32'h10408000;
      2575: inst = 32'hc404419;
      2576: inst = 32'h8220000;
      2577: inst = 32'h10408000;
      2578: inst = 32'hc40441a;
      2579: inst = 32'h8220000;
      2580: inst = 32'h10408000;
      2581: inst = 32'hc40441b;
      2582: inst = 32'h8220000;
      2583: inst = 32'h10408000;
      2584: inst = 32'hc404444;
      2585: inst = 32'h8220000;
      2586: inst = 32'h10408000;
      2587: inst = 32'hc404445;
      2588: inst = 32'h8220000;
      2589: inst = 32'h10408000;
      2590: inst = 32'hc404446;
      2591: inst = 32'h8220000;
      2592: inst = 32'h10408000;
      2593: inst = 32'hc404447;
      2594: inst = 32'h8220000;
      2595: inst = 32'h10408000;
      2596: inst = 32'hc404448;
      2597: inst = 32'h8220000;
      2598: inst = 32'h10408000;
      2599: inst = 32'hc404449;
      2600: inst = 32'h8220000;
      2601: inst = 32'h10408000;
      2602: inst = 32'hc40444a;
      2603: inst = 32'h8220000;
      2604: inst = 32'h10408000;
      2605: inst = 32'hc40444b;
      2606: inst = 32'h8220000;
      2607: inst = 32'h10408000;
      2608: inst = 32'hc40444c;
      2609: inst = 32'h8220000;
      2610: inst = 32'h10408000;
      2611: inst = 32'hc40444d;
      2612: inst = 32'h8220000;
      2613: inst = 32'h10408000;
      2614: inst = 32'hc40444e;
      2615: inst = 32'h8220000;
      2616: inst = 32'h10408000;
      2617: inst = 32'hc40444f;
      2618: inst = 32'h8220000;
      2619: inst = 32'h10408000;
      2620: inst = 32'hc404450;
      2621: inst = 32'h8220000;
      2622: inst = 32'h10408000;
      2623: inst = 32'hc404451;
      2624: inst = 32'h8220000;
      2625: inst = 32'h10408000;
      2626: inst = 32'hc404452;
      2627: inst = 32'h8220000;
      2628: inst = 32'h10408000;
      2629: inst = 32'hc404453;
      2630: inst = 32'h8220000;
      2631: inst = 32'h10408000;
      2632: inst = 32'hc404454;
      2633: inst = 32'h8220000;
      2634: inst = 32'h10408000;
      2635: inst = 32'hc404455;
      2636: inst = 32'h8220000;
      2637: inst = 32'h10408000;
      2638: inst = 32'hc404456;
      2639: inst = 32'h8220000;
      2640: inst = 32'h10408000;
      2641: inst = 32'hc404457;
      2642: inst = 32'h8220000;
      2643: inst = 32'h10408000;
      2644: inst = 32'hc404458;
      2645: inst = 32'h8220000;
      2646: inst = 32'h10408000;
      2647: inst = 32'hc404459;
      2648: inst = 32'h8220000;
      2649: inst = 32'h10408000;
      2650: inst = 32'hc40445a;
      2651: inst = 32'h8220000;
      2652: inst = 32'h10408000;
      2653: inst = 32'hc40445b;
      2654: inst = 32'h8220000;
      2655: inst = 32'h10408000;
      2656: inst = 32'hc40445c;
      2657: inst = 32'h8220000;
      2658: inst = 32'h10408000;
      2659: inst = 32'hc40445d;
      2660: inst = 32'h8220000;
      2661: inst = 32'h10408000;
      2662: inst = 32'hc40445e;
      2663: inst = 32'h8220000;
      2664: inst = 32'h10408000;
      2665: inst = 32'hc40445f;
      2666: inst = 32'h8220000;
      2667: inst = 32'h10408000;
      2668: inst = 32'hc404460;
      2669: inst = 32'h8220000;
      2670: inst = 32'h10408000;
      2671: inst = 32'hc404461;
      2672: inst = 32'h8220000;
      2673: inst = 32'h10408000;
      2674: inst = 32'hc404462;
      2675: inst = 32'h8220000;
      2676: inst = 32'h10408000;
      2677: inst = 32'hc404463;
      2678: inst = 32'h8220000;
      2679: inst = 32'h10408000;
      2680: inst = 32'hc404464;
      2681: inst = 32'h8220000;
      2682: inst = 32'h10408000;
      2683: inst = 32'hc404465;
      2684: inst = 32'h8220000;
      2685: inst = 32'h10408000;
      2686: inst = 32'hc404466;
      2687: inst = 32'h8220000;
      2688: inst = 32'h10408000;
      2689: inst = 32'hc404467;
      2690: inst = 32'h8220000;
      2691: inst = 32'h10408000;
      2692: inst = 32'hc404468;
      2693: inst = 32'h8220000;
      2694: inst = 32'h10408000;
      2695: inst = 32'hc404469;
      2696: inst = 32'h8220000;
      2697: inst = 32'h10408000;
      2698: inst = 32'hc40446e;
      2699: inst = 32'h8220000;
      2700: inst = 32'h10408000;
      2701: inst = 32'hc40446f;
      2702: inst = 32'h8220000;
      2703: inst = 32'h10408000;
      2704: inst = 32'hc404470;
      2705: inst = 32'h8220000;
      2706: inst = 32'h10408000;
      2707: inst = 32'hc404471;
      2708: inst = 32'h8220000;
      2709: inst = 32'h10408000;
      2710: inst = 32'hc404472;
      2711: inst = 32'h8220000;
      2712: inst = 32'h10408000;
      2713: inst = 32'hc404473;
      2714: inst = 32'h8220000;
      2715: inst = 32'h10408000;
      2716: inst = 32'hc404474;
      2717: inst = 32'h8220000;
      2718: inst = 32'h10408000;
      2719: inst = 32'hc404475;
      2720: inst = 32'h8220000;
      2721: inst = 32'h10408000;
      2722: inst = 32'hc404476;
      2723: inst = 32'h8220000;
      2724: inst = 32'h10408000;
      2725: inst = 32'hc404477;
      2726: inst = 32'h8220000;
      2727: inst = 32'h10408000;
      2728: inst = 32'hc404478;
      2729: inst = 32'h8220000;
      2730: inst = 32'h10408000;
      2731: inst = 32'hc404479;
      2732: inst = 32'h8220000;
      2733: inst = 32'h10408000;
      2734: inst = 32'hc40447a;
      2735: inst = 32'h8220000;
      2736: inst = 32'h10408000;
      2737: inst = 32'hc40447b;
      2738: inst = 32'h8220000;
      2739: inst = 32'h10408000;
      2740: inst = 32'hc4044a4;
      2741: inst = 32'h8220000;
      2742: inst = 32'h10408000;
      2743: inst = 32'hc4044a5;
      2744: inst = 32'h8220000;
      2745: inst = 32'h10408000;
      2746: inst = 32'hc4044a6;
      2747: inst = 32'h8220000;
      2748: inst = 32'h10408000;
      2749: inst = 32'hc4044a7;
      2750: inst = 32'h8220000;
      2751: inst = 32'h10408000;
      2752: inst = 32'hc4044a8;
      2753: inst = 32'h8220000;
      2754: inst = 32'h10408000;
      2755: inst = 32'hc4044a9;
      2756: inst = 32'h8220000;
      2757: inst = 32'h10408000;
      2758: inst = 32'hc4044aa;
      2759: inst = 32'h8220000;
      2760: inst = 32'h10408000;
      2761: inst = 32'hc4044ab;
      2762: inst = 32'h8220000;
      2763: inst = 32'h10408000;
      2764: inst = 32'hc4044ac;
      2765: inst = 32'h8220000;
      2766: inst = 32'h10408000;
      2767: inst = 32'hc4044ad;
      2768: inst = 32'h8220000;
      2769: inst = 32'h10408000;
      2770: inst = 32'hc4044ae;
      2771: inst = 32'h8220000;
      2772: inst = 32'h10408000;
      2773: inst = 32'hc4044af;
      2774: inst = 32'h8220000;
      2775: inst = 32'h10408000;
      2776: inst = 32'hc4044b0;
      2777: inst = 32'h8220000;
      2778: inst = 32'h10408000;
      2779: inst = 32'hc4044b1;
      2780: inst = 32'h8220000;
      2781: inst = 32'h10408000;
      2782: inst = 32'hc4044b6;
      2783: inst = 32'h8220000;
      2784: inst = 32'h10408000;
      2785: inst = 32'hc4044b7;
      2786: inst = 32'h8220000;
      2787: inst = 32'h10408000;
      2788: inst = 32'hc4044b8;
      2789: inst = 32'h8220000;
      2790: inst = 32'h10408000;
      2791: inst = 32'hc4044b9;
      2792: inst = 32'h8220000;
      2793: inst = 32'h10408000;
      2794: inst = 32'hc4044ba;
      2795: inst = 32'h8220000;
      2796: inst = 32'h10408000;
      2797: inst = 32'hc4044bb;
      2798: inst = 32'h8220000;
      2799: inst = 32'h10408000;
      2800: inst = 32'hc4044bc;
      2801: inst = 32'h8220000;
      2802: inst = 32'h10408000;
      2803: inst = 32'hc4044bd;
      2804: inst = 32'h8220000;
      2805: inst = 32'h10408000;
      2806: inst = 32'hc4044be;
      2807: inst = 32'h8220000;
      2808: inst = 32'h10408000;
      2809: inst = 32'hc4044bf;
      2810: inst = 32'h8220000;
      2811: inst = 32'h10408000;
      2812: inst = 32'hc4044c0;
      2813: inst = 32'h8220000;
      2814: inst = 32'h10408000;
      2815: inst = 32'hc4044c1;
      2816: inst = 32'h8220000;
      2817: inst = 32'h10408000;
      2818: inst = 32'hc4044c2;
      2819: inst = 32'h8220000;
      2820: inst = 32'h10408000;
      2821: inst = 32'hc4044c3;
      2822: inst = 32'h8220000;
      2823: inst = 32'h10408000;
      2824: inst = 32'hc4044c4;
      2825: inst = 32'h8220000;
      2826: inst = 32'h10408000;
      2827: inst = 32'hc4044c5;
      2828: inst = 32'h8220000;
      2829: inst = 32'h10408000;
      2830: inst = 32'hc4044c6;
      2831: inst = 32'h8220000;
      2832: inst = 32'h10408000;
      2833: inst = 32'hc4044c7;
      2834: inst = 32'h8220000;
      2835: inst = 32'h10408000;
      2836: inst = 32'hc4044c8;
      2837: inst = 32'h8220000;
      2838: inst = 32'h10408000;
      2839: inst = 32'hc4044c9;
      2840: inst = 32'h8220000;
      2841: inst = 32'h10408000;
      2842: inst = 32'hc4044ca;
      2843: inst = 32'h8220000;
      2844: inst = 32'h10408000;
      2845: inst = 32'hc4044cd;
      2846: inst = 32'h8220000;
      2847: inst = 32'h10408000;
      2848: inst = 32'hc4044ce;
      2849: inst = 32'h8220000;
      2850: inst = 32'h10408000;
      2851: inst = 32'hc4044cf;
      2852: inst = 32'h8220000;
      2853: inst = 32'h10408000;
      2854: inst = 32'hc4044d0;
      2855: inst = 32'h8220000;
      2856: inst = 32'h10408000;
      2857: inst = 32'hc4044d1;
      2858: inst = 32'h8220000;
      2859: inst = 32'h10408000;
      2860: inst = 32'hc4044d2;
      2861: inst = 32'h8220000;
      2862: inst = 32'h10408000;
      2863: inst = 32'hc4044d3;
      2864: inst = 32'h8220000;
      2865: inst = 32'h10408000;
      2866: inst = 32'hc4044d4;
      2867: inst = 32'h8220000;
      2868: inst = 32'h10408000;
      2869: inst = 32'hc4044d5;
      2870: inst = 32'h8220000;
      2871: inst = 32'h10408000;
      2872: inst = 32'hc4044d6;
      2873: inst = 32'h8220000;
      2874: inst = 32'h10408000;
      2875: inst = 32'hc4044d7;
      2876: inst = 32'h8220000;
      2877: inst = 32'h10408000;
      2878: inst = 32'hc4044d8;
      2879: inst = 32'h8220000;
      2880: inst = 32'h10408000;
      2881: inst = 32'hc4044d9;
      2882: inst = 32'h8220000;
      2883: inst = 32'h10408000;
      2884: inst = 32'hc4044da;
      2885: inst = 32'h8220000;
      2886: inst = 32'h10408000;
      2887: inst = 32'hc4044db;
      2888: inst = 32'h8220000;
      2889: inst = 32'h10408000;
      2890: inst = 32'hc404504;
      2891: inst = 32'h8220000;
      2892: inst = 32'h10408000;
      2893: inst = 32'hc404505;
      2894: inst = 32'h8220000;
      2895: inst = 32'h10408000;
      2896: inst = 32'hc404506;
      2897: inst = 32'h8220000;
      2898: inst = 32'h10408000;
      2899: inst = 32'hc404507;
      2900: inst = 32'h8220000;
      2901: inst = 32'h10408000;
      2902: inst = 32'hc404508;
      2903: inst = 32'h8220000;
      2904: inst = 32'h10408000;
      2905: inst = 32'hc404509;
      2906: inst = 32'h8220000;
      2907: inst = 32'h10408000;
      2908: inst = 32'hc40450a;
      2909: inst = 32'h8220000;
      2910: inst = 32'h10408000;
      2911: inst = 32'hc40450b;
      2912: inst = 32'h8220000;
      2913: inst = 32'h10408000;
      2914: inst = 32'hc40450c;
      2915: inst = 32'h8220000;
      2916: inst = 32'h10408000;
      2917: inst = 32'hc40450d;
      2918: inst = 32'h8220000;
      2919: inst = 32'h10408000;
      2920: inst = 32'hc40450e;
      2921: inst = 32'h8220000;
      2922: inst = 32'h10408000;
      2923: inst = 32'hc40450f;
      2924: inst = 32'h8220000;
      2925: inst = 32'h10408000;
      2926: inst = 32'hc404510;
      2927: inst = 32'h8220000;
      2928: inst = 32'h10408000;
      2929: inst = 32'hc404511;
      2930: inst = 32'h8220000;
      2931: inst = 32'h10408000;
      2932: inst = 32'hc404512;
      2933: inst = 32'h8220000;
      2934: inst = 32'h10408000;
      2935: inst = 32'hc404515;
      2936: inst = 32'h8220000;
      2937: inst = 32'h10408000;
      2938: inst = 32'hc404516;
      2939: inst = 32'h8220000;
      2940: inst = 32'h10408000;
      2941: inst = 32'hc404517;
      2942: inst = 32'h8220000;
      2943: inst = 32'h10408000;
      2944: inst = 32'hc404518;
      2945: inst = 32'h8220000;
      2946: inst = 32'h10408000;
      2947: inst = 32'hc404519;
      2948: inst = 32'h8220000;
      2949: inst = 32'h10408000;
      2950: inst = 32'hc40451a;
      2951: inst = 32'h8220000;
      2952: inst = 32'h10408000;
      2953: inst = 32'hc40451b;
      2954: inst = 32'h8220000;
      2955: inst = 32'h10408000;
      2956: inst = 32'hc40451c;
      2957: inst = 32'h8220000;
      2958: inst = 32'h10408000;
      2959: inst = 32'hc40451d;
      2960: inst = 32'h8220000;
      2961: inst = 32'h10408000;
      2962: inst = 32'hc40451e;
      2963: inst = 32'h8220000;
      2964: inst = 32'h10408000;
      2965: inst = 32'hc40451f;
      2966: inst = 32'h8220000;
      2967: inst = 32'h10408000;
      2968: inst = 32'hc404520;
      2969: inst = 32'h8220000;
      2970: inst = 32'h10408000;
      2971: inst = 32'hc404521;
      2972: inst = 32'h8220000;
      2973: inst = 32'h10408000;
      2974: inst = 32'hc404522;
      2975: inst = 32'h8220000;
      2976: inst = 32'h10408000;
      2977: inst = 32'hc404523;
      2978: inst = 32'h8220000;
      2979: inst = 32'h10408000;
      2980: inst = 32'hc404524;
      2981: inst = 32'h8220000;
      2982: inst = 32'h10408000;
      2983: inst = 32'hc404525;
      2984: inst = 32'h8220000;
      2985: inst = 32'h10408000;
      2986: inst = 32'hc404526;
      2987: inst = 32'h8220000;
      2988: inst = 32'h10408000;
      2989: inst = 32'hc404527;
      2990: inst = 32'h8220000;
      2991: inst = 32'h10408000;
      2992: inst = 32'hc404528;
      2993: inst = 32'h8220000;
      2994: inst = 32'h10408000;
      2995: inst = 32'hc404529;
      2996: inst = 32'h8220000;
      2997: inst = 32'h10408000;
      2998: inst = 32'hc40452a;
      2999: inst = 32'h8220000;
      3000: inst = 32'h10408000;
      3001: inst = 32'hc40452b;
      3002: inst = 32'h8220000;
      3003: inst = 32'h10408000;
      3004: inst = 32'hc40452c;
      3005: inst = 32'h8220000;
      3006: inst = 32'h10408000;
      3007: inst = 32'hc40452d;
      3008: inst = 32'h8220000;
      3009: inst = 32'h10408000;
      3010: inst = 32'hc40452e;
      3011: inst = 32'h8220000;
      3012: inst = 32'h10408000;
      3013: inst = 32'hc40452f;
      3014: inst = 32'h8220000;
      3015: inst = 32'h10408000;
      3016: inst = 32'hc404530;
      3017: inst = 32'h8220000;
      3018: inst = 32'h10408000;
      3019: inst = 32'hc404531;
      3020: inst = 32'h8220000;
      3021: inst = 32'h10408000;
      3022: inst = 32'hc404532;
      3023: inst = 32'h8220000;
      3024: inst = 32'h10408000;
      3025: inst = 32'hc404533;
      3026: inst = 32'h8220000;
      3027: inst = 32'h10408000;
      3028: inst = 32'hc404534;
      3029: inst = 32'h8220000;
      3030: inst = 32'h10408000;
      3031: inst = 32'hc404535;
      3032: inst = 32'h8220000;
      3033: inst = 32'h10408000;
      3034: inst = 32'hc404536;
      3035: inst = 32'h8220000;
      3036: inst = 32'h10408000;
      3037: inst = 32'hc404537;
      3038: inst = 32'h8220000;
      3039: inst = 32'h10408000;
      3040: inst = 32'hc404538;
      3041: inst = 32'h8220000;
      3042: inst = 32'h10408000;
      3043: inst = 32'hc404539;
      3044: inst = 32'h8220000;
      3045: inst = 32'h10408000;
      3046: inst = 32'hc40453a;
      3047: inst = 32'h8220000;
      3048: inst = 32'h10408000;
      3049: inst = 32'hc40453b;
      3050: inst = 32'h8220000;
      3051: inst = 32'h10408000;
      3052: inst = 32'hc404564;
      3053: inst = 32'h8220000;
      3054: inst = 32'h10408000;
      3055: inst = 32'hc404565;
      3056: inst = 32'h8220000;
      3057: inst = 32'h10408000;
      3058: inst = 32'hc404566;
      3059: inst = 32'h8220000;
      3060: inst = 32'h10408000;
      3061: inst = 32'hc404567;
      3062: inst = 32'h8220000;
      3063: inst = 32'h10408000;
      3064: inst = 32'hc404568;
      3065: inst = 32'h8220000;
      3066: inst = 32'h10408000;
      3067: inst = 32'hc404569;
      3068: inst = 32'h8220000;
      3069: inst = 32'h10408000;
      3070: inst = 32'hc40456a;
      3071: inst = 32'h8220000;
      3072: inst = 32'h10408000;
      3073: inst = 32'hc40456b;
      3074: inst = 32'h8220000;
      3075: inst = 32'h10408000;
      3076: inst = 32'hc40456c;
      3077: inst = 32'h8220000;
      3078: inst = 32'h10408000;
      3079: inst = 32'hc40456d;
      3080: inst = 32'h8220000;
      3081: inst = 32'h10408000;
      3082: inst = 32'hc40456e;
      3083: inst = 32'h8220000;
      3084: inst = 32'h10408000;
      3085: inst = 32'hc40456f;
      3086: inst = 32'h8220000;
      3087: inst = 32'h10408000;
      3088: inst = 32'hc404570;
      3089: inst = 32'h8220000;
      3090: inst = 32'h10408000;
      3091: inst = 32'hc404571;
      3092: inst = 32'h8220000;
      3093: inst = 32'h10408000;
      3094: inst = 32'hc404572;
      3095: inst = 32'h8220000;
      3096: inst = 32'h10408000;
      3097: inst = 32'hc404573;
      3098: inst = 32'h8220000;
      3099: inst = 32'h10408000;
      3100: inst = 32'hc404574;
      3101: inst = 32'h8220000;
      3102: inst = 32'h10408000;
      3103: inst = 32'hc404575;
      3104: inst = 32'h8220000;
      3105: inst = 32'h10408000;
      3106: inst = 32'hc404576;
      3107: inst = 32'h8220000;
      3108: inst = 32'h10408000;
      3109: inst = 32'hc404577;
      3110: inst = 32'h8220000;
      3111: inst = 32'h10408000;
      3112: inst = 32'hc404578;
      3113: inst = 32'h8220000;
      3114: inst = 32'h10408000;
      3115: inst = 32'hc404579;
      3116: inst = 32'h8220000;
      3117: inst = 32'h10408000;
      3118: inst = 32'hc40457a;
      3119: inst = 32'h8220000;
      3120: inst = 32'h10408000;
      3121: inst = 32'hc40457b;
      3122: inst = 32'h8220000;
      3123: inst = 32'h10408000;
      3124: inst = 32'hc40457c;
      3125: inst = 32'h8220000;
      3126: inst = 32'h10408000;
      3127: inst = 32'hc40457d;
      3128: inst = 32'h8220000;
      3129: inst = 32'h10408000;
      3130: inst = 32'hc40457e;
      3131: inst = 32'h8220000;
      3132: inst = 32'h10408000;
      3133: inst = 32'hc40457f;
      3134: inst = 32'h8220000;
      3135: inst = 32'h10408000;
      3136: inst = 32'hc404580;
      3137: inst = 32'h8220000;
      3138: inst = 32'h10408000;
      3139: inst = 32'hc404581;
      3140: inst = 32'h8220000;
      3141: inst = 32'h10408000;
      3142: inst = 32'hc404582;
      3143: inst = 32'h8220000;
      3144: inst = 32'h10408000;
      3145: inst = 32'hc404583;
      3146: inst = 32'h8220000;
      3147: inst = 32'h10408000;
      3148: inst = 32'hc404584;
      3149: inst = 32'h8220000;
      3150: inst = 32'h10408000;
      3151: inst = 32'hc404585;
      3152: inst = 32'h8220000;
      3153: inst = 32'h10408000;
      3154: inst = 32'hc404586;
      3155: inst = 32'h8220000;
      3156: inst = 32'h10408000;
      3157: inst = 32'hc404587;
      3158: inst = 32'h8220000;
      3159: inst = 32'h10408000;
      3160: inst = 32'hc404588;
      3161: inst = 32'h8220000;
      3162: inst = 32'h10408000;
      3163: inst = 32'hc404589;
      3164: inst = 32'h8220000;
      3165: inst = 32'h10408000;
      3166: inst = 32'hc40458a;
      3167: inst = 32'h8220000;
      3168: inst = 32'h10408000;
      3169: inst = 32'hc40458b;
      3170: inst = 32'h8220000;
      3171: inst = 32'h10408000;
      3172: inst = 32'hc40458c;
      3173: inst = 32'h8220000;
      3174: inst = 32'h10408000;
      3175: inst = 32'hc40458d;
      3176: inst = 32'h8220000;
      3177: inst = 32'h10408000;
      3178: inst = 32'hc40458e;
      3179: inst = 32'h8220000;
      3180: inst = 32'h10408000;
      3181: inst = 32'hc40458f;
      3182: inst = 32'h8220000;
      3183: inst = 32'h10408000;
      3184: inst = 32'hc404590;
      3185: inst = 32'h8220000;
      3186: inst = 32'h10408000;
      3187: inst = 32'hc404591;
      3188: inst = 32'h8220000;
      3189: inst = 32'h10408000;
      3190: inst = 32'hc404592;
      3191: inst = 32'h8220000;
      3192: inst = 32'h10408000;
      3193: inst = 32'hc404593;
      3194: inst = 32'h8220000;
      3195: inst = 32'h10408000;
      3196: inst = 32'hc404594;
      3197: inst = 32'h8220000;
      3198: inst = 32'h10408000;
      3199: inst = 32'hc404595;
      3200: inst = 32'h8220000;
      3201: inst = 32'h10408000;
      3202: inst = 32'hc404596;
      3203: inst = 32'h8220000;
      3204: inst = 32'h10408000;
      3205: inst = 32'hc404597;
      3206: inst = 32'h8220000;
      3207: inst = 32'h10408000;
      3208: inst = 32'hc404598;
      3209: inst = 32'h8220000;
      3210: inst = 32'h10408000;
      3211: inst = 32'hc404599;
      3212: inst = 32'h8220000;
      3213: inst = 32'h10408000;
      3214: inst = 32'hc40459a;
      3215: inst = 32'h8220000;
      3216: inst = 32'h10408000;
      3217: inst = 32'hc40459b;
      3218: inst = 32'h8220000;
      3219: inst = 32'h10408000;
      3220: inst = 32'hc4045c4;
      3221: inst = 32'h8220000;
      3222: inst = 32'h10408000;
      3223: inst = 32'hc4045c5;
      3224: inst = 32'h8220000;
      3225: inst = 32'h10408000;
      3226: inst = 32'hc4045c6;
      3227: inst = 32'h8220000;
      3228: inst = 32'h10408000;
      3229: inst = 32'hc4045c7;
      3230: inst = 32'h8220000;
      3231: inst = 32'h10408000;
      3232: inst = 32'hc4045c8;
      3233: inst = 32'h8220000;
      3234: inst = 32'h10408000;
      3235: inst = 32'hc4045c9;
      3236: inst = 32'h8220000;
      3237: inst = 32'h10408000;
      3238: inst = 32'hc4045ca;
      3239: inst = 32'h8220000;
      3240: inst = 32'h10408000;
      3241: inst = 32'hc4045cb;
      3242: inst = 32'h8220000;
      3243: inst = 32'h10408000;
      3244: inst = 32'hc4045cc;
      3245: inst = 32'h8220000;
      3246: inst = 32'h10408000;
      3247: inst = 32'hc4045cd;
      3248: inst = 32'h8220000;
      3249: inst = 32'h10408000;
      3250: inst = 32'hc4045ce;
      3251: inst = 32'h8220000;
      3252: inst = 32'h10408000;
      3253: inst = 32'hc4045cf;
      3254: inst = 32'h8220000;
      3255: inst = 32'h10408000;
      3256: inst = 32'hc4045d0;
      3257: inst = 32'h8220000;
      3258: inst = 32'h10408000;
      3259: inst = 32'hc4045d1;
      3260: inst = 32'h8220000;
      3261: inst = 32'h10408000;
      3262: inst = 32'hc4045d2;
      3263: inst = 32'h8220000;
      3264: inst = 32'h10408000;
      3265: inst = 32'hc4045d3;
      3266: inst = 32'h8220000;
      3267: inst = 32'h10408000;
      3268: inst = 32'hc4045d4;
      3269: inst = 32'h8220000;
      3270: inst = 32'h10408000;
      3271: inst = 32'hc4045d5;
      3272: inst = 32'h8220000;
      3273: inst = 32'h10408000;
      3274: inst = 32'hc4045d6;
      3275: inst = 32'h8220000;
      3276: inst = 32'h10408000;
      3277: inst = 32'hc4045d7;
      3278: inst = 32'h8220000;
      3279: inst = 32'h10408000;
      3280: inst = 32'hc4045d8;
      3281: inst = 32'h8220000;
      3282: inst = 32'h10408000;
      3283: inst = 32'hc4045d9;
      3284: inst = 32'h8220000;
      3285: inst = 32'h10408000;
      3286: inst = 32'hc4045da;
      3287: inst = 32'h8220000;
      3288: inst = 32'h10408000;
      3289: inst = 32'hc4045db;
      3290: inst = 32'h8220000;
      3291: inst = 32'h10408000;
      3292: inst = 32'hc4045dc;
      3293: inst = 32'h8220000;
      3294: inst = 32'h10408000;
      3295: inst = 32'hc4045dd;
      3296: inst = 32'h8220000;
      3297: inst = 32'h10408000;
      3298: inst = 32'hc4045de;
      3299: inst = 32'h8220000;
      3300: inst = 32'h10408000;
      3301: inst = 32'hc4045df;
      3302: inst = 32'h8220000;
      3303: inst = 32'h10408000;
      3304: inst = 32'hc4045e0;
      3305: inst = 32'h8220000;
      3306: inst = 32'h10408000;
      3307: inst = 32'hc4045e1;
      3308: inst = 32'h8220000;
      3309: inst = 32'h10408000;
      3310: inst = 32'hc4045e2;
      3311: inst = 32'h8220000;
      3312: inst = 32'h10408000;
      3313: inst = 32'hc4045e3;
      3314: inst = 32'h8220000;
      3315: inst = 32'h10408000;
      3316: inst = 32'hc4045e4;
      3317: inst = 32'h8220000;
      3318: inst = 32'h10408000;
      3319: inst = 32'hc4045e5;
      3320: inst = 32'h8220000;
      3321: inst = 32'h10408000;
      3322: inst = 32'hc4045e6;
      3323: inst = 32'h8220000;
      3324: inst = 32'h10408000;
      3325: inst = 32'hc4045e7;
      3326: inst = 32'h8220000;
      3327: inst = 32'h10408000;
      3328: inst = 32'hc4045e8;
      3329: inst = 32'h8220000;
      3330: inst = 32'h10408000;
      3331: inst = 32'hc4045e9;
      3332: inst = 32'h8220000;
      3333: inst = 32'h10408000;
      3334: inst = 32'hc4045ea;
      3335: inst = 32'h8220000;
      3336: inst = 32'h10408000;
      3337: inst = 32'hc4045eb;
      3338: inst = 32'h8220000;
      3339: inst = 32'h10408000;
      3340: inst = 32'hc4045ec;
      3341: inst = 32'h8220000;
      3342: inst = 32'h10408000;
      3343: inst = 32'hc4045ed;
      3344: inst = 32'h8220000;
      3345: inst = 32'h10408000;
      3346: inst = 32'hc4045ee;
      3347: inst = 32'h8220000;
      3348: inst = 32'h10408000;
      3349: inst = 32'hc4045ef;
      3350: inst = 32'h8220000;
      3351: inst = 32'h10408000;
      3352: inst = 32'hc4045f0;
      3353: inst = 32'h8220000;
      3354: inst = 32'h10408000;
      3355: inst = 32'hc4045f1;
      3356: inst = 32'h8220000;
      3357: inst = 32'h10408000;
      3358: inst = 32'hc4045f2;
      3359: inst = 32'h8220000;
      3360: inst = 32'h10408000;
      3361: inst = 32'hc4045f3;
      3362: inst = 32'h8220000;
      3363: inst = 32'h10408000;
      3364: inst = 32'hc4045f4;
      3365: inst = 32'h8220000;
      3366: inst = 32'h10408000;
      3367: inst = 32'hc4045f5;
      3368: inst = 32'h8220000;
      3369: inst = 32'h10408000;
      3370: inst = 32'hc4045f6;
      3371: inst = 32'h8220000;
      3372: inst = 32'h10408000;
      3373: inst = 32'hc4045f7;
      3374: inst = 32'h8220000;
      3375: inst = 32'h10408000;
      3376: inst = 32'hc4045f8;
      3377: inst = 32'h8220000;
      3378: inst = 32'h10408000;
      3379: inst = 32'hc4045f9;
      3380: inst = 32'h8220000;
      3381: inst = 32'h10408000;
      3382: inst = 32'hc4045fa;
      3383: inst = 32'h8220000;
      3384: inst = 32'h10408000;
      3385: inst = 32'hc4045fb;
      3386: inst = 32'h8220000;
      3387: inst = 32'h10408000;
      3388: inst = 32'hc404624;
      3389: inst = 32'h8220000;
      3390: inst = 32'h10408000;
      3391: inst = 32'hc404625;
      3392: inst = 32'h8220000;
      3393: inst = 32'h10408000;
      3394: inst = 32'hc404626;
      3395: inst = 32'h8220000;
      3396: inst = 32'h10408000;
      3397: inst = 32'hc404627;
      3398: inst = 32'h8220000;
      3399: inst = 32'h10408000;
      3400: inst = 32'hc404628;
      3401: inst = 32'h8220000;
      3402: inst = 32'h10408000;
      3403: inst = 32'hc404629;
      3404: inst = 32'h8220000;
      3405: inst = 32'h10408000;
      3406: inst = 32'hc40462a;
      3407: inst = 32'h8220000;
      3408: inst = 32'h10408000;
      3409: inst = 32'hc40462b;
      3410: inst = 32'h8220000;
      3411: inst = 32'h10408000;
      3412: inst = 32'hc40462c;
      3413: inst = 32'h8220000;
      3414: inst = 32'h10408000;
      3415: inst = 32'hc40462d;
      3416: inst = 32'h8220000;
      3417: inst = 32'h10408000;
      3418: inst = 32'hc40462e;
      3419: inst = 32'h8220000;
      3420: inst = 32'h10408000;
      3421: inst = 32'hc40462f;
      3422: inst = 32'h8220000;
      3423: inst = 32'h10408000;
      3424: inst = 32'hc404630;
      3425: inst = 32'h8220000;
      3426: inst = 32'h10408000;
      3427: inst = 32'hc404631;
      3428: inst = 32'h8220000;
      3429: inst = 32'h10408000;
      3430: inst = 32'hc404632;
      3431: inst = 32'h8220000;
      3432: inst = 32'h10408000;
      3433: inst = 32'hc404633;
      3434: inst = 32'h8220000;
      3435: inst = 32'h10408000;
      3436: inst = 32'hc404634;
      3437: inst = 32'h8220000;
      3438: inst = 32'h10408000;
      3439: inst = 32'hc404635;
      3440: inst = 32'h8220000;
      3441: inst = 32'h10408000;
      3442: inst = 32'hc404636;
      3443: inst = 32'h8220000;
      3444: inst = 32'h10408000;
      3445: inst = 32'hc404637;
      3446: inst = 32'h8220000;
      3447: inst = 32'h10408000;
      3448: inst = 32'hc404638;
      3449: inst = 32'h8220000;
      3450: inst = 32'h10408000;
      3451: inst = 32'hc404639;
      3452: inst = 32'h8220000;
      3453: inst = 32'h10408000;
      3454: inst = 32'hc40463a;
      3455: inst = 32'h8220000;
      3456: inst = 32'h10408000;
      3457: inst = 32'hc40463b;
      3458: inst = 32'h8220000;
      3459: inst = 32'h10408000;
      3460: inst = 32'hc40463c;
      3461: inst = 32'h8220000;
      3462: inst = 32'h10408000;
      3463: inst = 32'hc40463d;
      3464: inst = 32'h8220000;
      3465: inst = 32'h10408000;
      3466: inst = 32'hc40463e;
      3467: inst = 32'h8220000;
      3468: inst = 32'h10408000;
      3469: inst = 32'hc40463f;
      3470: inst = 32'h8220000;
      3471: inst = 32'h10408000;
      3472: inst = 32'hc404640;
      3473: inst = 32'h8220000;
      3474: inst = 32'h10408000;
      3475: inst = 32'hc404641;
      3476: inst = 32'h8220000;
      3477: inst = 32'h10408000;
      3478: inst = 32'hc404642;
      3479: inst = 32'h8220000;
      3480: inst = 32'h10408000;
      3481: inst = 32'hc404643;
      3482: inst = 32'h8220000;
      3483: inst = 32'h10408000;
      3484: inst = 32'hc404644;
      3485: inst = 32'h8220000;
      3486: inst = 32'h10408000;
      3487: inst = 32'hc404645;
      3488: inst = 32'h8220000;
      3489: inst = 32'h10408000;
      3490: inst = 32'hc404646;
      3491: inst = 32'h8220000;
      3492: inst = 32'h10408000;
      3493: inst = 32'hc404647;
      3494: inst = 32'h8220000;
      3495: inst = 32'h10408000;
      3496: inst = 32'hc404648;
      3497: inst = 32'h8220000;
      3498: inst = 32'h10408000;
      3499: inst = 32'hc404649;
      3500: inst = 32'h8220000;
      3501: inst = 32'h10408000;
      3502: inst = 32'hc40464a;
      3503: inst = 32'h8220000;
      3504: inst = 32'h10408000;
      3505: inst = 32'hc40464b;
      3506: inst = 32'h8220000;
      3507: inst = 32'h10408000;
      3508: inst = 32'hc40464c;
      3509: inst = 32'h8220000;
      3510: inst = 32'h10408000;
      3511: inst = 32'hc40464d;
      3512: inst = 32'h8220000;
      3513: inst = 32'h10408000;
      3514: inst = 32'hc40464e;
      3515: inst = 32'h8220000;
      3516: inst = 32'h10408000;
      3517: inst = 32'hc40464f;
      3518: inst = 32'h8220000;
      3519: inst = 32'h10408000;
      3520: inst = 32'hc404650;
      3521: inst = 32'h8220000;
      3522: inst = 32'h10408000;
      3523: inst = 32'hc404651;
      3524: inst = 32'h8220000;
      3525: inst = 32'h10408000;
      3526: inst = 32'hc404652;
      3527: inst = 32'h8220000;
      3528: inst = 32'h10408000;
      3529: inst = 32'hc404653;
      3530: inst = 32'h8220000;
      3531: inst = 32'h10408000;
      3532: inst = 32'hc404654;
      3533: inst = 32'h8220000;
      3534: inst = 32'h10408000;
      3535: inst = 32'hc404655;
      3536: inst = 32'h8220000;
      3537: inst = 32'h10408000;
      3538: inst = 32'hc404656;
      3539: inst = 32'h8220000;
      3540: inst = 32'h10408000;
      3541: inst = 32'hc404657;
      3542: inst = 32'h8220000;
      3543: inst = 32'h10408000;
      3544: inst = 32'hc404658;
      3545: inst = 32'h8220000;
      3546: inst = 32'h10408000;
      3547: inst = 32'hc404659;
      3548: inst = 32'h8220000;
      3549: inst = 32'h10408000;
      3550: inst = 32'hc40465a;
      3551: inst = 32'h8220000;
      3552: inst = 32'h10408000;
      3553: inst = 32'hc40465b;
      3554: inst = 32'h8220000;
      3555: inst = 32'h10408000;
      3556: inst = 32'hc404684;
      3557: inst = 32'h8220000;
      3558: inst = 32'h10408000;
      3559: inst = 32'hc404685;
      3560: inst = 32'h8220000;
      3561: inst = 32'h10408000;
      3562: inst = 32'hc404686;
      3563: inst = 32'h8220000;
      3564: inst = 32'h10408000;
      3565: inst = 32'hc404687;
      3566: inst = 32'h8220000;
      3567: inst = 32'h10408000;
      3568: inst = 32'hc404688;
      3569: inst = 32'h8220000;
      3570: inst = 32'h10408000;
      3571: inst = 32'hc404689;
      3572: inst = 32'h8220000;
      3573: inst = 32'h10408000;
      3574: inst = 32'hc40468a;
      3575: inst = 32'h8220000;
      3576: inst = 32'h10408000;
      3577: inst = 32'hc40468b;
      3578: inst = 32'h8220000;
      3579: inst = 32'h10408000;
      3580: inst = 32'hc40468c;
      3581: inst = 32'h8220000;
      3582: inst = 32'h10408000;
      3583: inst = 32'hc40468d;
      3584: inst = 32'h8220000;
      3585: inst = 32'h10408000;
      3586: inst = 32'hc40468e;
      3587: inst = 32'h8220000;
      3588: inst = 32'h10408000;
      3589: inst = 32'hc40468f;
      3590: inst = 32'h8220000;
      3591: inst = 32'h10408000;
      3592: inst = 32'hc404690;
      3593: inst = 32'h8220000;
      3594: inst = 32'h10408000;
      3595: inst = 32'hc404691;
      3596: inst = 32'h8220000;
      3597: inst = 32'h10408000;
      3598: inst = 32'hc404692;
      3599: inst = 32'h8220000;
      3600: inst = 32'h10408000;
      3601: inst = 32'hc404693;
      3602: inst = 32'h8220000;
      3603: inst = 32'h10408000;
      3604: inst = 32'hc404694;
      3605: inst = 32'h8220000;
      3606: inst = 32'h10408000;
      3607: inst = 32'hc404695;
      3608: inst = 32'h8220000;
      3609: inst = 32'h10408000;
      3610: inst = 32'hc404696;
      3611: inst = 32'h8220000;
      3612: inst = 32'h10408000;
      3613: inst = 32'hc404697;
      3614: inst = 32'h8220000;
      3615: inst = 32'h10408000;
      3616: inst = 32'hc404698;
      3617: inst = 32'h8220000;
      3618: inst = 32'h10408000;
      3619: inst = 32'hc404699;
      3620: inst = 32'h8220000;
      3621: inst = 32'h10408000;
      3622: inst = 32'hc40469a;
      3623: inst = 32'h8220000;
      3624: inst = 32'h10408000;
      3625: inst = 32'hc40469b;
      3626: inst = 32'h8220000;
      3627: inst = 32'h10408000;
      3628: inst = 32'hc40469c;
      3629: inst = 32'h8220000;
      3630: inst = 32'h10408000;
      3631: inst = 32'hc40469d;
      3632: inst = 32'h8220000;
      3633: inst = 32'h10408000;
      3634: inst = 32'hc40469e;
      3635: inst = 32'h8220000;
      3636: inst = 32'h10408000;
      3637: inst = 32'hc40469f;
      3638: inst = 32'h8220000;
      3639: inst = 32'h10408000;
      3640: inst = 32'hc4046a0;
      3641: inst = 32'h8220000;
      3642: inst = 32'h10408000;
      3643: inst = 32'hc4046a1;
      3644: inst = 32'h8220000;
      3645: inst = 32'h10408000;
      3646: inst = 32'hc4046a2;
      3647: inst = 32'h8220000;
      3648: inst = 32'h10408000;
      3649: inst = 32'hc4046a3;
      3650: inst = 32'h8220000;
      3651: inst = 32'h10408000;
      3652: inst = 32'hc4046a4;
      3653: inst = 32'h8220000;
      3654: inst = 32'h10408000;
      3655: inst = 32'hc4046a5;
      3656: inst = 32'h8220000;
      3657: inst = 32'h10408000;
      3658: inst = 32'hc4046a6;
      3659: inst = 32'h8220000;
      3660: inst = 32'h10408000;
      3661: inst = 32'hc4046a7;
      3662: inst = 32'h8220000;
      3663: inst = 32'h10408000;
      3664: inst = 32'hc4046a8;
      3665: inst = 32'h8220000;
      3666: inst = 32'h10408000;
      3667: inst = 32'hc4046a9;
      3668: inst = 32'h8220000;
      3669: inst = 32'h10408000;
      3670: inst = 32'hc4046aa;
      3671: inst = 32'h8220000;
      3672: inst = 32'h10408000;
      3673: inst = 32'hc4046ab;
      3674: inst = 32'h8220000;
      3675: inst = 32'h10408000;
      3676: inst = 32'hc4046ac;
      3677: inst = 32'h8220000;
      3678: inst = 32'h10408000;
      3679: inst = 32'hc4046ad;
      3680: inst = 32'h8220000;
      3681: inst = 32'h10408000;
      3682: inst = 32'hc4046ae;
      3683: inst = 32'h8220000;
      3684: inst = 32'h10408000;
      3685: inst = 32'hc4046af;
      3686: inst = 32'h8220000;
      3687: inst = 32'h10408000;
      3688: inst = 32'hc4046b0;
      3689: inst = 32'h8220000;
      3690: inst = 32'h10408000;
      3691: inst = 32'hc4046b1;
      3692: inst = 32'h8220000;
      3693: inst = 32'h10408000;
      3694: inst = 32'hc4046b2;
      3695: inst = 32'h8220000;
      3696: inst = 32'h10408000;
      3697: inst = 32'hc4046b3;
      3698: inst = 32'h8220000;
      3699: inst = 32'h10408000;
      3700: inst = 32'hc4046b4;
      3701: inst = 32'h8220000;
      3702: inst = 32'h10408000;
      3703: inst = 32'hc4046b5;
      3704: inst = 32'h8220000;
      3705: inst = 32'h10408000;
      3706: inst = 32'hc4046b6;
      3707: inst = 32'h8220000;
      3708: inst = 32'h10408000;
      3709: inst = 32'hc4046b7;
      3710: inst = 32'h8220000;
      3711: inst = 32'h10408000;
      3712: inst = 32'hc4046b8;
      3713: inst = 32'h8220000;
      3714: inst = 32'h10408000;
      3715: inst = 32'hc4046b9;
      3716: inst = 32'h8220000;
      3717: inst = 32'h10408000;
      3718: inst = 32'hc4046ba;
      3719: inst = 32'h8220000;
      3720: inst = 32'h10408000;
      3721: inst = 32'hc4046bb;
      3722: inst = 32'h8220000;
      3723: inst = 32'h10408000;
      3724: inst = 32'hc4046e4;
      3725: inst = 32'h8220000;
      3726: inst = 32'h10408000;
      3727: inst = 32'hc4046e5;
      3728: inst = 32'h8220000;
      3729: inst = 32'h10408000;
      3730: inst = 32'hc4046e6;
      3731: inst = 32'h8220000;
      3732: inst = 32'h10408000;
      3733: inst = 32'hc4046e7;
      3734: inst = 32'h8220000;
      3735: inst = 32'h10408000;
      3736: inst = 32'hc4046e8;
      3737: inst = 32'h8220000;
      3738: inst = 32'h10408000;
      3739: inst = 32'hc4046e9;
      3740: inst = 32'h8220000;
      3741: inst = 32'h10408000;
      3742: inst = 32'hc4046ea;
      3743: inst = 32'h8220000;
      3744: inst = 32'h10408000;
      3745: inst = 32'hc4046eb;
      3746: inst = 32'h8220000;
      3747: inst = 32'h10408000;
      3748: inst = 32'hc4046ec;
      3749: inst = 32'h8220000;
      3750: inst = 32'h10408000;
      3751: inst = 32'hc4046ed;
      3752: inst = 32'h8220000;
      3753: inst = 32'h10408000;
      3754: inst = 32'hc4046ee;
      3755: inst = 32'h8220000;
      3756: inst = 32'h10408000;
      3757: inst = 32'hc404700;
      3758: inst = 32'h8220000;
      3759: inst = 32'h10408000;
      3760: inst = 32'hc404701;
      3761: inst = 32'h8220000;
      3762: inst = 32'h10408000;
      3763: inst = 32'hc404702;
      3764: inst = 32'h8220000;
      3765: inst = 32'h10408000;
      3766: inst = 32'hc404703;
      3767: inst = 32'h8220000;
      3768: inst = 32'h10408000;
      3769: inst = 32'hc404704;
      3770: inst = 32'h8220000;
      3771: inst = 32'h10408000;
      3772: inst = 32'hc404705;
      3773: inst = 32'h8220000;
      3774: inst = 32'h10408000;
      3775: inst = 32'hc404706;
      3776: inst = 32'h8220000;
      3777: inst = 32'h10408000;
      3778: inst = 32'hc404707;
      3779: inst = 32'h8220000;
      3780: inst = 32'h10408000;
      3781: inst = 32'hc404708;
      3782: inst = 32'h8220000;
      3783: inst = 32'h10408000;
      3784: inst = 32'hc404709;
      3785: inst = 32'h8220000;
      3786: inst = 32'h10408000;
      3787: inst = 32'hc40470a;
      3788: inst = 32'h8220000;
      3789: inst = 32'h10408000;
      3790: inst = 32'hc40470b;
      3791: inst = 32'h8220000;
      3792: inst = 32'h10408000;
      3793: inst = 32'hc40470c;
      3794: inst = 32'h8220000;
      3795: inst = 32'h10408000;
      3796: inst = 32'hc40470d;
      3797: inst = 32'h8220000;
      3798: inst = 32'h10408000;
      3799: inst = 32'hc40470e;
      3800: inst = 32'h8220000;
      3801: inst = 32'h10408000;
      3802: inst = 32'hc40470f;
      3803: inst = 32'h8220000;
      3804: inst = 32'h10408000;
      3805: inst = 32'hc404710;
      3806: inst = 32'h8220000;
      3807: inst = 32'h10408000;
      3808: inst = 32'hc404711;
      3809: inst = 32'h8220000;
      3810: inst = 32'h10408000;
      3811: inst = 32'hc404712;
      3812: inst = 32'h8220000;
      3813: inst = 32'h10408000;
      3814: inst = 32'hc404713;
      3815: inst = 32'h8220000;
      3816: inst = 32'h10408000;
      3817: inst = 32'hc404714;
      3818: inst = 32'h8220000;
      3819: inst = 32'h10408000;
      3820: inst = 32'hc404715;
      3821: inst = 32'h8220000;
      3822: inst = 32'h10408000;
      3823: inst = 32'hc404716;
      3824: inst = 32'h8220000;
      3825: inst = 32'h10408000;
      3826: inst = 32'hc404717;
      3827: inst = 32'h8220000;
      3828: inst = 32'h10408000;
      3829: inst = 32'hc404718;
      3830: inst = 32'h8220000;
      3831: inst = 32'h10408000;
      3832: inst = 32'hc404719;
      3833: inst = 32'h8220000;
      3834: inst = 32'h10408000;
      3835: inst = 32'hc40471a;
      3836: inst = 32'h8220000;
      3837: inst = 32'h10408000;
      3838: inst = 32'hc40471b;
      3839: inst = 32'h8220000;
      3840: inst = 32'h10408000;
      3841: inst = 32'hc404744;
      3842: inst = 32'h8220000;
      3843: inst = 32'h10408000;
      3844: inst = 32'hc404745;
      3845: inst = 32'h8220000;
      3846: inst = 32'h10408000;
      3847: inst = 32'hc404746;
      3848: inst = 32'h8220000;
      3849: inst = 32'h10408000;
      3850: inst = 32'hc404747;
      3851: inst = 32'h8220000;
      3852: inst = 32'h10408000;
      3853: inst = 32'hc404748;
      3854: inst = 32'h8220000;
      3855: inst = 32'h10408000;
      3856: inst = 32'hc404749;
      3857: inst = 32'h8220000;
      3858: inst = 32'h10408000;
      3859: inst = 32'hc40474a;
      3860: inst = 32'h8220000;
      3861: inst = 32'h10408000;
      3862: inst = 32'hc40474b;
      3863: inst = 32'h8220000;
      3864: inst = 32'h10408000;
      3865: inst = 32'hc40474c;
      3866: inst = 32'h8220000;
      3867: inst = 32'h10408000;
      3868: inst = 32'hc40474d;
      3869: inst = 32'h8220000;
      3870: inst = 32'h10408000;
      3871: inst = 32'hc40474e;
      3872: inst = 32'h8220000;
      3873: inst = 32'h10408000;
      3874: inst = 32'hc404760;
      3875: inst = 32'h8220000;
      3876: inst = 32'h10408000;
      3877: inst = 32'hc404761;
      3878: inst = 32'h8220000;
      3879: inst = 32'h10408000;
      3880: inst = 32'hc404762;
      3881: inst = 32'h8220000;
      3882: inst = 32'h10408000;
      3883: inst = 32'hc404763;
      3884: inst = 32'h8220000;
      3885: inst = 32'h10408000;
      3886: inst = 32'hc404764;
      3887: inst = 32'h8220000;
      3888: inst = 32'h10408000;
      3889: inst = 32'hc404765;
      3890: inst = 32'h8220000;
      3891: inst = 32'h10408000;
      3892: inst = 32'hc404766;
      3893: inst = 32'h8220000;
      3894: inst = 32'h10408000;
      3895: inst = 32'hc404767;
      3896: inst = 32'h8220000;
      3897: inst = 32'h10408000;
      3898: inst = 32'hc404768;
      3899: inst = 32'h8220000;
      3900: inst = 32'h10408000;
      3901: inst = 32'hc404769;
      3902: inst = 32'h8220000;
      3903: inst = 32'h10408000;
      3904: inst = 32'hc40476a;
      3905: inst = 32'h8220000;
      3906: inst = 32'h10408000;
      3907: inst = 32'hc40476b;
      3908: inst = 32'h8220000;
      3909: inst = 32'h10408000;
      3910: inst = 32'hc40476c;
      3911: inst = 32'h8220000;
      3912: inst = 32'h10408000;
      3913: inst = 32'hc40476d;
      3914: inst = 32'h8220000;
      3915: inst = 32'h10408000;
      3916: inst = 32'hc40476e;
      3917: inst = 32'h8220000;
      3918: inst = 32'h10408000;
      3919: inst = 32'hc40476f;
      3920: inst = 32'h8220000;
      3921: inst = 32'h10408000;
      3922: inst = 32'hc404770;
      3923: inst = 32'h8220000;
      3924: inst = 32'h10408000;
      3925: inst = 32'hc404771;
      3926: inst = 32'h8220000;
      3927: inst = 32'h10408000;
      3928: inst = 32'hc404772;
      3929: inst = 32'h8220000;
      3930: inst = 32'h10408000;
      3931: inst = 32'hc404773;
      3932: inst = 32'h8220000;
      3933: inst = 32'h10408000;
      3934: inst = 32'hc404774;
      3935: inst = 32'h8220000;
      3936: inst = 32'h10408000;
      3937: inst = 32'hc404775;
      3938: inst = 32'h8220000;
      3939: inst = 32'h10408000;
      3940: inst = 32'hc404776;
      3941: inst = 32'h8220000;
      3942: inst = 32'h10408000;
      3943: inst = 32'hc404777;
      3944: inst = 32'h8220000;
      3945: inst = 32'h10408000;
      3946: inst = 32'hc404778;
      3947: inst = 32'h8220000;
      3948: inst = 32'h10408000;
      3949: inst = 32'hc404779;
      3950: inst = 32'h8220000;
      3951: inst = 32'h10408000;
      3952: inst = 32'hc40477a;
      3953: inst = 32'h8220000;
      3954: inst = 32'h10408000;
      3955: inst = 32'hc40477b;
      3956: inst = 32'h8220000;
      3957: inst = 32'h10408000;
      3958: inst = 32'hc4047a4;
      3959: inst = 32'h8220000;
      3960: inst = 32'h10408000;
      3961: inst = 32'hc4047a5;
      3962: inst = 32'h8220000;
      3963: inst = 32'h10408000;
      3964: inst = 32'hc4047a6;
      3965: inst = 32'h8220000;
      3966: inst = 32'h10408000;
      3967: inst = 32'hc4047a7;
      3968: inst = 32'h8220000;
      3969: inst = 32'h10408000;
      3970: inst = 32'hc4047a8;
      3971: inst = 32'h8220000;
      3972: inst = 32'h10408000;
      3973: inst = 32'hc4047a9;
      3974: inst = 32'h8220000;
      3975: inst = 32'h10408000;
      3976: inst = 32'hc4047aa;
      3977: inst = 32'h8220000;
      3978: inst = 32'h10408000;
      3979: inst = 32'hc4047ab;
      3980: inst = 32'h8220000;
      3981: inst = 32'h10408000;
      3982: inst = 32'hc4047ac;
      3983: inst = 32'h8220000;
      3984: inst = 32'h10408000;
      3985: inst = 32'hc4047ad;
      3986: inst = 32'h8220000;
      3987: inst = 32'h10408000;
      3988: inst = 32'hc4047ae;
      3989: inst = 32'h8220000;
      3990: inst = 32'h10408000;
      3991: inst = 32'hc4047c0;
      3992: inst = 32'h8220000;
      3993: inst = 32'h10408000;
      3994: inst = 32'hc4047c1;
      3995: inst = 32'h8220000;
      3996: inst = 32'h10408000;
      3997: inst = 32'hc4047c2;
      3998: inst = 32'h8220000;
      3999: inst = 32'h10408000;
      4000: inst = 32'hc4047c3;
      4001: inst = 32'h8220000;
      4002: inst = 32'h10408000;
      4003: inst = 32'hc4047c4;
      4004: inst = 32'h8220000;
      4005: inst = 32'h10408000;
      4006: inst = 32'hc4047c5;
      4007: inst = 32'h8220000;
      4008: inst = 32'h10408000;
      4009: inst = 32'hc4047c6;
      4010: inst = 32'h8220000;
      4011: inst = 32'h10408000;
      4012: inst = 32'hc4047c7;
      4013: inst = 32'h8220000;
      4014: inst = 32'h10408000;
      4015: inst = 32'hc4047c8;
      4016: inst = 32'h8220000;
      4017: inst = 32'h10408000;
      4018: inst = 32'hc4047c9;
      4019: inst = 32'h8220000;
      4020: inst = 32'h10408000;
      4021: inst = 32'hc4047ca;
      4022: inst = 32'h8220000;
      4023: inst = 32'h10408000;
      4024: inst = 32'hc4047cb;
      4025: inst = 32'h8220000;
      4026: inst = 32'h10408000;
      4027: inst = 32'hc4047cc;
      4028: inst = 32'h8220000;
      4029: inst = 32'h10408000;
      4030: inst = 32'hc4047cd;
      4031: inst = 32'h8220000;
      4032: inst = 32'h10408000;
      4033: inst = 32'hc4047ce;
      4034: inst = 32'h8220000;
      4035: inst = 32'h10408000;
      4036: inst = 32'hc4047cf;
      4037: inst = 32'h8220000;
      4038: inst = 32'h10408000;
      4039: inst = 32'hc4047d0;
      4040: inst = 32'h8220000;
      4041: inst = 32'h10408000;
      4042: inst = 32'hc4047d1;
      4043: inst = 32'h8220000;
      4044: inst = 32'h10408000;
      4045: inst = 32'hc4047d2;
      4046: inst = 32'h8220000;
      4047: inst = 32'h10408000;
      4048: inst = 32'hc4047d3;
      4049: inst = 32'h8220000;
      4050: inst = 32'h10408000;
      4051: inst = 32'hc4047d4;
      4052: inst = 32'h8220000;
      4053: inst = 32'h10408000;
      4054: inst = 32'hc4047d5;
      4055: inst = 32'h8220000;
      4056: inst = 32'h10408000;
      4057: inst = 32'hc4047d6;
      4058: inst = 32'h8220000;
      4059: inst = 32'h10408000;
      4060: inst = 32'hc4047d7;
      4061: inst = 32'h8220000;
      4062: inst = 32'h10408000;
      4063: inst = 32'hc4047d8;
      4064: inst = 32'h8220000;
      4065: inst = 32'h10408000;
      4066: inst = 32'hc4047d9;
      4067: inst = 32'h8220000;
      4068: inst = 32'h10408000;
      4069: inst = 32'hc4047da;
      4070: inst = 32'h8220000;
      4071: inst = 32'h10408000;
      4072: inst = 32'hc4047db;
      4073: inst = 32'h8220000;
      4074: inst = 32'h10408000;
      4075: inst = 32'hc404804;
      4076: inst = 32'h8220000;
      4077: inst = 32'h10408000;
      4078: inst = 32'hc404805;
      4079: inst = 32'h8220000;
      4080: inst = 32'h10408000;
      4081: inst = 32'hc404806;
      4082: inst = 32'h8220000;
      4083: inst = 32'h10408000;
      4084: inst = 32'hc404807;
      4085: inst = 32'h8220000;
      4086: inst = 32'h10408000;
      4087: inst = 32'hc404808;
      4088: inst = 32'h8220000;
      4089: inst = 32'h10408000;
      4090: inst = 32'hc404809;
      4091: inst = 32'h8220000;
      4092: inst = 32'h10408000;
      4093: inst = 32'hc40480a;
      4094: inst = 32'h8220000;
      4095: inst = 32'h10408000;
      4096: inst = 32'hc40480b;
      4097: inst = 32'h8220000;
      4098: inst = 32'h10408000;
      4099: inst = 32'hc40480c;
      4100: inst = 32'h8220000;
      4101: inst = 32'h10408000;
      4102: inst = 32'hc40480d;
      4103: inst = 32'h8220000;
      4104: inst = 32'h10408000;
      4105: inst = 32'hc40480e;
      4106: inst = 32'h8220000;
      4107: inst = 32'h10408000;
      4108: inst = 32'hc404820;
      4109: inst = 32'h8220000;
      4110: inst = 32'h10408000;
      4111: inst = 32'hc404821;
      4112: inst = 32'h8220000;
      4113: inst = 32'h10408000;
      4114: inst = 32'hc404822;
      4115: inst = 32'h8220000;
      4116: inst = 32'h10408000;
      4117: inst = 32'hc404823;
      4118: inst = 32'h8220000;
      4119: inst = 32'h10408000;
      4120: inst = 32'hc404824;
      4121: inst = 32'h8220000;
      4122: inst = 32'h10408000;
      4123: inst = 32'hc404825;
      4124: inst = 32'h8220000;
      4125: inst = 32'h10408000;
      4126: inst = 32'hc404826;
      4127: inst = 32'h8220000;
      4128: inst = 32'h10408000;
      4129: inst = 32'hc404827;
      4130: inst = 32'h8220000;
      4131: inst = 32'h10408000;
      4132: inst = 32'hc404828;
      4133: inst = 32'h8220000;
      4134: inst = 32'h10408000;
      4135: inst = 32'hc404829;
      4136: inst = 32'h8220000;
      4137: inst = 32'h10408000;
      4138: inst = 32'hc40482a;
      4139: inst = 32'h8220000;
      4140: inst = 32'h10408000;
      4141: inst = 32'hc40482b;
      4142: inst = 32'h8220000;
      4143: inst = 32'h10408000;
      4144: inst = 32'hc40482c;
      4145: inst = 32'h8220000;
      4146: inst = 32'h10408000;
      4147: inst = 32'hc40482d;
      4148: inst = 32'h8220000;
      4149: inst = 32'h10408000;
      4150: inst = 32'hc40482e;
      4151: inst = 32'h8220000;
      4152: inst = 32'h10408000;
      4153: inst = 32'hc40482f;
      4154: inst = 32'h8220000;
      4155: inst = 32'h10408000;
      4156: inst = 32'hc404830;
      4157: inst = 32'h8220000;
      4158: inst = 32'h10408000;
      4159: inst = 32'hc404831;
      4160: inst = 32'h8220000;
      4161: inst = 32'h10408000;
      4162: inst = 32'hc404832;
      4163: inst = 32'h8220000;
      4164: inst = 32'h10408000;
      4165: inst = 32'hc404833;
      4166: inst = 32'h8220000;
      4167: inst = 32'h10408000;
      4168: inst = 32'hc404834;
      4169: inst = 32'h8220000;
      4170: inst = 32'h10408000;
      4171: inst = 32'hc404835;
      4172: inst = 32'h8220000;
      4173: inst = 32'h10408000;
      4174: inst = 32'hc404836;
      4175: inst = 32'h8220000;
      4176: inst = 32'h10408000;
      4177: inst = 32'hc404837;
      4178: inst = 32'h8220000;
      4179: inst = 32'h10408000;
      4180: inst = 32'hc404838;
      4181: inst = 32'h8220000;
      4182: inst = 32'h10408000;
      4183: inst = 32'hc404839;
      4184: inst = 32'h8220000;
      4185: inst = 32'h10408000;
      4186: inst = 32'hc40483a;
      4187: inst = 32'h8220000;
      4188: inst = 32'h10408000;
      4189: inst = 32'hc40483b;
      4190: inst = 32'h8220000;
      4191: inst = 32'h10408000;
      4192: inst = 32'hc404864;
      4193: inst = 32'h8220000;
      4194: inst = 32'h10408000;
      4195: inst = 32'hc404865;
      4196: inst = 32'h8220000;
      4197: inst = 32'h10408000;
      4198: inst = 32'hc404866;
      4199: inst = 32'h8220000;
      4200: inst = 32'h10408000;
      4201: inst = 32'hc404867;
      4202: inst = 32'h8220000;
      4203: inst = 32'h10408000;
      4204: inst = 32'hc404868;
      4205: inst = 32'h8220000;
      4206: inst = 32'h10408000;
      4207: inst = 32'hc404869;
      4208: inst = 32'h8220000;
      4209: inst = 32'h10408000;
      4210: inst = 32'hc40486a;
      4211: inst = 32'h8220000;
      4212: inst = 32'h10408000;
      4213: inst = 32'hc40486b;
      4214: inst = 32'h8220000;
      4215: inst = 32'h10408000;
      4216: inst = 32'hc40486c;
      4217: inst = 32'h8220000;
      4218: inst = 32'h10408000;
      4219: inst = 32'hc40486d;
      4220: inst = 32'h8220000;
      4221: inst = 32'h10408000;
      4222: inst = 32'hc40486e;
      4223: inst = 32'h8220000;
      4224: inst = 32'h10408000;
      4225: inst = 32'hc404880;
      4226: inst = 32'h8220000;
      4227: inst = 32'h10408000;
      4228: inst = 32'hc404881;
      4229: inst = 32'h8220000;
      4230: inst = 32'h10408000;
      4231: inst = 32'hc404882;
      4232: inst = 32'h8220000;
      4233: inst = 32'h10408000;
      4234: inst = 32'hc404883;
      4235: inst = 32'h8220000;
      4236: inst = 32'h10408000;
      4237: inst = 32'hc404884;
      4238: inst = 32'h8220000;
      4239: inst = 32'h10408000;
      4240: inst = 32'hc404885;
      4241: inst = 32'h8220000;
      4242: inst = 32'h10408000;
      4243: inst = 32'hc404886;
      4244: inst = 32'h8220000;
      4245: inst = 32'h10408000;
      4246: inst = 32'hc404887;
      4247: inst = 32'h8220000;
      4248: inst = 32'h10408000;
      4249: inst = 32'hc404888;
      4250: inst = 32'h8220000;
      4251: inst = 32'h10408000;
      4252: inst = 32'hc404889;
      4253: inst = 32'h8220000;
      4254: inst = 32'h10408000;
      4255: inst = 32'hc40488a;
      4256: inst = 32'h8220000;
      4257: inst = 32'h10408000;
      4258: inst = 32'hc40488b;
      4259: inst = 32'h8220000;
      4260: inst = 32'h10408000;
      4261: inst = 32'hc40488c;
      4262: inst = 32'h8220000;
      4263: inst = 32'h10408000;
      4264: inst = 32'hc40488d;
      4265: inst = 32'h8220000;
      4266: inst = 32'h10408000;
      4267: inst = 32'hc40488e;
      4268: inst = 32'h8220000;
      4269: inst = 32'h10408000;
      4270: inst = 32'hc40488f;
      4271: inst = 32'h8220000;
      4272: inst = 32'h10408000;
      4273: inst = 32'hc404890;
      4274: inst = 32'h8220000;
      4275: inst = 32'h10408000;
      4276: inst = 32'hc404891;
      4277: inst = 32'h8220000;
      4278: inst = 32'h10408000;
      4279: inst = 32'hc404892;
      4280: inst = 32'h8220000;
      4281: inst = 32'h10408000;
      4282: inst = 32'hc404893;
      4283: inst = 32'h8220000;
      4284: inst = 32'h10408000;
      4285: inst = 32'hc404894;
      4286: inst = 32'h8220000;
      4287: inst = 32'h10408000;
      4288: inst = 32'hc404895;
      4289: inst = 32'h8220000;
      4290: inst = 32'h10408000;
      4291: inst = 32'hc404896;
      4292: inst = 32'h8220000;
      4293: inst = 32'h10408000;
      4294: inst = 32'hc404897;
      4295: inst = 32'h8220000;
      4296: inst = 32'h10408000;
      4297: inst = 32'hc404898;
      4298: inst = 32'h8220000;
      4299: inst = 32'h10408000;
      4300: inst = 32'hc404899;
      4301: inst = 32'h8220000;
      4302: inst = 32'h10408000;
      4303: inst = 32'hc40489a;
      4304: inst = 32'h8220000;
      4305: inst = 32'h10408000;
      4306: inst = 32'hc40489b;
      4307: inst = 32'h8220000;
      4308: inst = 32'h10408000;
      4309: inst = 32'hc4048c4;
      4310: inst = 32'h8220000;
      4311: inst = 32'h10408000;
      4312: inst = 32'hc4048c5;
      4313: inst = 32'h8220000;
      4314: inst = 32'h10408000;
      4315: inst = 32'hc4048c6;
      4316: inst = 32'h8220000;
      4317: inst = 32'h10408000;
      4318: inst = 32'hc4048c7;
      4319: inst = 32'h8220000;
      4320: inst = 32'h10408000;
      4321: inst = 32'hc4048c8;
      4322: inst = 32'h8220000;
      4323: inst = 32'h10408000;
      4324: inst = 32'hc4048c9;
      4325: inst = 32'h8220000;
      4326: inst = 32'h10408000;
      4327: inst = 32'hc4048ca;
      4328: inst = 32'h8220000;
      4329: inst = 32'h10408000;
      4330: inst = 32'hc4048cb;
      4331: inst = 32'h8220000;
      4332: inst = 32'h10408000;
      4333: inst = 32'hc4048cc;
      4334: inst = 32'h8220000;
      4335: inst = 32'h10408000;
      4336: inst = 32'hc4048cd;
      4337: inst = 32'h8220000;
      4338: inst = 32'h10408000;
      4339: inst = 32'hc4048ce;
      4340: inst = 32'h8220000;
      4341: inst = 32'h10408000;
      4342: inst = 32'hc4048e0;
      4343: inst = 32'h8220000;
      4344: inst = 32'h10408000;
      4345: inst = 32'hc4048e1;
      4346: inst = 32'h8220000;
      4347: inst = 32'h10408000;
      4348: inst = 32'hc4048e2;
      4349: inst = 32'h8220000;
      4350: inst = 32'h10408000;
      4351: inst = 32'hc4048e3;
      4352: inst = 32'h8220000;
      4353: inst = 32'h10408000;
      4354: inst = 32'hc4048e4;
      4355: inst = 32'h8220000;
      4356: inst = 32'h10408000;
      4357: inst = 32'hc4048e5;
      4358: inst = 32'h8220000;
      4359: inst = 32'h10408000;
      4360: inst = 32'hc4048e6;
      4361: inst = 32'h8220000;
      4362: inst = 32'h10408000;
      4363: inst = 32'hc4048e7;
      4364: inst = 32'h8220000;
      4365: inst = 32'h10408000;
      4366: inst = 32'hc4048e8;
      4367: inst = 32'h8220000;
      4368: inst = 32'h10408000;
      4369: inst = 32'hc4048e9;
      4370: inst = 32'h8220000;
      4371: inst = 32'h10408000;
      4372: inst = 32'hc4048ea;
      4373: inst = 32'h8220000;
      4374: inst = 32'h10408000;
      4375: inst = 32'hc4048eb;
      4376: inst = 32'h8220000;
      4377: inst = 32'h10408000;
      4378: inst = 32'hc4048ec;
      4379: inst = 32'h8220000;
      4380: inst = 32'h10408000;
      4381: inst = 32'hc4048ed;
      4382: inst = 32'h8220000;
      4383: inst = 32'h10408000;
      4384: inst = 32'hc4048ee;
      4385: inst = 32'h8220000;
      4386: inst = 32'h10408000;
      4387: inst = 32'hc4048ef;
      4388: inst = 32'h8220000;
      4389: inst = 32'h10408000;
      4390: inst = 32'hc4048f0;
      4391: inst = 32'h8220000;
      4392: inst = 32'h10408000;
      4393: inst = 32'hc4048f1;
      4394: inst = 32'h8220000;
      4395: inst = 32'h10408000;
      4396: inst = 32'hc4048f2;
      4397: inst = 32'h8220000;
      4398: inst = 32'h10408000;
      4399: inst = 32'hc4048f3;
      4400: inst = 32'h8220000;
      4401: inst = 32'h10408000;
      4402: inst = 32'hc4048f4;
      4403: inst = 32'h8220000;
      4404: inst = 32'h10408000;
      4405: inst = 32'hc4048f5;
      4406: inst = 32'h8220000;
      4407: inst = 32'h10408000;
      4408: inst = 32'hc4048f6;
      4409: inst = 32'h8220000;
      4410: inst = 32'h10408000;
      4411: inst = 32'hc4048f7;
      4412: inst = 32'h8220000;
      4413: inst = 32'h10408000;
      4414: inst = 32'hc4048f8;
      4415: inst = 32'h8220000;
      4416: inst = 32'h10408000;
      4417: inst = 32'hc4048f9;
      4418: inst = 32'h8220000;
      4419: inst = 32'h10408000;
      4420: inst = 32'hc4048fa;
      4421: inst = 32'h8220000;
      4422: inst = 32'h10408000;
      4423: inst = 32'hc4048fb;
      4424: inst = 32'h8220000;
      4425: inst = 32'h10408000;
      4426: inst = 32'hc404924;
      4427: inst = 32'h8220000;
      4428: inst = 32'h10408000;
      4429: inst = 32'hc404925;
      4430: inst = 32'h8220000;
      4431: inst = 32'h10408000;
      4432: inst = 32'hc404926;
      4433: inst = 32'h8220000;
      4434: inst = 32'h10408000;
      4435: inst = 32'hc404927;
      4436: inst = 32'h8220000;
      4437: inst = 32'h10408000;
      4438: inst = 32'hc404928;
      4439: inst = 32'h8220000;
      4440: inst = 32'h10408000;
      4441: inst = 32'hc404929;
      4442: inst = 32'h8220000;
      4443: inst = 32'h10408000;
      4444: inst = 32'hc40492a;
      4445: inst = 32'h8220000;
      4446: inst = 32'h10408000;
      4447: inst = 32'hc40492b;
      4448: inst = 32'h8220000;
      4449: inst = 32'h10408000;
      4450: inst = 32'hc40492c;
      4451: inst = 32'h8220000;
      4452: inst = 32'h10408000;
      4453: inst = 32'hc40492d;
      4454: inst = 32'h8220000;
      4455: inst = 32'h10408000;
      4456: inst = 32'hc40492e;
      4457: inst = 32'h8220000;
      4458: inst = 32'h10408000;
      4459: inst = 32'hc404940;
      4460: inst = 32'h8220000;
      4461: inst = 32'h10408000;
      4462: inst = 32'hc404941;
      4463: inst = 32'h8220000;
      4464: inst = 32'h10408000;
      4465: inst = 32'hc404942;
      4466: inst = 32'h8220000;
      4467: inst = 32'h10408000;
      4468: inst = 32'hc404943;
      4469: inst = 32'h8220000;
      4470: inst = 32'h10408000;
      4471: inst = 32'hc404944;
      4472: inst = 32'h8220000;
      4473: inst = 32'h10408000;
      4474: inst = 32'hc404945;
      4475: inst = 32'h8220000;
      4476: inst = 32'h10408000;
      4477: inst = 32'hc404946;
      4478: inst = 32'h8220000;
      4479: inst = 32'h10408000;
      4480: inst = 32'hc404947;
      4481: inst = 32'h8220000;
      4482: inst = 32'h10408000;
      4483: inst = 32'hc404948;
      4484: inst = 32'h8220000;
      4485: inst = 32'h10408000;
      4486: inst = 32'hc404949;
      4487: inst = 32'h8220000;
      4488: inst = 32'h10408000;
      4489: inst = 32'hc40494a;
      4490: inst = 32'h8220000;
      4491: inst = 32'h10408000;
      4492: inst = 32'hc40494b;
      4493: inst = 32'h8220000;
      4494: inst = 32'h10408000;
      4495: inst = 32'hc40494c;
      4496: inst = 32'h8220000;
      4497: inst = 32'h10408000;
      4498: inst = 32'hc40494d;
      4499: inst = 32'h8220000;
      4500: inst = 32'h10408000;
      4501: inst = 32'hc40494e;
      4502: inst = 32'h8220000;
      4503: inst = 32'h10408000;
      4504: inst = 32'hc40494f;
      4505: inst = 32'h8220000;
      4506: inst = 32'h10408000;
      4507: inst = 32'hc404950;
      4508: inst = 32'h8220000;
      4509: inst = 32'h10408000;
      4510: inst = 32'hc404951;
      4511: inst = 32'h8220000;
      4512: inst = 32'h10408000;
      4513: inst = 32'hc404952;
      4514: inst = 32'h8220000;
      4515: inst = 32'h10408000;
      4516: inst = 32'hc404953;
      4517: inst = 32'h8220000;
      4518: inst = 32'h10408000;
      4519: inst = 32'hc404954;
      4520: inst = 32'h8220000;
      4521: inst = 32'h10408000;
      4522: inst = 32'hc404955;
      4523: inst = 32'h8220000;
      4524: inst = 32'h10408000;
      4525: inst = 32'hc404956;
      4526: inst = 32'h8220000;
      4527: inst = 32'h10408000;
      4528: inst = 32'hc404957;
      4529: inst = 32'h8220000;
      4530: inst = 32'h10408000;
      4531: inst = 32'hc404958;
      4532: inst = 32'h8220000;
      4533: inst = 32'h10408000;
      4534: inst = 32'hc404959;
      4535: inst = 32'h8220000;
      4536: inst = 32'h10408000;
      4537: inst = 32'hc40495a;
      4538: inst = 32'h8220000;
      4539: inst = 32'h10408000;
      4540: inst = 32'hc40495b;
      4541: inst = 32'h8220000;
      4542: inst = 32'h10408000;
      4543: inst = 32'hc404984;
      4544: inst = 32'h8220000;
      4545: inst = 32'h10408000;
      4546: inst = 32'hc404985;
      4547: inst = 32'h8220000;
      4548: inst = 32'h10408000;
      4549: inst = 32'hc404986;
      4550: inst = 32'h8220000;
      4551: inst = 32'h10408000;
      4552: inst = 32'hc404987;
      4553: inst = 32'h8220000;
      4554: inst = 32'h10408000;
      4555: inst = 32'hc404988;
      4556: inst = 32'h8220000;
      4557: inst = 32'h10408000;
      4558: inst = 32'hc404989;
      4559: inst = 32'h8220000;
      4560: inst = 32'h10408000;
      4561: inst = 32'hc40498a;
      4562: inst = 32'h8220000;
      4563: inst = 32'h10408000;
      4564: inst = 32'hc40498b;
      4565: inst = 32'h8220000;
      4566: inst = 32'h10408000;
      4567: inst = 32'hc40498c;
      4568: inst = 32'h8220000;
      4569: inst = 32'h10408000;
      4570: inst = 32'hc40498d;
      4571: inst = 32'h8220000;
      4572: inst = 32'h10408000;
      4573: inst = 32'hc40498e;
      4574: inst = 32'h8220000;
      4575: inst = 32'h10408000;
      4576: inst = 32'hc4049a0;
      4577: inst = 32'h8220000;
      4578: inst = 32'h10408000;
      4579: inst = 32'hc4049a1;
      4580: inst = 32'h8220000;
      4581: inst = 32'h10408000;
      4582: inst = 32'hc4049a2;
      4583: inst = 32'h8220000;
      4584: inst = 32'h10408000;
      4585: inst = 32'hc4049a3;
      4586: inst = 32'h8220000;
      4587: inst = 32'h10408000;
      4588: inst = 32'hc4049a4;
      4589: inst = 32'h8220000;
      4590: inst = 32'h10408000;
      4591: inst = 32'hc4049a5;
      4592: inst = 32'h8220000;
      4593: inst = 32'h10408000;
      4594: inst = 32'hc4049a6;
      4595: inst = 32'h8220000;
      4596: inst = 32'h10408000;
      4597: inst = 32'hc4049a7;
      4598: inst = 32'h8220000;
      4599: inst = 32'h10408000;
      4600: inst = 32'hc4049a8;
      4601: inst = 32'h8220000;
      4602: inst = 32'h10408000;
      4603: inst = 32'hc4049a9;
      4604: inst = 32'h8220000;
      4605: inst = 32'h10408000;
      4606: inst = 32'hc4049aa;
      4607: inst = 32'h8220000;
      4608: inst = 32'h10408000;
      4609: inst = 32'hc4049ab;
      4610: inst = 32'h8220000;
      4611: inst = 32'h10408000;
      4612: inst = 32'hc4049ac;
      4613: inst = 32'h8220000;
      4614: inst = 32'h10408000;
      4615: inst = 32'hc4049ad;
      4616: inst = 32'h8220000;
      4617: inst = 32'h10408000;
      4618: inst = 32'hc4049ae;
      4619: inst = 32'h8220000;
      4620: inst = 32'h10408000;
      4621: inst = 32'hc4049af;
      4622: inst = 32'h8220000;
      4623: inst = 32'h10408000;
      4624: inst = 32'hc4049b0;
      4625: inst = 32'h8220000;
      4626: inst = 32'h10408000;
      4627: inst = 32'hc4049b1;
      4628: inst = 32'h8220000;
      4629: inst = 32'h10408000;
      4630: inst = 32'hc4049b2;
      4631: inst = 32'h8220000;
      4632: inst = 32'h10408000;
      4633: inst = 32'hc4049b3;
      4634: inst = 32'h8220000;
      4635: inst = 32'h10408000;
      4636: inst = 32'hc4049b4;
      4637: inst = 32'h8220000;
      4638: inst = 32'h10408000;
      4639: inst = 32'hc4049b5;
      4640: inst = 32'h8220000;
      4641: inst = 32'h10408000;
      4642: inst = 32'hc4049b6;
      4643: inst = 32'h8220000;
      4644: inst = 32'h10408000;
      4645: inst = 32'hc4049b7;
      4646: inst = 32'h8220000;
      4647: inst = 32'h10408000;
      4648: inst = 32'hc4049b8;
      4649: inst = 32'h8220000;
      4650: inst = 32'h10408000;
      4651: inst = 32'hc4049b9;
      4652: inst = 32'h8220000;
      4653: inst = 32'h10408000;
      4654: inst = 32'hc4049ba;
      4655: inst = 32'h8220000;
      4656: inst = 32'h10408000;
      4657: inst = 32'hc4049bb;
      4658: inst = 32'h8220000;
      4659: inst = 32'h10408000;
      4660: inst = 32'hc4049e4;
      4661: inst = 32'h8220000;
      4662: inst = 32'h10408000;
      4663: inst = 32'hc4049e5;
      4664: inst = 32'h8220000;
      4665: inst = 32'h10408000;
      4666: inst = 32'hc4049e6;
      4667: inst = 32'h8220000;
      4668: inst = 32'h10408000;
      4669: inst = 32'hc4049e7;
      4670: inst = 32'h8220000;
      4671: inst = 32'h10408000;
      4672: inst = 32'hc4049e8;
      4673: inst = 32'h8220000;
      4674: inst = 32'h10408000;
      4675: inst = 32'hc4049e9;
      4676: inst = 32'h8220000;
      4677: inst = 32'h10408000;
      4678: inst = 32'hc4049ea;
      4679: inst = 32'h8220000;
      4680: inst = 32'h10408000;
      4681: inst = 32'hc4049eb;
      4682: inst = 32'h8220000;
      4683: inst = 32'h10408000;
      4684: inst = 32'hc4049ec;
      4685: inst = 32'h8220000;
      4686: inst = 32'h10408000;
      4687: inst = 32'hc4049ed;
      4688: inst = 32'h8220000;
      4689: inst = 32'h10408000;
      4690: inst = 32'hc4049ee;
      4691: inst = 32'h8220000;
      4692: inst = 32'h10408000;
      4693: inst = 32'hc404a00;
      4694: inst = 32'h8220000;
      4695: inst = 32'h10408000;
      4696: inst = 32'hc404a01;
      4697: inst = 32'h8220000;
      4698: inst = 32'h10408000;
      4699: inst = 32'hc404a02;
      4700: inst = 32'h8220000;
      4701: inst = 32'h10408000;
      4702: inst = 32'hc404a03;
      4703: inst = 32'h8220000;
      4704: inst = 32'h10408000;
      4705: inst = 32'hc404a04;
      4706: inst = 32'h8220000;
      4707: inst = 32'h10408000;
      4708: inst = 32'hc404a05;
      4709: inst = 32'h8220000;
      4710: inst = 32'h10408000;
      4711: inst = 32'hc404a06;
      4712: inst = 32'h8220000;
      4713: inst = 32'h10408000;
      4714: inst = 32'hc404a07;
      4715: inst = 32'h8220000;
      4716: inst = 32'h10408000;
      4717: inst = 32'hc404a0f;
      4718: inst = 32'h8220000;
      4719: inst = 32'h10408000;
      4720: inst = 32'hc404a10;
      4721: inst = 32'h8220000;
      4722: inst = 32'h10408000;
      4723: inst = 32'hc404a11;
      4724: inst = 32'h8220000;
      4725: inst = 32'h10408000;
      4726: inst = 32'hc404a12;
      4727: inst = 32'h8220000;
      4728: inst = 32'h10408000;
      4729: inst = 32'hc404a13;
      4730: inst = 32'h8220000;
      4731: inst = 32'h10408000;
      4732: inst = 32'hc404a14;
      4733: inst = 32'h8220000;
      4734: inst = 32'h10408000;
      4735: inst = 32'hc404a15;
      4736: inst = 32'h8220000;
      4737: inst = 32'h10408000;
      4738: inst = 32'hc404a16;
      4739: inst = 32'h8220000;
      4740: inst = 32'h10408000;
      4741: inst = 32'hc404a17;
      4742: inst = 32'h8220000;
      4743: inst = 32'h10408000;
      4744: inst = 32'hc404a18;
      4745: inst = 32'h8220000;
      4746: inst = 32'h10408000;
      4747: inst = 32'hc404a19;
      4748: inst = 32'h8220000;
      4749: inst = 32'h10408000;
      4750: inst = 32'hc404a1a;
      4751: inst = 32'h8220000;
      4752: inst = 32'h10408000;
      4753: inst = 32'hc404a1b;
      4754: inst = 32'h8220000;
      4755: inst = 32'h10408000;
      4756: inst = 32'hc404a44;
      4757: inst = 32'h8220000;
      4758: inst = 32'h10408000;
      4759: inst = 32'hc404a45;
      4760: inst = 32'h8220000;
      4761: inst = 32'h10408000;
      4762: inst = 32'hc404a46;
      4763: inst = 32'h8220000;
      4764: inst = 32'h10408000;
      4765: inst = 32'hc404a47;
      4766: inst = 32'h8220000;
      4767: inst = 32'h10408000;
      4768: inst = 32'hc404a48;
      4769: inst = 32'h8220000;
      4770: inst = 32'h10408000;
      4771: inst = 32'hc404a49;
      4772: inst = 32'h8220000;
      4773: inst = 32'h10408000;
      4774: inst = 32'hc404a4a;
      4775: inst = 32'h8220000;
      4776: inst = 32'h10408000;
      4777: inst = 32'hc404a4b;
      4778: inst = 32'h8220000;
      4779: inst = 32'h10408000;
      4780: inst = 32'hc404a4c;
      4781: inst = 32'h8220000;
      4782: inst = 32'h10408000;
      4783: inst = 32'hc404a4d;
      4784: inst = 32'h8220000;
      4785: inst = 32'h10408000;
      4786: inst = 32'hc404a4e;
      4787: inst = 32'h8220000;
      4788: inst = 32'h10408000;
      4789: inst = 32'hc404a60;
      4790: inst = 32'h8220000;
      4791: inst = 32'h10408000;
      4792: inst = 32'hc404a61;
      4793: inst = 32'h8220000;
      4794: inst = 32'h10408000;
      4795: inst = 32'hc404a62;
      4796: inst = 32'h8220000;
      4797: inst = 32'h10408000;
      4798: inst = 32'hc404a63;
      4799: inst = 32'h8220000;
      4800: inst = 32'h10408000;
      4801: inst = 32'hc404a64;
      4802: inst = 32'h8220000;
      4803: inst = 32'h10408000;
      4804: inst = 32'hc404a65;
      4805: inst = 32'h8220000;
      4806: inst = 32'h10408000;
      4807: inst = 32'hc404a66;
      4808: inst = 32'h8220000;
      4809: inst = 32'h10408000;
      4810: inst = 32'hc404a70;
      4811: inst = 32'h8220000;
      4812: inst = 32'h10408000;
      4813: inst = 32'hc404a71;
      4814: inst = 32'h8220000;
      4815: inst = 32'h10408000;
      4816: inst = 32'hc404a72;
      4817: inst = 32'h8220000;
      4818: inst = 32'h10408000;
      4819: inst = 32'hc404a73;
      4820: inst = 32'h8220000;
      4821: inst = 32'h10408000;
      4822: inst = 32'hc404a74;
      4823: inst = 32'h8220000;
      4824: inst = 32'h10408000;
      4825: inst = 32'hc404a75;
      4826: inst = 32'h8220000;
      4827: inst = 32'h10408000;
      4828: inst = 32'hc404a76;
      4829: inst = 32'h8220000;
      4830: inst = 32'h10408000;
      4831: inst = 32'hc404a77;
      4832: inst = 32'h8220000;
      4833: inst = 32'h10408000;
      4834: inst = 32'hc404a78;
      4835: inst = 32'h8220000;
      4836: inst = 32'h10408000;
      4837: inst = 32'hc404a79;
      4838: inst = 32'h8220000;
      4839: inst = 32'h10408000;
      4840: inst = 32'hc404a7a;
      4841: inst = 32'h8220000;
      4842: inst = 32'h10408000;
      4843: inst = 32'hc404a7b;
      4844: inst = 32'h8220000;
      4845: inst = 32'h10408000;
      4846: inst = 32'hc404aa4;
      4847: inst = 32'h8220000;
      4848: inst = 32'h10408000;
      4849: inst = 32'hc404aa5;
      4850: inst = 32'h8220000;
      4851: inst = 32'h10408000;
      4852: inst = 32'hc404aa6;
      4853: inst = 32'h8220000;
      4854: inst = 32'h10408000;
      4855: inst = 32'hc404aa7;
      4856: inst = 32'h8220000;
      4857: inst = 32'h10408000;
      4858: inst = 32'hc404aa8;
      4859: inst = 32'h8220000;
      4860: inst = 32'h10408000;
      4861: inst = 32'hc404aa9;
      4862: inst = 32'h8220000;
      4863: inst = 32'h10408000;
      4864: inst = 32'hc404aaa;
      4865: inst = 32'h8220000;
      4866: inst = 32'h10408000;
      4867: inst = 32'hc404aab;
      4868: inst = 32'h8220000;
      4869: inst = 32'h10408000;
      4870: inst = 32'hc404aac;
      4871: inst = 32'h8220000;
      4872: inst = 32'h10408000;
      4873: inst = 32'hc404aad;
      4874: inst = 32'h8220000;
      4875: inst = 32'h10408000;
      4876: inst = 32'hc404aae;
      4877: inst = 32'h8220000;
      4878: inst = 32'h10408000;
      4879: inst = 32'hc404ac0;
      4880: inst = 32'h8220000;
      4881: inst = 32'h10408000;
      4882: inst = 32'hc404ac1;
      4883: inst = 32'h8220000;
      4884: inst = 32'h10408000;
      4885: inst = 32'hc404ac2;
      4886: inst = 32'h8220000;
      4887: inst = 32'h10408000;
      4888: inst = 32'hc404ac3;
      4889: inst = 32'h8220000;
      4890: inst = 32'h10408000;
      4891: inst = 32'hc404ac4;
      4892: inst = 32'h8220000;
      4893: inst = 32'h10408000;
      4894: inst = 32'hc404ac5;
      4895: inst = 32'h8220000;
      4896: inst = 32'h10408000;
      4897: inst = 32'hc404ac6;
      4898: inst = 32'h8220000;
      4899: inst = 32'h10408000;
      4900: inst = 32'hc404ad0;
      4901: inst = 32'h8220000;
      4902: inst = 32'h10408000;
      4903: inst = 32'hc404ad1;
      4904: inst = 32'h8220000;
      4905: inst = 32'h10408000;
      4906: inst = 32'hc404ad2;
      4907: inst = 32'h8220000;
      4908: inst = 32'h10408000;
      4909: inst = 32'hc404ad3;
      4910: inst = 32'h8220000;
      4911: inst = 32'h10408000;
      4912: inst = 32'hc404ad4;
      4913: inst = 32'h8220000;
      4914: inst = 32'h10408000;
      4915: inst = 32'hc404ad5;
      4916: inst = 32'h8220000;
      4917: inst = 32'h10408000;
      4918: inst = 32'hc404ad6;
      4919: inst = 32'h8220000;
      4920: inst = 32'h10408000;
      4921: inst = 32'hc404ad7;
      4922: inst = 32'h8220000;
      4923: inst = 32'h10408000;
      4924: inst = 32'hc404ad8;
      4925: inst = 32'h8220000;
      4926: inst = 32'h10408000;
      4927: inst = 32'hc404ad9;
      4928: inst = 32'h8220000;
      4929: inst = 32'h10408000;
      4930: inst = 32'hc404ada;
      4931: inst = 32'h8220000;
      4932: inst = 32'h10408000;
      4933: inst = 32'hc404adb;
      4934: inst = 32'h8220000;
      4935: inst = 32'h10408000;
      4936: inst = 32'hc404b04;
      4937: inst = 32'h8220000;
      4938: inst = 32'h10408000;
      4939: inst = 32'hc404b05;
      4940: inst = 32'h8220000;
      4941: inst = 32'h10408000;
      4942: inst = 32'hc404b06;
      4943: inst = 32'h8220000;
      4944: inst = 32'h10408000;
      4945: inst = 32'hc404b07;
      4946: inst = 32'h8220000;
      4947: inst = 32'h10408000;
      4948: inst = 32'hc404b08;
      4949: inst = 32'h8220000;
      4950: inst = 32'h10408000;
      4951: inst = 32'hc404b09;
      4952: inst = 32'h8220000;
      4953: inst = 32'h10408000;
      4954: inst = 32'hc404b0a;
      4955: inst = 32'h8220000;
      4956: inst = 32'h10408000;
      4957: inst = 32'hc404b0b;
      4958: inst = 32'h8220000;
      4959: inst = 32'h10408000;
      4960: inst = 32'hc404b0c;
      4961: inst = 32'h8220000;
      4962: inst = 32'h10408000;
      4963: inst = 32'hc404b0d;
      4964: inst = 32'h8220000;
      4965: inst = 32'h10408000;
      4966: inst = 32'hc404b0e;
      4967: inst = 32'h8220000;
      4968: inst = 32'h10408000;
      4969: inst = 32'hc404b20;
      4970: inst = 32'h8220000;
      4971: inst = 32'h10408000;
      4972: inst = 32'hc404b21;
      4973: inst = 32'h8220000;
      4974: inst = 32'h10408000;
      4975: inst = 32'hc404b22;
      4976: inst = 32'h8220000;
      4977: inst = 32'h10408000;
      4978: inst = 32'hc404b23;
      4979: inst = 32'h8220000;
      4980: inst = 32'h10408000;
      4981: inst = 32'hc404b24;
      4982: inst = 32'h8220000;
      4983: inst = 32'h10408000;
      4984: inst = 32'hc404b25;
      4985: inst = 32'h8220000;
      4986: inst = 32'h10408000;
      4987: inst = 32'hc404b26;
      4988: inst = 32'h8220000;
      4989: inst = 32'h10408000;
      4990: inst = 32'hc404b30;
      4991: inst = 32'h8220000;
      4992: inst = 32'h10408000;
      4993: inst = 32'hc404b31;
      4994: inst = 32'h8220000;
      4995: inst = 32'h10408000;
      4996: inst = 32'hc404b32;
      4997: inst = 32'h8220000;
      4998: inst = 32'h10408000;
      4999: inst = 32'hc404b33;
      5000: inst = 32'h8220000;
      5001: inst = 32'h10408000;
      5002: inst = 32'hc404b34;
      5003: inst = 32'h8220000;
      5004: inst = 32'h10408000;
      5005: inst = 32'hc404b35;
      5006: inst = 32'h8220000;
      5007: inst = 32'h10408000;
      5008: inst = 32'hc404b36;
      5009: inst = 32'h8220000;
      5010: inst = 32'h10408000;
      5011: inst = 32'hc404b37;
      5012: inst = 32'h8220000;
      5013: inst = 32'h10408000;
      5014: inst = 32'hc404b38;
      5015: inst = 32'h8220000;
      5016: inst = 32'h10408000;
      5017: inst = 32'hc404b39;
      5018: inst = 32'h8220000;
      5019: inst = 32'h10408000;
      5020: inst = 32'hc404b3a;
      5021: inst = 32'h8220000;
      5022: inst = 32'h10408000;
      5023: inst = 32'hc404b3b;
      5024: inst = 32'h8220000;
      5025: inst = 32'h10408000;
      5026: inst = 32'hc404b64;
      5027: inst = 32'h8220000;
      5028: inst = 32'h10408000;
      5029: inst = 32'hc404b65;
      5030: inst = 32'h8220000;
      5031: inst = 32'h10408000;
      5032: inst = 32'hc404b66;
      5033: inst = 32'h8220000;
      5034: inst = 32'h10408000;
      5035: inst = 32'hc404b67;
      5036: inst = 32'h8220000;
      5037: inst = 32'h10408000;
      5038: inst = 32'hc404b68;
      5039: inst = 32'h8220000;
      5040: inst = 32'h10408000;
      5041: inst = 32'hc404b69;
      5042: inst = 32'h8220000;
      5043: inst = 32'h10408000;
      5044: inst = 32'hc404b6a;
      5045: inst = 32'h8220000;
      5046: inst = 32'h10408000;
      5047: inst = 32'hc404b6b;
      5048: inst = 32'h8220000;
      5049: inst = 32'h10408000;
      5050: inst = 32'hc404b6c;
      5051: inst = 32'h8220000;
      5052: inst = 32'h10408000;
      5053: inst = 32'hc404b6d;
      5054: inst = 32'h8220000;
      5055: inst = 32'h10408000;
      5056: inst = 32'hc404b6e;
      5057: inst = 32'h8220000;
      5058: inst = 32'h10408000;
      5059: inst = 32'hc404b80;
      5060: inst = 32'h8220000;
      5061: inst = 32'h10408000;
      5062: inst = 32'hc404b81;
      5063: inst = 32'h8220000;
      5064: inst = 32'h10408000;
      5065: inst = 32'hc404b82;
      5066: inst = 32'h8220000;
      5067: inst = 32'h10408000;
      5068: inst = 32'hc404b83;
      5069: inst = 32'h8220000;
      5070: inst = 32'h10408000;
      5071: inst = 32'hc404b84;
      5072: inst = 32'h8220000;
      5073: inst = 32'h10408000;
      5074: inst = 32'hc404b85;
      5075: inst = 32'h8220000;
      5076: inst = 32'h10408000;
      5077: inst = 32'hc404b86;
      5078: inst = 32'h8220000;
      5079: inst = 32'h10408000;
      5080: inst = 32'hc404b90;
      5081: inst = 32'h8220000;
      5082: inst = 32'h10408000;
      5083: inst = 32'hc404b91;
      5084: inst = 32'h8220000;
      5085: inst = 32'h10408000;
      5086: inst = 32'hc404b92;
      5087: inst = 32'h8220000;
      5088: inst = 32'h10408000;
      5089: inst = 32'hc404b93;
      5090: inst = 32'h8220000;
      5091: inst = 32'h10408000;
      5092: inst = 32'hc404b94;
      5093: inst = 32'h8220000;
      5094: inst = 32'h10408000;
      5095: inst = 32'hc404b95;
      5096: inst = 32'h8220000;
      5097: inst = 32'h10408000;
      5098: inst = 32'hc404b96;
      5099: inst = 32'h8220000;
      5100: inst = 32'h10408000;
      5101: inst = 32'hc404b97;
      5102: inst = 32'h8220000;
      5103: inst = 32'h10408000;
      5104: inst = 32'hc404b98;
      5105: inst = 32'h8220000;
      5106: inst = 32'h10408000;
      5107: inst = 32'hc404b99;
      5108: inst = 32'h8220000;
      5109: inst = 32'h10408000;
      5110: inst = 32'hc404b9a;
      5111: inst = 32'h8220000;
      5112: inst = 32'h10408000;
      5113: inst = 32'hc404b9b;
      5114: inst = 32'h8220000;
      5115: inst = 32'h10408000;
      5116: inst = 32'hc404bc4;
      5117: inst = 32'h8220000;
      5118: inst = 32'h10408000;
      5119: inst = 32'hc404bc5;
      5120: inst = 32'h8220000;
      5121: inst = 32'h10408000;
      5122: inst = 32'hc404bc6;
      5123: inst = 32'h8220000;
      5124: inst = 32'h10408000;
      5125: inst = 32'hc404bc7;
      5126: inst = 32'h8220000;
      5127: inst = 32'h10408000;
      5128: inst = 32'hc404bc8;
      5129: inst = 32'h8220000;
      5130: inst = 32'h10408000;
      5131: inst = 32'hc404bc9;
      5132: inst = 32'h8220000;
      5133: inst = 32'h10408000;
      5134: inst = 32'hc404bca;
      5135: inst = 32'h8220000;
      5136: inst = 32'h10408000;
      5137: inst = 32'hc404bcb;
      5138: inst = 32'h8220000;
      5139: inst = 32'h10408000;
      5140: inst = 32'hc404bcc;
      5141: inst = 32'h8220000;
      5142: inst = 32'h10408000;
      5143: inst = 32'hc404bcd;
      5144: inst = 32'h8220000;
      5145: inst = 32'h10408000;
      5146: inst = 32'hc404bce;
      5147: inst = 32'h8220000;
      5148: inst = 32'h10408000;
      5149: inst = 32'hc404be0;
      5150: inst = 32'h8220000;
      5151: inst = 32'h10408000;
      5152: inst = 32'hc404be1;
      5153: inst = 32'h8220000;
      5154: inst = 32'h10408000;
      5155: inst = 32'hc404be2;
      5156: inst = 32'h8220000;
      5157: inst = 32'h10408000;
      5158: inst = 32'hc404be3;
      5159: inst = 32'h8220000;
      5160: inst = 32'h10408000;
      5161: inst = 32'hc404be4;
      5162: inst = 32'h8220000;
      5163: inst = 32'h10408000;
      5164: inst = 32'hc404be5;
      5165: inst = 32'h8220000;
      5166: inst = 32'h10408000;
      5167: inst = 32'hc404be6;
      5168: inst = 32'h8220000;
      5169: inst = 32'h10408000;
      5170: inst = 32'hc404bf0;
      5171: inst = 32'h8220000;
      5172: inst = 32'h10408000;
      5173: inst = 32'hc404bf1;
      5174: inst = 32'h8220000;
      5175: inst = 32'h10408000;
      5176: inst = 32'hc404bf2;
      5177: inst = 32'h8220000;
      5178: inst = 32'h10408000;
      5179: inst = 32'hc404bf3;
      5180: inst = 32'h8220000;
      5181: inst = 32'h10408000;
      5182: inst = 32'hc404bf4;
      5183: inst = 32'h8220000;
      5184: inst = 32'h10408000;
      5185: inst = 32'hc404bf5;
      5186: inst = 32'h8220000;
      5187: inst = 32'h10408000;
      5188: inst = 32'hc404bf6;
      5189: inst = 32'h8220000;
      5190: inst = 32'h10408000;
      5191: inst = 32'hc404bf7;
      5192: inst = 32'h8220000;
      5193: inst = 32'h10408000;
      5194: inst = 32'hc404bf8;
      5195: inst = 32'h8220000;
      5196: inst = 32'h10408000;
      5197: inst = 32'hc404bf9;
      5198: inst = 32'h8220000;
      5199: inst = 32'h10408000;
      5200: inst = 32'hc404c26;
      5201: inst = 32'h8220000;
      5202: inst = 32'h10408000;
      5203: inst = 32'hc404c27;
      5204: inst = 32'h8220000;
      5205: inst = 32'h10408000;
      5206: inst = 32'hc404c28;
      5207: inst = 32'h8220000;
      5208: inst = 32'h10408000;
      5209: inst = 32'hc404c29;
      5210: inst = 32'h8220000;
      5211: inst = 32'h10408000;
      5212: inst = 32'hc404c2a;
      5213: inst = 32'h8220000;
      5214: inst = 32'h10408000;
      5215: inst = 32'hc404c2b;
      5216: inst = 32'h8220000;
      5217: inst = 32'h10408000;
      5218: inst = 32'hc404c2c;
      5219: inst = 32'h8220000;
      5220: inst = 32'h10408000;
      5221: inst = 32'hc404c2d;
      5222: inst = 32'h8220000;
      5223: inst = 32'h10408000;
      5224: inst = 32'hc404c2e;
      5225: inst = 32'h8220000;
      5226: inst = 32'h10408000;
      5227: inst = 32'hc404c40;
      5228: inst = 32'h8220000;
      5229: inst = 32'h10408000;
      5230: inst = 32'hc404c41;
      5231: inst = 32'h8220000;
      5232: inst = 32'h10408000;
      5233: inst = 32'hc404c42;
      5234: inst = 32'h8220000;
      5235: inst = 32'h10408000;
      5236: inst = 32'hc404c43;
      5237: inst = 32'h8220000;
      5238: inst = 32'h10408000;
      5239: inst = 32'hc404c44;
      5240: inst = 32'h8220000;
      5241: inst = 32'h10408000;
      5242: inst = 32'hc404c45;
      5243: inst = 32'h8220000;
      5244: inst = 32'h10408000;
      5245: inst = 32'hc404c46;
      5246: inst = 32'h8220000;
      5247: inst = 32'h10408000;
      5248: inst = 32'hc404c4f;
      5249: inst = 32'h8220000;
      5250: inst = 32'h10408000;
      5251: inst = 32'hc404c50;
      5252: inst = 32'h8220000;
      5253: inst = 32'h10408000;
      5254: inst = 32'hc404c51;
      5255: inst = 32'h8220000;
      5256: inst = 32'h10408000;
      5257: inst = 32'hc404c52;
      5258: inst = 32'h8220000;
      5259: inst = 32'h10408000;
      5260: inst = 32'hc404c53;
      5261: inst = 32'h8220000;
      5262: inst = 32'h10408000;
      5263: inst = 32'hc404c54;
      5264: inst = 32'h8220000;
      5265: inst = 32'h10408000;
      5266: inst = 32'hc404c55;
      5267: inst = 32'h8220000;
      5268: inst = 32'h10408000;
      5269: inst = 32'hc404c56;
      5270: inst = 32'h8220000;
      5271: inst = 32'h10408000;
      5272: inst = 32'hc404c57;
      5273: inst = 32'h8220000;
      5274: inst = 32'h10408000;
      5275: inst = 32'hc404c58;
      5276: inst = 32'h8220000;
      5277: inst = 32'h10408000;
      5278: inst = 32'hc404c59;
      5279: inst = 32'h8220000;
      5280: inst = 32'h10408000;
      5281: inst = 32'hc404c5a;
      5282: inst = 32'h8220000;
      5283: inst = 32'h10408000;
      5284: inst = 32'hc404c5b;
      5285: inst = 32'h8220000;
      5286: inst = 32'h10408000;
      5287: inst = 32'hc404c5c;
      5288: inst = 32'h8220000;
      5289: inst = 32'h10408000;
      5290: inst = 32'hc404c5d;
      5291: inst = 32'h8220000;
      5292: inst = 32'h10408000;
      5293: inst = 32'hc404c5e;
      5294: inst = 32'h8220000;
      5295: inst = 32'h10408000;
      5296: inst = 32'hc404c5f;
      5297: inst = 32'h8220000;
      5298: inst = 32'h10408000;
      5299: inst = 32'hc404c60;
      5300: inst = 32'h8220000;
      5301: inst = 32'h10408000;
      5302: inst = 32'hc404c61;
      5303: inst = 32'h8220000;
      5304: inst = 32'h10408000;
      5305: inst = 32'hc404c62;
      5306: inst = 32'h8220000;
      5307: inst = 32'h10408000;
      5308: inst = 32'hc404c63;
      5309: inst = 32'h8220000;
      5310: inst = 32'h10408000;
      5311: inst = 32'hc404c64;
      5312: inst = 32'h8220000;
      5313: inst = 32'h10408000;
      5314: inst = 32'hc404c65;
      5315: inst = 32'h8220000;
      5316: inst = 32'h10408000;
      5317: inst = 32'hc404c66;
      5318: inst = 32'h8220000;
      5319: inst = 32'h10408000;
      5320: inst = 32'hc404c67;
      5321: inst = 32'h8220000;
      5322: inst = 32'h10408000;
      5323: inst = 32'hc404c68;
      5324: inst = 32'h8220000;
      5325: inst = 32'h10408000;
      5326: inst = 32'hc404c69;
      5327: inst = 32'h8220000;
      5328: inst = 32'h10408000;
      5329: inst = 32'hc404c6a;
      5330: inst = 32'h8220000;
      5331: inst = 32'h10408000;
      5332: inst = 32'hc404c6b;
      5333: inst = 32'h8220000;
      5334: inst = 32'h10408000;
      5335: inst = 32'hc404c6c;
      5336: inst = 32'h8220000;
      5337: inst = 32'h10408000;
      5338: inst = 32'hc404c6d;
      5339: inst = 32'h8220000;
      5340: inst = 32'h10408000;
      5341: inst = 32'hc404c6e;
      5342: inst = 32'h8220000;
      5343: inst = 32'h10408000;
      5344: inst = 32'hc404c6f;
      5345: inst = 32'h8220000;
      5346: inst = 32'h10408000;
      5347: inst = 32'hc404c70;
      5348: inst = 32'h8220000;
      5349: inst = 32'h10408000;
      5350: inst = 32'hc404c71;
      5351: inst = 32'h8220000;
      5352: inst = 32'h10408000;
      5353: inst = 32'hc404c72;
      5354: inst = 32'h8220000;
      5355: inst = 32'h10408000;
      5356: inst = 32'hc404c73;
      5357: inst = 32'h8220000;
      5358: inst = 32'h10408000;
      5359: inst = 32'hc404c74;
      5360: inst = 32'h8220000;
      5361: inst = 32'h10408000;
      5362: inst = 32'hc404c75;
      5363: inst = 32'h8220000;
      5364: inst = 32'h10408000;
      5365: inst = 32'hc404c76;
      5366: inst = 32'h8220000;
      5367: inst = 32'h10408000;
      5368: inst = 32'hc404c77;
      5369: inst = 32'h8220000;
      5370: inst = 32'h10408000;
      5371: inst = 32'hc404c78;
      5372: inst = 32'h8220000;
      5373: inst = 32'h10408000;
      5374: inst = 32'hc404c79;
      5375: inst = 32'h8220000;
      5376: inst = 32'h10408000;
      5377: inst = 32'hc404c7a;
      5378: inst = 32'h8220000;
      5379: inst = 32'h10408000;
      5380: inst = 32'hc404c7b;
      5381: inst = 32'h8220000;
      5382: inst = 32'h10408000;
      5383: inst = 32'hc404c7c;
      5384: inst = 32'h8220000;
      5385: inst = 32'h10408000;
      5386: inst = 32'hc404c7d;
      5387: inst = 32'h8220000;
      5388: inst = 32'h10408000;
      5389: inst = 32'hc404c7e;
      5390: inst = 32'h8220000;
      5391: inst = 32'h10408000;
      5392: inst = 32'hc404c7f;
      5393: inst = 32'h8220000;
      5394: inst = 32'h10408000;
      5395: inst = 32'hc404c80;
      5396: inst = 32'h8220000;
      5397: inst = 32'h10408000;
      5398: inst = 32'hc404c81;
      5399: inst = 32'h8220000;
      5400: inst = 32'h10408000;
      5401: inst = 32'hc404c82;
      5402: inst = 32'h8220000;
      5403: inst = 32'h10408000;
      5404: inst = 32'hc404c83;
      5405: inst = 32'h8220000;
      5406: inst = 32'h10408000;
      5407: inst = 32'hc404c84;
      5408: inst = 32'h8220000;
      5409: inst = 32'h10408000;
      5410: inst = 32'hc404c85;
      5411: inst = 32'h8220000;
      5412: inst = 32'h10408000;
      5413: inst = 32'hc404c86;
      5414: inst = 32'h8220000;
      5415: inst = 32'h10408000;
      5416: inst = 32'hc404c87;
      5417: inst = 32'h8220000;
      5418: inst = 32'h10408000;
      5419: inst = 32'hc404c88;
      5420: inst = 32'h8220000;
      5421: inst = 32'h10408000;
      5422: inst = 32'hc404c89;
      5423: inst = 32'h8220000;
      5424: inst = 32'h10408000;
      5425: inst = 32'hc404c8a;
      5426: inst = 32'h8220000;
      5427: inst = 32'h10408000;
      5428: inst = 32'hc404c8b;
      5429: inst = 32'h8220000;
      5430: inst = 32'h10408000;
      5431: inst = 32'hc404c8c;
      5432: inst = 32'h8220000;
      5433: inst = 32'h10408000;
      5434: inst = 32'hc404c8d;
      5435: inst = 32'h8220000;
      5436: inst = 32'h10408000;
      5437: inst = 32'hc404c8e;
      5438: inst = 32'h8220000;
      5439: inst = 32'h10408000;
      5440: inst = 32'hc404ca0;
      5441: inst = 32'h8220000;
      5442: inst = 32'h10408000;
      5443: inst = 32'hc404ca1;
      5444: inst = 32'h8220000;
      5445: inst = 32'h10408000;
      5446: inst = 32'hc404cb7;
      5447: inst = 32'h8220000;
      5448: inst = 32'h10408000;
      5449: inst = 32'hc404cb8;
      5450: inst = 32'h8220000;
      5451: inst = 32'h10408000;
      5452: inst = 32'hc404cb9;
      5453: inst = 32'h8220000;
      5454: inst = 32'h10408000;
      5455: inst = 32'hc404cba;
      5456: inst = 32'h8220000;
      5457: inst = 32'h10408000;
      5458: inst = 32'hc404cbb;
      5459: inst = 32'h8220000;
      5460: inst = 32'h10408000;
      5461: inst = 32'hc404cbc;
      5462: inst = 32'h8220000;
      5463: inst = 32'h10408000;
      5464: inst = 32'hc404cbd;
      5465: inst = 32'h8220000;
      5466: inst = 32'h10408000;
      5467: inst = 32'hc404cbe;
      5468: inst = 32'h8220000;
      5469: inst = 32'h10408000;
      5470: inst = 32'hc404cbf;
      5471: inst = 32'h8220000;
      5472: inst = 32'h10408000;
      5473: inst = 32'hc404cc0;
      5474: inst = 32'h8220000;
      5475: inst = 32'h10408000;
      5476: inst = 32'hc404cc1;
      5477: inst = 32'h8220000;
      5478: inst = 32'h10408000;
      5479: inst = 32'hc404cc2;
      5480: inst = 32'h8220000;
      5481: inst = 32'h10408000;
      5482: inst = 32'hc404cc3;
      5483: inst = 32'h8220000;
      5484: inst = 32'h10408000;
      5485: inst = 32'hc404cc4;
      5486: inst = 32'h8220000;
      5487: inst = 32'h10408000;
      5488: inst = 32'hc404cc5;
      5489: inst = 32'h8220000;
      5490: inst = 32'h10408000;
      5491: inst = 32'hc404cc6;
      5492: inst = 32'h8220000;
      5493: inst = 32'h10408000;
      5494: inst = 32'hc404cc7;
      5495: inst = 32'h8220000;
      5496: inst = 32'h10408000;
      5497: inst = 32'hc404cc8;
      5498: inst = 32'h8220000;
      5499: inst = 32'h10408000;
      5500: inst = 32'hc404cc9;
      5501: inst = 32'h8220000;
      5502: inst = 32'h10408000;
      5503: inst = 32'hc404cca;
      5504: inst = 32'h8220000;
      5505: inst = 32'h10408000;
      5506: inst = 32'hc404ccb;
      5507: inst = 32'h8220000;
      5508: inst = 32'h10408000;
      5509: inst = 32'hc404ccc;
      5510: inst = 32'h8220000;
      5511: inst = 32'h10408000;
      5512: inst = 32'hc404ccd;
      5513: inst = 32'h8220000;
      5514: inst = 32'h10408000;
      5515: inst = 32'hc404cce;
      5516: inst = 32'h8220000;
      5517: inst = 32'h10408000;
      5518: inst = 32'hc404ccf;
      5519: inst = 32'h8220000;
      5520: inst = 32'h10408000;
      5521: inst = 32'hc404cd0;
      5522: inst = 32'h8220000;
      5523: inst = 32'h10408000;
      5524: inst = 32'hc404cd1;
      5525: inst = 32'h8220000;
      5526: inst = 32'h10408000;
      5527: inst = 32'hc404cd2;
      5528: inst = 32'h8220000;
      5529: inst = 32'h10408000;
      5530: inst = 32'hc404cd3;
      5531: inst = 32'h8220000;
      5532: inst = 32'h10408000;
      5533: inst = 32'hc404cd4;
      5534: inst = 32'h8220000;
      5535: inst = 32'h10408000;
      5536: inst = 32'hc404cd5;
      5537: inst = 32'h8220000;
      5538: inst = 32'h10408000;
      5539: inst = 32'hc404cd6;
      5540: inst = 32'h8220000;
      5541: inst = 32'h10408000;
      5542: inst = 32'hc404cd7;
      5543: inst = 32'h8220000;
      5544: inst = 32'h10408000;
      5545: inst = 32'hc404cd8;
      5546: inst = 32'h8220000;
      5547: inst = 32'h10408000;
      5548: inst = 32'hc404cd9;
      5549: inst = 32'h8220000;
      5550: inst = 32'h10408000;
      5551: inst = 32'hc404cda;
      5552: inst = 32'h8220000;
      5553: inst = 32'h10408000;
      5554: inst = 32'hc404cdb;
      5555: inst = 32'h8220000;
      5556: inst = 32'h10408000;
      5557: inst = 32'hc404cdc;
      5558: inst = 32'h8220000;
      5559: inst = 32'h10408000;
      5560: inst = 32'hc404cdd;
      5561: inst = 32'h8220000;
      5562: inst = 32'h10408000;
      5563: inst = 32'hc404cde;
      5564: inst = 32'h8220000;
      5565: inst = 32'h10408000;
      5566: inst = 32'hc404cdf;
      5567: inst = 32'h8220000;
      5568: inst = 32'h10408000;
      5569: inst = 32'hc404ce0;
      5570: inst = 32'h8220000;
      5571: inst = 32'h10408000;
      5572: inst = 32'hc404ce1;
      5573: inst = 32'h8220000;
      5574: inst = 32'h10408000;
      5575: inst = 32'hc404ce2;
      5576: inst = 32'h8220000;
      5577: inst = 32'h10408000;
      5578: inst = 32'hc404ce3;
      5579: inst = 32'h8220000;
      5580: inst = 32'h10408000;
      5581: inst = 32'hc404ce4;
      5582: inst = 32'h8220000;
      5583: inst = 32'h10408000;
      5584: inst = 32'hc404ce5;
      5585: inst = 32'h8220000;
      5586: inst = 32'h10408000;
      5587: inst = 32'hc404ce6;
      5588: inst = 32'h8220000;
      5589: inst = 32'h10408000;
      5590: inst = 32'hc404ce7;
      5591: inst = 32'h8220000;
      5592: inst = 32'h10408000;
      5593: inst = 32'hc404ce8;
      5594: inst = 32'h8220000;
      5595: inst = 32'h10408000;
      5596: inst = 32'hc404ce9;
      5597: inst = 32'h8220000;
      5598: inst = 32'h10408000;
      5599: inst = 32'hc404cea;
      5600: inst = 32'h8220000;
      5601: inst = 32'h10408000;
      5602: inst = 32'hc404ceb;
      5603: inst = 32'h8220000;
      5604: inst = 32'h10408000;
      5605: inst = 32'hc404cec;
      5606: inst = 32'h8220000;
      5607: inst = 32'h10408000;
      5608: inst = 32'hc404ced;
      5609: inst = 32'h8220000;
      5610: inst = 32'h10408000;
      5611: inst = 32'hc404cee;
      5612: inst = 32'h8220000;
      5613: inst = 32'h10408000;
      5614: inst = 32'hc404d17;
      5615: inst = 32'h8220000;
      5616: inst = 32'h10408000;
      5617: inst = 32'hc404d18;
      5618: inst = 32'h8220000;
      5619: inst = 32'h10408000;
      5620: inst = 32'hc404d19;
      5621: inst = 32'h8220000;
      5622: inst = 32'h10408000;
      5623: inst = 32'hc404d1a;
      5624: inst = 32'h8220000;
      5625: inst = 32'h10408000;
      5626: inst = 32'hc404d1b;
      5627: inst = 32'h8220000;
      5628: inst = 32'h10408000;
      5629: inst = 32'hc404d1c;
      5630: inst = 32'h8220000;
      5631: inst = 32'h10408000;
      5632: inst = 32'hc404d1d;
      5633: inst = 32'h8220000;
      5634: inst = 32'h10408000;
      5635: inst = 32'hc404d1e;
      5636: inst = 32'h8220000;
      5637: inst = 32'h10408000;
      5638: inst = 32'hc404d1f;
      5639: inst = 32'h8220000;
      5640: inst = 32'h10408000;
      5641: inst = 32'hc404d20;
      5642: inst = 32'h8220000;
      5643: inst = 32'h10408000;
      5644: inst = 32'hc404d21;
      5645: inst = 32'h8220000;
      5646: inst = 32'h10408000;
      5647: inst = 32'hc404d22;
      5648: inst = 32'h8220000;
      5649: inst = 32'h10408000;
      5650: inst = 32'hc404d23;
      5651: inst = 32'h8220000;
      5652: inst = 32'h10408000;
      5653: inst = 32'hc404d24;
      5654: inst = 32'h8220000;
      5655: inst = 32'h10408000;
      5656: inst = 32'hc404d25;
      5657: inst = 32'h8220000;
      5658: inst = 32'h10408000;
      5659: inst = 32'hc404d26;
      5660: inst = 32'h8220000;
      5661: inst = 32'h10408000;
      5662: inst = 32'hc404d27;
      5663: inst = 32'h8220000;
      5664: inst = 32'h10408000;
      5665: inst = 32'hc404d28;
      5666: inst = 32'h8220000;
      5667: inst = 32'h10408000;
      5668: inst = 32'hc404d29;
      5669: inst = 32'h8220000;
      5670: inst = 32'h10408000;
      5671: inst = 32'hc404d2a;
      5672: inst = 32'h8220000;
      5673: inst = 32'h10408000;
      5674: inst = 32'hc404d2b;
      5675: inst = 32'h8220000;
      5676: inst = 32'h10408000;
      5677: inst = 32'hc404d2c;
      5678: inst = 32'h8220000;
      5679: inst = 32'h10408000;
      5680: inst = 32'hc404d2d;
      5681: inst = 32'h8220000;
      5682: inst = 32'h10408000;
      5683: inst = 32'hc404d2e;
      5684: inst = 32'h8220000;
      5685: inst = 32'h10408000;
      5686: inst = 32'hc404d2f;
      5687: inst = 32'h8220000;
      5688: inst = 32'h10408000;
      5689: inst = 32'hc404d30;
      5690: inst = 32'h8220000;
      5691: inst = 32'h10408000;
      5692: inst = 32'hc404d31;
      5693: inst = 32'h8220000;
      5694: inst = 32'h10408000;
      5695: inst = 32'hc404d32;
      5696: inst = 32'h8220000;
      5697: inst = 32'h10408000;
      5698: inst = 32'hc404d33;
      5699: inst = 32'h8220000;
      5700: inst = 32'h10408000;
      5701: inst = 32'hc404d34;
      5702: inst = 32'h8220000;
      5703: inst = 32'h10408000;
      5704: inst = 32'hc404d35;
      5705: inst = 32'h8220000;
      5706: inst = 32'h10408000;
      5707: inst = 32'hc404d36;
      5708: inst = 32'h8220000;
      5709: inst = 32'h10408000;
      5710: inst = 32'hc404d37;
      5711: inst = 32'h8220000;
      5712: inst = 32'h10408000;
      5713: inst = 32'hc404d38;
      5714: inst = 32'h8220000;
      5715: inst = 32'h10408000;
      5716: inst = 32'hc404d39;
      5717: inst = 32'h8220000;
      5718: inst = 32'h10408000;
      5719: inst = 32'hc404d3a;
      5720: inst = 32'h8220000;
      5721: inst = 32'h10408000;
      5722: inst = 32'hc404d3b;
      5723: inst = 32'h8220000;
      5724: inst = 32'h10408000;
      5725: inst = 32'hc404d3c;
      5726: inst = 32'h8220000;
      5727: inst = 32'h10408000;
      5728: inst = 32'hc404d3d;
      5729: inst = 32'h8220000;
      5730: inst = 32'h10408000;
      5731: inst = 32'hc404d3e;
      5732: inst = 32'h8220000;
      5733: inst = 32'h10408000;
      5734: inst = 32'hc404d3f;
      5735: inst = 32'h8220000;
      5736: inst = 32'h10408000;
      5737: inst = 32'hc404d40;
      5738: inst = 32'h8220000;
      5739: inst = 32'h10408000;
      5740: inst = 32'hc404d41;
      5741: inst = 32'h8220000;
      5742: inst = 32'h10408000;
      5743: inst = 32'hc404d42;
      5744: inst = 32'h8220000;
      5745: inst = 32'h10408000;
      5746: inst = 32'hc404d43;
      5747: inst = 32'h8220000;
      5748: inst = 32'h10408000;
      5749: inst = 32'hc404d44;
      5750: inst = 32'h8220000;
      5751: inst = 32'h10408000;
      5752: inst = 32'hc404d45;
      5753: inst = 32'h8220000;
      5754: inst = 32'h10408000;
      5755: inst = 32'hc404d46;
      5756: inst = 32'h8220000;
      5757: inst = 32'h10408000;
      5758: inst = 32'hc404d47;
      5759: inst = 32'h8220000;
      5760: inst = 32'h10408000;
      5761: inst = 32'hc404d48;
      5762: inst = 32'h8220000;
      5763: inst = 32'h10408000;
      5764: inst = 32'hc404d49;
      5765: inst = 32'h8220000;
      5766: inst = 32'h10408000;
      5767: inst = 32'hc404d4a;
      5768: inst = 32'h8220000;
      5769: inst = 32'h10408000;
      5770: inst = 32'hc404d4b;
      5771: inst = 32'h8220000;
      5772: inst = 32'h10408000;
      5773: inst = 32'hc404d4c;
      5774: inst = 32'h8220000;
      5775: inst = 32'h10408000;
      5776: inst = 32'hc404d4d;
      5777: inst = 32'h8220000;
      5778: inst = 32'h10408000;
      5779: inst = 32'hc404d4e;
      5780: inst = 32'h8220000;
      5781: inst = 32'h10408000;
      5782: inst = 32'hc404d77;
      5783: inst = 32'h8220000;
      5784: inst = 32'h10408000;
      5785: inst = 32'hc404d78;
      5786: inst = 32'h8220000;
      5787: inst = 32'h10408000;
      5788: inst = 32'hc404d79;
      5789: inst = 32'h8220000;
      5790: inst = 32'h10408000;
      5791: inst = 32'hc404d7a;
      5792: inst = 32'h8220000;
      5793: inst = 32'h10408000;
      5794: inst = 32'hc404d7b;
      5795: inst = 32'h8220000;
      5796: inst = 32'h10408000;
      5797: inst = 32'hc404d7c;
      5798: inst = 32'h8220000;
      5799: inst = 32'h10408000;
      5800: inst = 32'hc404d7d;
      5801: inst = 32'h8220000;
      5802: inst = 32'h10408000;
      5803: inst = 32'hc404d7e;
      5804: inst = 32'h8220000;
      5805: inst = 32'h10408000;
      5806: inst = 32'hc404d7f;
      5807: inst = 32'h8220000;
      5808: inst = 32'h10408000;
      5809: inst = 32'hc404d80;
      5810: inst = 32'h8220000;
      5811: inst = 32'h10408000;
      5812: inst = 32'hc404d81;
      5813: inst = 32'h8220000;
      5814: inst = 32'h10408000;
      5815: inst = 32'hc404d82;
      5816: inst = 32'h8220000;
      5817: inst = 32'h10408000;
      5818: inst = 32'hc404d83;
      5819: inst = 32'h8220000;
      5820: inst = 32'h10408000;
      5821: inst = 32'hc404d84;
      5822: inst = 32'h8220000;
      5823: inst = 32'h10408000;
      5824: inst = 32'hc404d85;
      5825: inst = 32'h8220000;
      5826: inst = 32'h10408000;
      5827: inst = 32'hc404d86;
      5828: inst = 32'h8220000;
      5829: inst = 32'h10408000;
      5830: inst = 32'hc404d87;
      5831: inst = 32'h8220000;
      5832: inst = 32'h10408000;
      5833: inst = 32'hc404d88;
      5834: inst = 32'h8220000;
      5835: inst = 32'h10408000;
      5836: inst = 32'hc404d89;
      5837: inst = 32'h8220000;
      5838: inst = 32'h10408000;
      5839: inst = 32'hc404d8a;
      5840: inst = 32'h8220000;
      5841: inst = 32'h10408000;
      5842: inst = 32'hc404d8b;
      5843: inst = 32'h8220000;
      5844: inst = 32'h10408000;
      5845: inst = 32'hc404d8c;
      5846: inst = 32'h8220000;
      5847: inst = 32'h10408000;
      5848: inst = 32'hc404d8d;
      5849: inst = 32'h8220000;
      5850: inst = 32'h10408000;
      5851: inst = 32'hc404d8e;
      5852: inst = 32'h8220000;
      5853: inst = 32'h10408000;
      5854: inst = 32'hc404d8f;
      5855: inst = 32'h8220000;
      5856: inst = 32'h10408000;
      5857: inst = 32'hc404d90;
      5858: inst = 32'h8220000;
      5859: inst = 32'h10408000;
      5860: inst = 32'hc404d91;
      5861: inst = 32'h8220000;
      5862: inst = 32'h10408000;
      5863: inst = 32'hc404d92;
      5864: inst = 32'h8220000;
      5865: inst = 32'h10408000;
      5866: inst = 32'hc404d93;
      5867: inst = 32'h8220000;
      5868: inst = 32'h10408000;
      5869: inst = 32'hc404d94;
      5870: inst = 32'h8220000;
      5871: inst = 32'h10408000;
      5872: inst = 32'hc404d95;
      5873: inst = 32'h8220000;
      5874: inst = 32'h10408000;
      5875: inst = 32'hc404d96;
      5876: inst = 32'h8220000;
      5877: inst = 32'h10408000;
      5878: inst = 32'hc404d97;
      5879: inst = 32'h8220000;
      5880: inst = 32'h10408000;
      5881: inst = 32'hc404d98;
      5882: inst = 32'h8220000;
      5883: inst = 32'h10408000;
      5884: inst = 32'hc404d99;
      5885: inst = 32'h8220000;
      5886: inst = 32'h10408000;
      5887: inst = 32'hc404d9a;
      5888: inst = 32'h8220000;
      5889: inst = 32'h10408000;
      5890: inst = 32'hc404d9b;
      5891: inst = 32'h8220000;
      5892: inst = 32'h10408000;
      5893: inst = 32'hc404d9c;
      5894: inst = 32'h8220000;
      5895: inst = 32'h10408000;
      5896: inst = 32'hc404d9d;
      5897: inst = 32'h8220000;
      5898: inst = 32'h10408000;
      5899: inst = 32'hc404d9e;
      5900: inst = 32'h8220000;
      5901: inst = 32'h10408000;
      5902: inst = 32'hc404d9f;
      5903: inst = 32'h8220000;
      5904: inst = 32'h10408000;
      5905: inst = 32'hc404da0;
      5906: inst = 32'h8220000;
      5907: inst = 32'h10408000;
      5908: inst = 32'hc404da1;
      5909: inst = 32'h8220000;
      5910: inst = 32'h10408000;
      5911: inst = 32'hc404da2;
      5912: inst = 32'h8220000;
      5913: inst = 32'h10408000;
      5914: inst = 32'hc404da3;
      5915: inst = 32'h8220000;
      5916: inst = 32'h10408000;
      5917: inst = 32'hc404da4;
      5918: inst = 32'h8220000;
      5919: inst = 32'h10408000;
      5920: inst = 32'hc404da5;
      5921: inst = 32'h8220000;
      5922: inst = 32'h10408000;
      5923: inst = 32'hc404da6;
      5924: inst = 32'h8220000;
      5925: inst = 32'h10408000;
      5926: inst = 32'hc404da7;
      5927: inst = 32'h8220000;
      5928: inst = 32'h10408000;
      5929: inst = 32'hc404da8;
      5930: inst = 32'h8220000;
      5931: inst = 32'h10408000;
      5932: inst = 32'hc404da9;
      5933: inst = 32'h8220000;
      5934: inst = 32'h10408000;
      5935: inst = 32'hc404daa;
      5936: inst = 32'h8220000;
      5937: inst = 32'h10408000;
      5938: inst = 32'hc404dab;
      5939: inst = 32'h8220000;
      5940: inst = 32'h10408000;
      5941: inst = 32'hc404dac;
      5942: inst = 32'h8220000;
      5943: inst = 32'h10408000;
      5944: inst = 32'hc404dad;
      5945: inst = 32'h8220000;
      5946: inst = 32'h10408000;
      5947: inst = 32'hc404dae;
      5948: inst = 32'h8220000;
      5949: inst = 32'h10408000;
      5950: inst = 32'hc404dd7;
      5951: inst = 32'h8220000;
      5952: inst = 32'h10408000;
      5953: inst = 32'hc404dd8;
      5954: inst = 32'h8220000;
      5955: inst = 32'h10408000;
      5956: inst = 32'hc404dd9;
      5957: inst = 32'h8220000;
      5958: inst = 32'h10408000;
      5959: inst = 32'hc404dda;
      5960: inst = 32'h8220000;
      5961: inst = 32'h10408000;
      5962: inst = 32'hc404ddb;
      5963: inst = 32'h8220000;
      5964: inst = 32'h10408000;
      5965: inst = 32'hc404ddc;
      5966: inst = 32'h8220000;
      5967: inst = 32'h10408000;
      5968: inst = 32'hc404ddd;
      5969: inst = 32'h8220000;
      5970: inst = 32'h10408000;
      5971: inst = 32'hc404dde;
      5972: inst = 32'h8220000;
      5973: inst = 32'h10408000;
      5974: inst = 32'hc404ddf;
      5975: inst = 32'h8220000;
      5976: inst = 32'h10408000;
      5977: inst = 32'hc404de0;
      5978: inst = 32'h8220000;
      5979: inst = 32'h10408000;
      5980: inst = 32'hc404de1;
      5981: inst = 32'h8220000;
      5982: inst = 32'h10408000;
      5983: inst = 32'hc404de2;
      5984: inst = 32'h8220000;
      5985: inst = 32'h10408000;
      5986: inst = 32'hc404de3;
      5987: inst = 32'h8220000;
      5988: inst = 32'h10408000;
      5989: inst = 32'hc404de4;
      5990: inst = 32'h8220000;
      5991: inst = 32'h10408000;
      5992: inst = 32'hc404de5;
      5993: inst = 32'h8220000;
      5994: inst = 32'h10408000;
      5995: inst = 32'hc404de6;
      5996: inst = 32'h8220000;
      5997: inst = 32'h10408000;
      5998: inst = 32'hc404de7;
      5999: inst = 32'h8220000;
      6000: inst = 32'h10408000;
      6001: inst = 32'hc404de8;
      6002: inst = 32'h8220000;
      6003: inst = 32'h10408000;
      6004: inst = 32'hc404de9;
      6005: inst = 32'h8220000;
      6006: inst = 32'h10408000;
      6007: inst = 32'hc404dea;
      6008: inst = 32'h8220000;
      6009: inst = 32'h10408000;
      6010: inst = 32'hc404deb;
      6011: inst = 32'h8220000;
      6012: inst = 32'h10408000;
      6013: inst = 32'hc404dec;
      6014: inst = 32'h8220000;
      6015: inst = 32'h10408000;
      6016: inst = 32'hc404ded;
      6017: inst = 32'h8220000;
      6018: inst = 32'h10408000;
      6019: inst = 32'hc404dee;
      6020: inst = 32'h8220000;
      6021: inst = 32'h10408000;
      6022: inst = 32'hc404def;
      6023: inst = 32'h8220000;
      6024: inst = 32'h10408000;
      6025: inst = 32'hc404df0;
      6026: inst = 32'h8220000;
      6027: inst = 32'h10408000;
      6028: inst = 32'hc404df1;
      6029: inst = 32'h8220000;
      6030: inst = 32'h10408000;
      6031: inst = 32'hc404df2;
      6032: inst = 32'h8220000;
      6033: inst = 32'h10408000;
      6034: inst = 32'hc404df3;
      6035: inst = 32'h8220000;
      6036: inst = 32'h10408000;
      6037: inst = 32'hc404df4;
      6038: inst = 32'h8220000;
      6039: inst = 32'h10408000;
      6040: inst = 32'hc404df5;
      6041: inst = 32'h8220000;
      6042: inst = 32'h10408000;
      6043: inst = 32'hc404df6;
      6044: inst = 32'h8220000;
      6045: inst = 32'h10408000;
      6046: inst = 32'hc404df7;
      6047: inst = 32'h8220000;
      6048: inst = 32'h10408000;
      6049: inst = 32'hc404df8;
      6050: inst = 32'h8220000;
      6051: inst = 32'h10408000;
      6052: inst = 32'hc404df9;
      6053: inst = 32'h8220000;
      6054: inst = 32'h10408000;
      6055: inst = 32'hc404dfa;
      6056: inst = 32'h8220000;
      6057: inst = 32'h10408000;
      6058: inst = 32'hc404dfb;
      6059: inst = 32'h8220000;
      6060: inst = 32'h10408000;
      6061: inst = 32'hc404dfc;
      6062: inst = 32'h8220000;
      6063: inst = 32'h10408000;
      6064: inst = 32'hc404dfd;
      6065: inst = 32'h8220000;
      6066: inst = 32'h10408000;
      6067: inst = 32'hc404dfe;
      6068: inst = 32'h8220000;
      6069: inst = 32'h10408000;
      6070: inst = 32'hc404dff;
      6071: inst = 32'h8220000;
      6072: inst = 32'h10408000;
      6073: inst = 32'hc404e00;
      6074: inst = 32'h8220000;
      6075: inst = 32'h10408000;
      6076: inst = 32'hc404e01;
      6077: inst = 32'h8220000;
      6078: inst = 32'h10408000;
      6079: inst = 32'hc404e02;
      6080: inst = 32'h8220000;
      6081: inst = 32'h10408000;
      6082: inst = 32'hc404e03;
      6083: inst = 32'h8220000;
      6084: inst = 32'h10408000;
      6085: inst = 32'hc404e04;
      6086: inst = 32'h8220000;
      6087: inst = 32'h10408000;
      6088: inst = 32'hc404e05;
      6089: inst = 32'h8220000;
      6090: inst = 32'h10408000;
      6091: inst = 32'hc404e06;
      6092: inst = 32'h8220000;
      6093: inst = 32'h10408000;
      6094: inst = 32'hc404e07;
      6095: inst = 32'h8220000;
      6096: inst = 32'h10408000;
      6097: inst = 32'hc404e08;
      6098: inst = 32'h8220000;
      6099: inst = 32'h10408000;
      6100: inst = 32'hc404e09;
      6101: inst = 32'h8220000;
      6102: inst = 32'h10408000;
      6103: inst = 32'hc404e0a;
      6104: inst = 32'h8220000;
      6105: inst = 32'h10408000;
      6106: inst = 32'hc404e0b;
      6107: inst = 32'h8220000;
      6108: inst = 32'h10408000;
      6109: inst = 32'hc404e0c;
      6110: inst = 32'h8220000;
      6111: inst = 32'h10408000;
      6112: inst = 32'hc404e0d;
      6113: inst = 32'h8220000;
      6114: inst = 32'h10408000;
      6115: inst = 32'hc404e0e;
      6116: inst = 32'h8220000;
      6117: inst = 32'h10408000;
      6118: inst = 32'hc404e37;
      6119: inst = 32'h8220000;
      6120: inst = 32'h10408000;
      6121: inst = 32'hc404e38;
      6122: inst = 32'h8220000;
      6123: inst = 32'h10408000;
      6124: inst = 32'hc404e39;
      6125: inst = 32'h8220000;
      6126: inst = 32'h10408000;
      6127: inst = 32'hc404e3a;
      6128: inst = 32'h8220000;
      6129: inst = 32'h10408000;
      6130: inst = 32'hc404e3b;
      6131: inst = 32'h8220000;
      6132: inst = 32'h10408000;
      6133: inst = 32'hc404e3c;
      6134: inst = 32'h8220000;
      6135: inst = 32'h10408000;
      6136: inst = 32'hc404e3d;
      6137: inst = 32'h8220000;
      6138: inst = 32'h10408000;
      6139: inst = 32'hc404e3e;
      6140: inst = 32'h8220000;
      6141: inst = 32'h10408000;
      6142: inst = 32'hc404e3f;
      6143: inst = 32'h8220000;
      6144: inst = 32'h10408000;
      6145: inst = 32'hc404e40;
      6146: inst = 32'h8220000;
      6147: inst = 32'h10408000;
      6148: inst = 32'hc404e41;
      6149: inst = 32'h8220000;
      6150: inst = 32'h10408000;
      6151: inst = 32'hc404e42;
      6152: inst = 32'h8220000;
      6153: inst = 32'h10408000;
      6154: inst = 32'hc404e43;
      6155: inst = 32'h8220000;
      6156: inst = 32'h10408000;
      6157: inst = 32'hc404e44;
      6158: inst = 32'h8220000;
      6159: inst = 32'h10408000;
      6160: inst = 32'hc404e45;
      6161: inst = 32'h8220000;
      6162: inst = 32'h10408000;
      6163: inst = 32'hc404e46;
      6164: inst = 32'h8220000;
      6165: inst = 32'h10408000;
      6166: inst = 32'hc404e47;
      6167: inst = 32'h8220000;
      6168: inst = 32'h10408000;
      6169: inst = 32'hc404e48;
      6170: inst = 32'h8220000;
      6171: inst = 32'h10408000;
      6172: inst = 32'hc404e49;
      6173: inst = 32'h8220000;
      6174: inst = 32'h10408000;
      6175: inst = 32'hc404e4a;
      6176: inst = 32'h8220000;
      6177: inst = 32'h10408000;
      6178: inst = 32'hc404e4b;
      6179: inst = 32'h8220000;
      6180: inst = 32'h10408000;
      6181: inst = 32'hc404e4c;
      6182: inst = 32'h8220000;
      6183: inst = 32'h10408000;
      6184: inst = 32'hc404e4d;
      6185: inst = 32'h8220000;
      6186: inst = 32'h10408000;
      6187: inst = 32'hc404e4e;
      6188: inst = 32'h8220000;
      6189: inst = 32'h10408000;
      6190: inst = 32'hc404e4f;
      6191: inst = 32'h8220000;
      6192: inst = 32'h10408000;
      6193: inst = 32'hc404e50;
      6194: inst = 32'h8220000;
      6195: inst = 32'h10408000;
      6196: inst = 32'hc404e51;
      6197: inst = 32'h8220000;
      6198: inst = 32'h10408000;
      6199: inst = 32'hc404e52;
      6200: inst = 32'h8220000;
      6201: inst = 32'h10408000;
      6202: inst = 32'hc404e53;
      6203: inst = 32'h8220000;
      6204: inst = 32'h10408000;
      6205: inst = 32'hc404e54;
      6206: inst = 32'h8220000;
      6207: inst = 32'h10408000;
      6208: inst = 32'hc404e55;
      6209: inst = 32'h8220000;
      6210: inst = 32'h10408000;
      6211: inst = 32'hc404e56;
      6212: inst = 32'h8220000;
      6213: inst = 32'h10408000;
      6214: inst = 32'hc404e57;
      6215: inst = 32'h8220000;
      6216: inst = 32'h10408000;
      6217: inst = 32'hc404e58;
      6218: inst = 32'h8220000;
      6219: inst = 32'h10408000;
      6220: inst = 32'hc404e59;
      6221: inst = 32'h8220000;
      6222: inst = 32'h10408000;
      6223: inst = 32'hc404e5a;
      6224: inst = 32'h8220000;
      6225: inst = 32'h10408000;
      6226: inst = 32'hc404e5b;
      6227: inst = 32'h8220000;
      6228: inst = 32'h10408000;
      6229: inst = 32'hc404e5c;
      6230: inst = 32'h8220000;
      6231: inst = 32'h10408000;
      6232: inst = 32'hc404e5d;
      6233: inst = 32'h8220000;
      6234: inst = 32'h10408000;
      6235: inst = 32'hc404e5e;
      6236: inst = 32'h8220000;
      6237: inst = 32'h10408000;
      6238: inst = 32'hc404e5f;
      6239: inst = 32'h8220000;
      6240: inst = 32'h10408000;
      6241: inst = 32'hc404e60;
      6242: inst = 32'h8220000;
      6243: inst = 32'h10408000;
      6244: inst = 32'hc404e61;
      6245: inst = 32'h8220000;
      6246: inst = 32'h10408000;
      6247: inst = 32'hc404e62;
      6248: inst = 32'h8220000;
      6249: inst = 32'h10408000;
      6250: inst = 32'hc404e63;
      6251: inst = 32'h8220000;
      6252: inst = 32'h10408000;
      6253: inst = 32'hc404e64;
      6254: inst = 32'h8220000;
      6255: inst = 32'h10408000;
      6256: inst = 32'hc404e65;
      6257: inst = 32'h8220000;
      6258: inst = 32'h10408000;
      6259: inst = 32'hc404e66;
      6260: inst = 32'h8220000;
      6261: inst = 32'h10408000;
      6262: inst = 32'hc404e67;
      6263: inst = 32'h8220000;
      6264: inst = 32'h10408000;
      6265: inst = 32'hc404e68;
      6266: inst = 32'h8220000;
      6267: inst = 32'h10408000;
      6268: inst = 32'hc404e69;
      6269: inst = 32'h8220000;
      6270: inst = 32'h10408000;
      6271: inst = 32'hc404e6a;
      6272: inst = 32'h8220000;
      6273: inst = 32'h10408000;
      6274: inst = 32'hc404e6b;
      6275: inst = 32'h8220000;
      6276: inst = 32'h10408000;
      6277: inst = 32'hc404e6c;
      6278: inst = 32'h8220000;
      6279: inst = 32'h10408000;
      6280: inst = 32'hc404e6d;
      6281: inst = 32'h8220000;
      6282: inst = 32'h10408000;
      6283: inst = 32'hc404e6e;
      6284: inst = 32'h8220000;
      6285: inst = 32'h10408000;
      6286: inst = 32'hc404e97;
      6287: inst = 32'h8220000;
      6288: inst = 32'h10408000;
      6289: inst = 32'hc404e98;
      6290: inst = 32'h8220000;
      6291: inst = 32'h10408000;
      6292: inst = 32'hc404e99;
      6293: inst = 32'h8220000;
      6294: inst = 32'h10408000;
      6295: inst = 32'hc404e9a;
      6296: inst = 32'h8220000;
      6297: inst = 32'h10408000;
      6298: inst = 32'hc404e9b;
      6299: inst = 32'h8220000;
      6300: inst = 32'h10408000;
      6301: inst = 32'hc404e9c;
      6302: inst = 32'h8220000;
      6303: inst = 32'h10408000;
      6304: inst = 32'hc404e9d;
      6305: inst = 32'h8220000;
      6306: inst = 32'h10408000;
      6307: inst = 32'hc404e9e;
      6308: inst = 32'h8220000;
      6309: inst = 32'h10408000;
      6310: inst = 32'hc404ea8;
      6311: inst = 32'h8220000;
      6312: inst = 32'h10408000;
      6313: inst = 32'hc404ea9;
      6314: inst = 32'h8220000;
      6315: inst = 32'h10408000;
      6316: inst = 32'hc404eaa;
      6317: inst = 32'h8220000;
      6318: inst = 32'h10408000;
      6319: inst = 32'hc404eab;
      6320: inst = 32'h8220000;
      6321: inst = 32'h10408000;
      6322: inst = 32'hc404eac;
      6323: inst = 32'h8220000;
      6324: inst = 32'h10408000;
      6325: inst = 32'hc404ead;
      6326: inst = 32'h8220000;
      6327: inst = 32'h10408000;
      6328: inst = 32'hc404eae;
      6329: inst = 32'h8220000;
      6330: inst = 32'h10408000;
      6331: inst = 32'hc404eaf;
      6332: inst = 32'h8220000;
      6333: inst = 32'h10408000;
      6334: inst = 32'hc404eb0;
      6335: inst = 32'h8220000;
      6336: inst = 32'h10408000;
      6337: inst = 32'hc404eb1;
      6338: inst = 32'h8220000;
      6339: inst = 32'h10408000;
      6340: inst = 32'hc404eb2;
      6341: inst = 32'h8220000;
      6342: inst = 32'h10408000;
      6343: inst = 32'hc404eb3;
      6344: inst = 32'h8220000;
      6345: inst = 32'h10408000;
      6346: inst = 32'hc404eb4;
      6347: inst = 32'h8220000;
      6348: inst = 32'h10408000;
      6349: inst = 32'hc404eb5;
      6350: inst = 32'h8220000;
      6351: inst = 32'h10408000;
      6352: inst = 32'hc404eb6;
      6353: inst = 32'h8220000;
      6354: inst = 32'h10408000;
      6355: inst = 32'hc404eb7;
      6356: inst = 32'h8220000;
      6357: inst = 32'h10408000;
      6358: inst = 32'hc404ec1;
      6359: inst = 32'h8220000;
      6360: inst = 32'h10408000;
      6361: inst = 32'hc404ec2;
      6362: inst = 32'h8220000;
      6363: inst = 32'h10408000;
      6364: inst = 32'hc404ec3;
      6365: inst = 32'h8220000;
      6366: inst = 32'h10408000;
      6367: inst = 32'hc404ec4;
      6368: inst = 32'h8220000;
      6369: inst = 32'h10408000;
      6370: inst = 32'hc404ec5;
      6371: inst = 32'h8220000;
      6372: inst = 32'h10408000;
      6373: inst = 32'hc404ec6;
      6374: inst = 32'h8220000;
      6375: inst = 32'h10408000;
      6376: inst = 32'hc404ec7;
      6377: inst = 32'h8220000;
      6378: inst = 32'h10408000;
      6379: inst = 32'hc404ec8;
      6380: inst = 32'h8220000;
      6381: inst = 32'h10408000;
      6382: inst = 32'hc404ec9;
      6383: inst = 32'h8220000;
      6384: inst = 32'h10408000;
      6385: inst = 32'hc404eca;
      6386: inst = 32'h8220000;
      6387: inst = 32'h10408000;
      6388: inst = 32'hc404ecb;
      6389: inst = 32'h8220000;
      6390: inst = 32'h10408000;
      6391: inst = 32'hc404ecc;
      6392: inst = 32'h8220000;
      6393: inst = 32'h10408000;
      6394: inst = 32'hc404ecd;
      6395: inst = 32'h8220000;
      6396: inst = 32'h10408000;
      6397: inst = 32'hc404ece;
      6398: inst = 32'h8220000;
      6399: inst = 32'h10408000;
      6400: inst = 32'hc404ef7;
      6401: inst = 32'h8220000;
      6402: inst = 32'h10408000;
      6403: inst = 32'hc404ef8;
      6404: inst = 32'h8220000;
      6405: inst = 32'h10408000;
      6406: inst = 32'hc404ef9;
      6407: inst = 32'h8220000;
      6408: inst = 32'h10408000;
      6409: inst = 32'hc404efa;
      6410: inst = 32'h8220000;
      6411: inst = 32'h10408000;
      6412: inst = 32'hc404efb;
      6413: inst = 32'h8220000;
      6414: inst = 32'h10408000;
      6415: inst = 32'hc404efc;
      6416: inst = 32'h8220000;
      6417: inst = 32'h10408000;
      6418: inst = 32'hc404efd;
      6419: inst = 32'h8220000;
      6420: inst = 32'h10408000;
      6421: inst = 32'hc404efe;
      6422: inst = 32'h8220000;
      6423: inst = 32'h10408000;
      6424: inst = 32'hc404f08;
      6425: inst = 32'h8220000;
      6426: inst = 32'h10408000;
      6427: inst = 32'hc404f09;
      6428: inst = 32'h8220000;
      6429: inst = 32'h10408000;
      6430: inst = 32'hc404f0a;
      6431: inst = 32'h8220000;
      6432: inst = 32'h10408000;
      6433: inst = 32'hc404f0b;
      6434: inst = 32'h8220000;
      6435: inst = 32'h10408000;
      6436: inst = 32'hc404f0c;
      6437: inst = 32'h8220000;
      6438: inst = 32'h10408000;
      6439: inst = 32'hc404f0d;
      6440: inst = 32'h8220000;
      6441: inst = 32'h10408000;
      6442: inst = 32'hc404f0e;
      6443: inst = 32'h8220000;
      6444: inst = 32'h10408000;
      6445: inst = 32'hc404f0f;
      6446: inst = 32'h8220000;
      6447: inst = 32'h10408000;
      6448: inst = 32'hc404f10;
      6449: inst = 32'h8220000;
      6450: inst = 32'h10408000;
      6451: inst = 32'hc404f11;
      6452: inst = 32'h8220000;
      6453: inst = 32'h10408000;
      6454: inst = 32'hc404f12;
      6455: inst = 32'h8220000;
      6456: inst = 32'h10408000;
      6457: inst = 32'hc404f13;
      6458: inst = 32'h8220000;
      6459: inst = 32'h10408000;
      6460: inst = 32'hc404f14;
      6461: inst = 32'h8220000;
      6462: inst = 32'h10408000;
      6463: inst = 32'hc404f15;
      6464: inst = 32'h8220000;
      6465: inst = 32'h10408000;
      6466: inst = 32'hc404f16;
      6467: inst = 32'h8220000;
      6468: inst = 32'h10408000;
      6469: inst = 32'hc404f17;
      6470: inst = 32'h8220000;
      6471: inst = 32'h10408000;
      6472: inst = 32'hc404f21;
      6473: inst = 32'h8220000;
      6474: inst = 32'h10408000;
      6475: inst = 32'hc404f22;
      6476: inst = 32'h8220000;
      6477: inst = 32'h10408000;
      6478: inst = 32'hc404f23;
      6479: inst = 32'h8220000;
      6480: inst = 32'h10408000;
      6481: inst = 32'hc404f24;
      6482: inst = 32'h8220000;
      6483: inst = 32'h10408000;
      6484: inst = 32'hc404f25;
      6485: inst = 32'h8220000;
      6486: inst = 32'h10408000;
      6487: inst = 32'hc404f26;
      6488: inst = 32'h8220000;
      6489: inst = 32'h10408000;
      6490: inst = 32'hc404f27;
      6491: inst = 32'h8220000;
      6492: inst = 32'h10408000;
      6493: inst = 32'hc404f28;
      6494: inst = 32'h8220000;
      6495: inst = 32'h10408000;
      6496: inst = 32'hc404f29;
      6497: inst = 32'h8220000;
      6498: inst = 32'h10408000;
      6499: inst = 32'hc404f2a;
      6500: inst = 32'h8220000;
      6501: inst = 32'h10408000;
      6502: inst = 32'hc404f2b;
      6503: inst = 32'h8220000;
      6504: inst = 32'h10408000;
      6505: inst = 32'hc404f2c;
      6506: inst = 32'h8220000;
      6507: inst = 32'h10408000;
      6508: inst = 32'hc404f2d;
      6509: inst = 32'h8220000;
      6510: inst = 32'h10408000;
      6511: inst = 32'hc404f2e;
      6512: inst = 32'h8220000;
      6513: inst = 32'h10408000;
      6514: inst = 32'hc404f57;
      6515: inst = 32'h8220000;
      6516: inst = 32'h10408000;
      6517: inst = 32'hc404f58;
      6518: inst = 32'h8220000;
      6519: inst = 32'h10408000;
      6520: inst = 32'hc404f59;
      6521: inst = 32'h8220000;
      6522: inst = 32'h10408000;
      6523: inst = 32'hc404f5a;
      6524: inst = 32'h8220000;
      6525: inst = 32'h10408000;
      6526: inst = 32'hc404f5b;
      6527: inst = 32'h8220000;
      6528: inst = 32'h10408000;
      6529: inst = 32'hc404f5c;
      6530: inst = 32'h8220000;
      6531: inst = 32'h10408000;
      6532: inst = 32'hc404f5d;
      6533: inst = 32'h8220000;
      6534: inst = 32'h10408000;
      6535: inst = 32'hc404f5e;
      6536: inst = 32'h8220000;
      6537: inst = 32'h10408000;
      6538: inst = 32'hc404f68;
      6539: inst = 32'h8220000;
      6540: inst = 32'h10408000;
      6541: inst = 32'hc404f69;
      6542: inst = 32'h8220000;
      6543: inst = 32'h10408000;
      6544: inst = 32'hc404f6a;
      6545: inst = 32'h8220000;
      6546: inst = 32'h10408000;
      6547: inst = 32'hc404f6b;
      6548: inst = 32'h8220000;
      6549: inst = 32'h10408000;
      6550: inst = 32'hc404f6c;
      6551: inst = 32'h8220000;
      6552: inst = 32'h10408000;
      6553: inst = 32'hc404f6d;
      6554: inst = 32'h8220000;
      6555: inst = 32'h10408000;
      6556: inst = 32'hc404f6e;
      6557: inst = 32'h8220000;
      6558: inst = 32'h10408000;
      6559: inst = 32'hc404f6f;
      6560: inst = 32'h8220000;
      6561: inst = 32'h10408000;
      6562: inst = 32'hc404f70;
      6563: inst = 32'h8220000;
      6564: inst = 32'h10408000;
      6565: inst = 32'hc404f71;
      6566: inst = 32'h8220000;
      6567: inst = 32'h10408000;
      6568: inst = 32'hc404f72;
      6569: inst = 32'h8220000;
      6570: inst = 32'h10408000;
      6571: inst = 32'hc404f73;
      6572: inst = 32'h8220000;
      6573: inst = 32'h10408000;
      6574: inst = 32'hc404f74;
      6575: inst = 32'h8220000;
      6576: inst = 32'h10408000;
      6577: inst = 32'hc404f75;
      6578: inst = 32'h8220000;
      6579: inst = 32'h10408000;
      6580: inst = 32'hc404f76;
      6581: inst = 32'h8220000;
      6582: inst = 32'h10408000;
      6583: inst = 32'hc404f77;
      6584: inst = 32'h8220000;
      6585: inst = 32'h10408000;
      6586: inst = 32'hc404f81;
      6587: inst = 32'h8220000;
      6588: inst = 32'h10408000;
      6589: inst = 32'hc404f82;
      6590: inst = 32'h8220000;
      6591: inst = 32'h10408000;
      6592: inst = 32'hc404f83;
      6593: inst = 32'h8220000;
      6594: inst = 32'h10408000;
      6595: inst = 32'hc404f84;
      6596: inst = 32'h8220000;
      6597: inst = 32'h10408000;
      6598: inst = 32'hc404f85;
      6599: inst = 32'h8220000;
      6600: inst = 32'h10408000;
      6601: inst = 32'hc404f86;
      6602: inst = 32'h8220000;
      6603: inst = 32'h10408000;
      6604: inst = 32'hc404f87;
      6605: inst = 32'h8220000;
      6606: inst = 32'h10408000;
      6607: inst = 32'hc404f88;
      6608: inst = 32'h8220000;
      6609: inst = 32'h10408000;
      6610: inst = 32'hc404f89;
      6611: inst = 32'h8220000;
      6612: inst = 32'h10408000;
      6613: inst = 32'hc404f8a;
      6614: inst = 32'h8220000;
      6615: inst = 32'h10408000;
      6616: inst = 32'hc404f8b;
      6617: inst = 32'h8220000;
      6618: inst = 32'h10408000;
      6619: inst = 32'hc404f8c;
      6620: inst = 32'h8220000;
      6621: inst = 32'h10408000;
      6622: inst = 32'hc404f8d;
      6623: inst = 32'h8220000;
      6624: inst = 32'h10408000;
      6625: inst = 32'hc404f8e;
      6626: inst = 32'h8220000;
      6627: inst = 32'h10408000;
      6628: inst = 32'hc404fb7;
      6629: inst = 32'h8220000;
      6630: inst = 32'h10408000;
      6631: inst = 32'hc404fb8;
      6632: inst = 32'h8220000;
      6633: inst = 32'h10408000;
      6634: inst = 32'hc404fb9;
      6635: inst = 32'h8220000;
      6636: inst = 32'h10408000;
      6637: inst = 32'hc404fba;
      6638: inst = 32'h8220000;
      6639: inst = 32'h10408000;
      6640: inst = 32'hc404fbb;
      6641: inst = 32'h8220000;
      6642: inst = 32'h10408000;
      6643: inst = 32'hc404fbc;
      6644: inst = 32'h8220000;
      6645: inst = 32'h10408000;
      6646: inst = 32'hc404fbd;
      6647: inst = 32'h8220000;
      6648: inst = 32'h10408000;
      6649: inst = 32'hc404fbe;
      6650: inst = 32'h8220000;
      6651: inst = 32'h10408000;
      6652: inst = 32'hc404fc8;
      6653: inst = 32'h8220000;
      6654: inst = 32'h10408000;
      6655: inst = 32'hc404fc9;
      6656: inst = 32'h8220000;
      6657: inst = 32'h10408000;
      6658: inst = 32'hc404fca;
      6659: inst = 32'h8220000;
      6660: inst = 32'h10408000;
      6661: inst = 32'hc404fcb;
      6662: inst = 32'h8220000;
      6663: inst = 32'h10408000;
      6664: inst = 32'hc404fcc;
      6665: inst = 32'h8220000;
      6666: inst = 32'h10408000;
      6667: inst = 32'hc404fcd;
      6668: inst = 32'h8220000;
      6669: inst = 32'h10408000;
      6670: inst = 32'hc404fce;
      6671: inst = 32'h8220000;
      6672: inst = 32'h10408000;
      6673: inst = 32'hc404fcf;
      6674: inst = 32'h8220000;
      6675: inst = 32'h10408000;
      6676: inst = 32'hc404fd0;
      6677: inst = 32'h8220000;
      6678: inst = 32'h10408000;
      6679: inst = 32'hc404fd1;
      6680: inst = 32'h8220000;
      6681: inst = 32'h10408000;
      6682: inst = 32'hc404fd2;
      6683: inst = 32'h8220000;
      6684: inst = 32'h10408000;
      6685: inst = 32'hc404fd3;
      6686: inst = 32'h8220000;
      6687: inst = 32'h10408000;
      6688: inst = 32'hc404fd4;
      6689: inst = 32'h8220000;
      6690: inst = 32'h10408000;
      6691: inst = 32'hc404fd5;
      6692: inst = 32'h8220000;
      6693: inst = 32'h10408000;
      6694: inst = 32'hc404fd6;
      6695: inst = 32'h8220000;
      6696: inst = 32'h10408000;
      6697: inst = 32'hc404fd7;
      6698: inst = 32'h8220000;
      6699: inst = 32'h10408000;
      6700: inst = 32'hc404fe1;
      6701: inst = 32'h8220000;
      6702: inst = 32'h10408000;
      6703: inst = 32'hc404fe2;
      6704: inst = 32'h8220000;
      6705: inst = 32'h10408000;
      6706: inst = 32'hc404fe3;
      6707: inst = 32'h8220000;
      6708: inst = 32'h10408000;
      6709: inst = 32'hc404fe4;
      6710: inst = 32'h8220000;
      6711: inst = 32'h10408000;
      6712: inst = 32'hc404fe5;
      6713: inst = 32'h8220000;
      6714: inst = 32'h10408000;
      6715: inst = 32'hc404fe6;
      6716: inst = 32'h8220000;
      6717: inst = 32'h10408000;
      6718: inst = 32'hc404fe7;
      6719: inst = 32'h8220000;
      6720: inst = 32'h10408000;
      6721: inst = 32'hc404fe8;
      6722: inst = 32'h8220000;
      6723: inst = 32'h10408000;
      6724: inst = 32'hc404fe9;
      6725: inst = 32'h8220000;
      6726: inst = 32'h10408000;
      6727: inst = 32'hc404fea;
      6728: inst = 32'h8220000;
      6729: inst = 32'h10408000;
      6730: inst = 32'hc404feb;
      6731: inst = 32'h8220000;
      6732: inst = 32'h10408000;
      6733: inst = 32'hc404fec;
      6734: inst = 32'h8220000;
      6735: inst = 32'h10408000;
      6736: inst = 32'hc404fed;
      6737: inst = 32'h8220000;
      6738: inst = 32'h10408000;
      6739: inst = 32'hc404fee;
      6740: inst = 32'h8220000;
      6741: inst = 32'h10408000;
      6742: inst = 32'hc405017;
      6743: inst = 32'h8220000;
      6744: inst = 32'h10408000;
      6745: inst = 32'hc405018;
      6746: inst = 32'h8220000;
      6747: inst = 32'h10408000;
      6748: inst = 32'hc405019;
      6749: inst = 32'h8220000;
      6750: inst = 32'h10408000;
      6751: inst = 32'hc40501a;
      6752: inst = 32'h8220000;
      6753: inst = 32'h10408000;
      6754: inst = 32'hc40501b;
      6755: inst = 32'h8220000;
      6756: inst = 32'h10408000;
      6757: inst = 32'hc40501c;
      6758: inst = 32'h8220000;
      6759: inst = 32'h10408000;
      6760: inst = 32'hc40501d;
      6761: inst = 32'h8220000;
      6762: inst = 32'h10408000;
      6763: inst = 32'hc40501e;
      6764: inst = 32'h8220000;
      6765: inst = 32'h10408000;
      6766: inst = 32'hc405028;
      6767: inst = 32'h8220000;
      6768: inst = 32'h10408000;
      6769: inst = 32'hc405029;
      6770: inst = 32'h8220000;
      6771: inst = 32'h10408000;
      6772: inst = 32'hc40502a;
      6773: inst = 32'h8220000;
      6774: inst = 32'h10408000;
      6775: inst = 32'hc40502b;
      6776: inst = 32'h8220000;
      6777: inst = 32'h10408000;
      6778: inst = 32'hc40502c;
      6779: inst = 32'h8220000;
      6780: inst = 32'h10408000;
      6781: inst = 32'hc40502d;
      6782: inst = 32'h8220000;
      6783: inst = 32'h10408000;
      6784: inst = 32'hc40502e;
      6785: inst = 32'h8220000;
      6786: inst = 32'h10408000;
      6787: inst = 32'hc40502f;
      6788: inst = 32'h8220000;
      6789: inst = 32'h10408000;
      6790: inst = 32'hc405030;
      6791: inst = 32'h8220000;
      6792: inst = 32'h10408000;
      6793: inst = 32'hc405031;
      6794: inst = 32'h8220000;
      6795: inst = 32'h10408000;
      6796: inst = 32'hc405032;
      6797: inst = 32'h8220000;
      6798: inst = 32'h10408000;
      6799: inst = 32'hc405033;
      6800: inst = 32'h8220000;
      6801: inst = 32'h10408000;
      6802: inst = 32'hc405034;
      6803: inst = 32'h8220000;
      6804: inst = 32'h10408000;
      6805: inst = 32'hc405035;
      6806: inst = 32'h8220000;
      6807: inst = 32'h10408000;
      6808: inst = 32'hc405036;
      6809: inst = 32'h8220000;
      6810: inst = 32'h10408000;
      6811: inst = 32'hc405037;
      6812: inst = 32'h8220000;
      6813: inst = 32'h10408000;
      6814: inst = 32'hc405041;
      6815: inst = 32'h8220000;
      6816: inst = 32'h10408000;
      6817: inst = 32'hc405042;
      6818: inst = 32'h8220000;
      6819: inst = 32'h10408000;
      6820: inst = 32'hc405043;
      6821: inst = 32'h8220000;
      6822: inst = 32'h10408000;
      6823: inst = 32'hc405044;
      6824: inst = 32'h8220000;
      6825: inst = 32'h10408000;
      6826: inst = 32'hc405045;
      6827: inst = 32'h8220000;
      6828: inst = 32'h10408000;
      6829: inst = 32'hc405046;
      6830: inst = 32'h8220000;
      6831: inst = 32'h10408000;
      6832: inst = 32'hc405047;
      6833: inst = 32'h8220000;
      6834: inst = 32'h10408000;
      6835: inst = 32'hc405048;
      6836: inst = 32'h8220000;
      6837: inst = 32'h10408000;
      6838: inst = 32'hc405049;
      6839: inst = 32'h8220000;
      6840: inst = 32'h10408000;
      6841: inst = 32'hc40504a;
      6842: inst = 32'h8220000;
      6843: inst = 32'h10408000;
      6844: inst = 32'hc40504b;
      6845: inst = 32'h8220000;
      6846: inst = 32'h10408000;
      6847: inst = 32'hc40504c;
      6848: inst = 32'h8220000;
      6849: inst = 32'h10408000;
      6850: inst = 32'hc40504d;
      6851: inst = 32'h8220000;
      6852: inst = 32'h10408000;
      6853: inst = 32'hc40504e;
      6854: inst = 32'h8220000;
      6855: inst = 32'h10408000;
      6856: inst = 32'hc405077;
      6857: inst = 32'h8220000;
      6858: inst = 32'h10408000;
      6859: inst = 32'hc405078;
      6860: inst = 32'h8220000;
      6861: inst = 32'h10408000;
      6862: inst = 32'hc405079;
      6863: inst = 32'h8220000;
      6864: inst = 32'h10408000;
      6865: inst = 32'hc40507a;
      6866: inst = 32'h8220000;
      6867: inst = 32'h10408000;
      6868: inst = 32'hc40507b;
      6869: inst = 32'h8220000;
      6870: inst = 32'h10408000;
      6871: inst = 32'hc40507c;
      6872: inst = 32'h8220000;
      6873: inst = 32'h10408000;
      6874: inst = 32'hc40507d;
      6875: inst = 32'h8220000;
      6876: inst = 32'h10408000;
      6877: inst = 32'hc40507e;
      6878: inst = 32'h8220000;
      6879: inst = 32'h10408000;
      6880: inst = 32'hc405088;
      6881: inst = 32'h8220000;
      6882: inst = 32'h10408000;
      6883: inst = 32'hc405089;
      6884: inst = 32'h8220000;
      6885: inst = 32'h10408000;
      6886: inst = 32'hc40508a;
      6887: inst = 32'h8220000;
      6888: inst = 32'h10408000;
      6889: inst = 32'hc40508b;
      6890: inst = 32'h8220000;
      6891: inst = 32'h10408000;
      6892: inst = 32'hc40508c;
      6893: inst = 32'h8220000;
      6894: inst = 32'h10408000;
      6895: inst = 32'hc40508d;
      6896: inst = 32'h8220000;
      6897: inst = 32'h10408000;
      6898: inst = 32'hc40508e;
      6899: inst = 32'h8220000;
      6900: inst = 32'h10408000;
      6901: inst = 32'hc40508f;
      6902: inst = 32'h8220000;
      6903: inst = 32'h10408000;
      6904: inst = 32'hc405090;
      6905: inst = 32'h8220000;
      6906: inst = 32'h10408000;
      6907: inst = 32'hc405091;
      6908: inst = 32'h8220000;
      6909: inst = 32'h10408000;
      6910: inst = 32'hc405092;
      6911: inst = 32'h8220000;
      6912: inst = 32'h10408000;
      6913: inst = 32'hc405093;
      6914: inst = 32'h8220000;
      6915: inst = 32'h10408000;
      6916: inst = 32'hc405094;
      6917: inst = 32'h8220000;
      6918: inst = 32'h10408000;
      6919: inst = 32'hc405095;
      6920: inst = 32'h8220000;
      6921: inst = 32'h10408000;
      6922: inst = 32'hc405096;
      6923: inst = 32'h8220000;
      6924: inst = 32'h10408000;
      6925: inst = 32'hc405097;
      6926: inst = 32'h8220000;
      6927: inst = 32'h10408000;
      6928: inst = 32'hc4050a1;
      6929: inst = 32'h8220000;
      6930: inst = 32'h10408000;
      6931: inst = 32'hc4050a2;
      6932: inst = 32'h8220000;
      6933: inst = 32'h10408000;
      6934: inst = 32'hc4050a3;
      6935: inst = 32'h8220000;
      6936: inst = 32'h10408000;
      6937: inst = 32'hc4050a4;
      6938: inst = 32'h8220000;
      6939: inst = 32'h10408000;
      6940: inst = 32'hc4050a5;
      6941: inst = 32'h8220000;
      6942: inst = 32'h10408000;
      6943: inst = 32'hc4050a6;
      6944: inst = 32'h8220000;
      6945: inst = 32'h10408000;
      6946: inst = 32'hc4050a7;
      6947: inst = 32'h8220000;
      6948: inst = 32'h10408000;
      6949: inst = 32'hc4050a8;
      6950: inst = 32'h8220000;
      6951: inst = 32'h10408000;
      6952: inst = 32'hc4050a9;
      6953: inst = 32'h8220000;
      6954: inst = 32'h10408000;
      6955: inst = 32'hc4050aa;
      6956: inst = 32'h8220000;
      6957: inst = 32'h10408000;
      6958: inst = 32'hc4050ab;
      6959: inst = 32'h8220000;
      6960: inst = 32'h10408000;
      6961: inst = 32'hc4050ac;
      6962: inst = 32'h8220000;
      6963: inst = 32'h10408000;
      6964: inst = 32'hc4050ad;
      6965: inst = 32'h8220000;
      6966: inst = 32'h10408000;
      6967: inst = 32'hc4050ae;
      6968: inst = 32'h8220000;
      6969: inst = 32'h10408000;
      6970: inst = 32'hc4050d7;
      6971: inst = 32'h8220000;
      6972: inst = 32'h10408000;
      6973: inst = 32'hc4050d8;
      6974: inst = 32'h8220000;
      6975: inst = 32'h10408000;
      6976: inst = 32'hc4050d9;
      6977: inst = 32'h8220000;
      6978: inst = 32'h10408000;
      6979: inst = 32'hc4050da;
      6980: inst = 32'h8220000;
      6981: inst = 32'h10408000;
      6982: inst = 32'hc4050db;
      6983: inst = 32'h8220000;
      6984: inst = 32'h10408000;
      6985: inst = 32'hc4050dc;
      6986: inst = 32'h8220000;
      6987: inst = 32'h10408000;
      6988: inst = 32'hc4050dd;
      6989: inst = 32'h8220000;
      6990: inst = 32'h10408000;
      6991: inst = 32'hc4050de;
      6992: inst = 32'h8220000;
      6993: inst = 32'h10408000;
      6994: inst = 32'hc4050e8;
      6995: inst = 32'h8220000;
      6996: inst = 32'h10408000;
      6997: inst = 32'hc4050e9;
      6998: inst = 32'h8220000;
      6999: inst = 32'h10408000;
      7000: inst = 32'hc4050ea;
      7001: inst = 32'h8220000;
      7002: inst = 32'h10408000;
      7003: inst = 32'hc4050eb;
      7004: inst = 32'h8220000;
      7005: inst = 32'h10408000;
      7006: inst = 32'hc4050ec;
      7007: inst = 32'h8220000;
      7008: inst = 32'h10408000;
      7009: inst = 32'hc4050ed;
      7010: inst = 32'h8220000;
      7011: inst = 32'h10408000;
      7012: inst = 32'hc4050ee;
      7013: inst = 32'h8220000;
      7014: inst = 32'h10408000;
      7015: inst = 32'hc4050ef;
      7016: inst = 32'h8220000;
      7017: inst = 32'h10408000;
      7018: inst = 32'hc4050f0;
      7019: inst = 32'h8220000;
      7020: inst = 32'h10408000;
      7021: inst = 32'hc4050f1;
      7022: inst = 32'h8220000;
      7023: inst = 32'h10408000;
      7024: inst = 32'hc4050f2;
      7025: inst = 32'h8220000;
      7026: inst = 32'h10408000;
      7027: inst = 32'hc4050f3;
      7028: inst = 32'h8220000;
      7029: inst = 32'h10408000;
      7030: inst = 32'hc4050f4;
      7031: inst = 32'h8220000;
      7032: inst = 32'h10408000;
      7033: inst = 32'hc4050f5;
      7034: inst = 32'h8220000;
      7035: inst = 32'h10408000;
      7036: inst = 32'hc4050f6;
      7037: inst = 32'h8220000;
      7038: inst = 32'h10408000;
      7039: inst = 32'hc4050f7;
      7040: inst = 32'h8220000;
      7041: inst = 32'h10408000;
      7042: inst = 32'hc405101;
      7043: inst = 32'h8220000;
      7044: inst = 32'h10408000;
      7045: inst = 32'hc405102;
      7046: inst = 32'h8220000;
      7047: inst = 32'h10408000;
      7048: inst = 32'hc405103;
      7049: inst = 32'h8220000;
      7050: inst = 32'h10408000;
      7051: inst = 32'hc405104;
      7052: inst = 32'h8220000;
      7053: inst = 32'h10408000;
      7054: inst = 32'hc405105;
      7055: inst = 32'h8220000;
      7056: inst = 32'h10408000;
      7057: inst = 32'hc405106;
      7058: inst = 32'h8220000;
      7059: inst = 32'h10408000;
      7060: inst = 32'hc405107;
      7061: inst = 32'h8220000;
      7062: inst = 32'h10408000;
      7063: inst = 32'hc405108;
      7064: inst = 32'h8220000;
      7065: inst = 32'h10408000;
      7066: inst = 32'hc405109;
      7067: inst = 32'h8220000;
      7068: inst = 32'h10408000;
      7069: inst = 32'hc40510a;
      7070: inst = 32'h8220000;
      7071: inst = 32'h10408000;
      7072: inst = 32'hc40510b;
      7073: inst = 32'h8220000;
      7074: inst = 32'h10408000;
      7075: inst = 32'hc40510c;
      7076: inst = 32'h8220000;
      7077: inst = 32'h10408000;
      7078: inst = 32'hc40510d;
      7079: inst = 32'h8220000;
      7080: inst = 32'h10408000;
      7081: inst = 32'hc40510e;
      7082: inst = 32'h8220000;
      7083: inst = 32'h10408000;
      7084: inst = 32'hc405137;
      7085: inst = 32'h8220000;
      7086: inst = 32'h10408000;
      7087: inst = 32'hc405138;
      7088: inst = 32'h8220000;
      7089: inst = 32'h10408000;
      7090: inst = 32'hc405139;
      7091: inst = 32'h8220000;
      7092: inst = 32'h10408000;
      7093: inst = 32'hc40513a;
      7094: inst = 32'h8220000;
      7095: inst = 32'h10408000;
      7096: inst = 32'hc40513b;
      7097: inst = 32'h8220000;
      7098: inst = 32'h10408000;
      7099: inst = 32'hc40513c;
      7100: inst = 32'h8220000;
      7101: inst = 32'h10408000;
      7102: inst = 32'hc40513d;
      7103: inst = 32'h8220000;
      7104: inst = 32'h10408000;
      7105: inst = 32'hc40513e;
      7106: inst = 32'h8220000;
      7107: inst = 32'h10408000;
      7108: inst = 32'hc405148;
      7109: inst = 32'h8220000;
      7110: inst = 32'h10408000;
      7111: inst = 32'hc405149;
      7112: inst = 32'h8220000;
      7113: inst = 32'h10408000;
      7114: inst = 32'hc40514a;
      7115: inst = 32'h8220000;
      7116: inst = 32'h10408000;
      7117: inst = 32'hc40514b;
      7118: inst = 32'h8220000;
      7119: inst = 32'h10408000;
      7120: inst = 32'hc40514c;
      7121: inst = 32'h8220000;
      7122: inst = 32'h10408000;
      7123: inst = 32'hc40514d;
      7124: inst = 32'h8220000;
      7125: inst = 32'h10408000;
      7126: inst = 32'hc40514e;
      7127: inst = 32'h8220000;
      7128: inst = 32'h10408000;
      7129: inst = 32'hc40514f;
      7130: inst = 32'h8220000;
      7131: inst = 32'h10408000;
      7132: inst = 32'hc405150;
      7133: inst = 32'h8220000;
      7134: inst = 32'h10408000;
      7135: inst = 32'hc405151;
      7136: inst = 32'h8220000;
      7137: inst = 32'h10408000;
      7138: inst = 32'hc405152;
      7139: inst = 32'h8220000;
      7140: inst = 32'h10408000;
      7141: inst = 32'hc405153;
      7142: inst = 32'h8220000;
      7143: inst = 32'h10408000;
      7144: inst = 32'hc405154;
      7145: inst = 32'h8220000;
      7146: inst = 32'h10408000;
      7147: inst = 32'hc405155;
      7148: inst = 32'h8220000;
      7149: inst = 32'h10408000;
      7150: inst = 32'hc405156;
      7151: inst = 32'h8220000;
      7152: inst = 32'h10408000;
      7153: inst = 32'hc405157;
      7154: inst = 32'h8220000;
      7155: inst = 32'h10408000;
      7156: inst = 32'hc405161;
      7157: inst = 32'h8220000;
      7158: inst = 32'h10408000;
      7159: inst = 32'hc405162;
      7160: inst = 32'h8220000;
      7161: inst = 32'h10408000;
      7162: inst = 32'hc405163;
      7163: inst = 32'h8220000;
      7164: inst = 32'h10408000;
      7165: inst = 32'hc405164;
      7166: inst = 32'h8220000;
      7167: inst = 32'h10408000;
      7168: inst = 32'hc405165;
      7169: inst = 32'h8220000;
      7170: inst = 32'h10408000;
      7171: inst = 32'hc405166;
      7172: inst = 32'h8220000;
      7173: inst = 32'h10408000;
      7174: inst = 32'hc405167;
      7175: inst = 32'h8220000;
      7176: inst = 32'h10408000;
      7177: inst = 32'hc405168;
      7178: inst = 32'h8220000;
      7179: inst = 32'h10408000;
      7180: inst = 32'hc405169;
      7181: inst = 32'h8220000;
      7182: inst = 32'h10408000;
      7183: inst = 32'hc40516a;
      7184: inst = 32'h8220000;
      7185: inst = 32'h10408000;
      7186: inst = 32'hc40516b;
      7187: inst = 32'h8220000;
      7188: inst = 32'h10408000;
      7189: inst = 32'hc40516c;
      7190: inst = 32'h8220000;
      7191: inst = 32'h10408000;
      7192: inst = 32'hc40516d;
      7193: inst = 32'h8220000;
      7194: inst = 32'h10408000;
      7195: inst = 32'hc40516e;
      7196: inst = 32'h8220000;
      7197: inst = 32'h10408000;
      7198: inst = 32'hc405197;
      7199: inst = 32'h8220000;
      7200: inst = 32'h10408000;
      7201: inst = 32'hc405198;
      7202: inst = 32'h8220000;
      7203: inst = 32'h10408000;
      7204: inst = 32'hc405199;
      7205: inst = 32'h8220000;
      7206: inst = 32'h10408000;
      7207: inst = 32'hc40519a;
      7208: inst = 32'h8220000;
      7209: inst = 32'h10408000;
      7210: inst = 32'hc40519b;
      7211: inst = 32'h8220000;
      7212: inst = 32'h10408000;
      7213: inst = 32'hc40519c;
      7214: inst = 32'h8220000;
      7215: inst = 32'h10408000;
      7216: inst = 32'hc40519d;
      7217: inst = 32'h8220000;
      7218: inst = 32'h10408000;
      7219: inst = 32'hc4051aa;
      7220: inst = 32'h8220000;
      7221: inst = 32'h10408000;
      7222: inst = 32'hc4051ab;
      7223: inst = 32'h8220000;
      7224: inst = 32'h10408000;
      7225: inst = 32'hc4051ac;
      7226: inst = 32'h8220000;
      7227: inst = 32'h10408000;
      7228: inst = 32'hc4051ad;
      7229: inst = 32'h8220000;
      7230: inst = 32'h10408000;
      7231: inst = 32'hc4051ae;
      7232: inst = 32'h8220000;
      7233: inst = 32'h10408000;
      7234: inst = 32'hc4051af;
      7235: inst = 32'h8220000;
      7236: inst = 32'h10408000;
      7237: inst = 32'hc4051b0;
      7238: inst = 32'h8220000;
      7239: inst = 32'h10408000;
      7240: inst = 32'hc4051b1;
      7241: inst = 32'h8220000;
      7242: inst = 32'h10408000;
      7243: inst = 32'hc4051b2;
      7244: inst = 32'h8220000;
      7245: inst = 32'h10408000;
      7246: inst = 32'hc4051b3;
      7247: inst = 32'h8220000;
      7248: inst = 32'h10408000;
      7249: inst = 32'hc4051b4;
      7250: inst = 32'h8220000;
      7251: inst = 32'h10408000;
      7252: inst = 32'hc4051b5;
      7253: inst = 32'h8220000;
      7254: inst = 32'h10408000;
      7255: inst = 32'hc4051c2;
      7256: inst = 32'h8220000;
      7257: inst = 32'h10408000;
      7258: inst = 32'hc4051c3;
      7259: inst = 32'h8220000;
      7260: inst = 32'h10408000;
      7261: inst = 32'hc4051c4;
      7262: inst = 32'h8220000;
      7263: inst = 32'h10408000;
      7264: inst = 32'hc4051c5;
      7265: inst = 32'h8220000;
      7266: inst = 32'h10408000;
      7267: inst = 32'hc4051c6;
      7268: inst = 32'h8220000;
      7269: inst = 32'h10408000;
      7270: inst = 32'hc4051c7;
      7271: inst = 32'h8220000;
      7272: inst = 32'h10408000;
      7273: inst = 32'hc4051c8;
      7274: inst = 32'h8220000;
      7275: inst = 32'h10408000;
      7276: inst = 32'hc4051c9;
      7277: inst = 32'h8220000;
      7278: inst = 32'h10408000;
      7279: inst = 32'hc4051ca;
      7280: inst = 32'h8220000;
      7281: inst = 32'h10408000;
      7282: inst = 32'hc4051cb;
      7283: inst = 32'h8220000;
      7284: inst = 32'h10408000;
      7285: inst = 32'hc4051cc;
      7286: inst = 32'h8220000;
      7287: inst = 32'h10408000;
      7288: inst = 32'hc4051cd;
      7289: inst = 32'h8220000;
      7290: inst = 32'h10408000;
      7291: inst = 32'hc4051ce;
      7292: inst = 32'h8220000;
      7293: inst = 32'h10408000;
      7294: inst = 32'hc4051f7;
      7295: inst = 32'h8220000;
      7296: inst = 32'h10408000;
      7297: inst = 32'hc4051f8;
      7298: inst = 32'h8220000;
      7299: inst = 32'h10408000;
      7300: inst = 32'hc4051f9;
      7301: inst = 32'h8220000;
      7302: inst = 32'h10408000;
      7303: inst = 32'hc4051fa;
      7304: inst = 32'h8220000;
      7305: inst = 32'h10408000;
      7306: inst = 32'hc4051fb;
      7307: inst = 32'h8220000;
      7308: inst = 32'h10408000;
      7309: inst = 32'hc4051fc;
      7310: inst = 32'h8220000;
      7311: inst = 32'h10408000;
      7312: inst = 32'hc40520a;
      7313: inst = 32'h8220000;
      7314: inst = 32'h10408000;
      7315: inst = 32'hc40520b;
      7316: inst = 32'h8220000;
      7317: inst = 32'h10408000;
      7318: inst = 32'hc40520c;
      7319: inst = 32'h8220000;
      7320: inst = 32'h10408000;
      7321: inst = 32'hc40520d;
      7322: inst = 32'h8220000;
      7323: inst = 32'h10408000;
      7324: inst = 32'hc40520e;
      7325: inst = 32'h8220000;
      7326: inst = 32'h10408000;
      7327: inst = 32'hc40520f;
      7328: inst = 32'h8220000;
      7329: inst = 32'h10408000;
      7330: inst = 32'hc405210;
      7331: inst = 32'h8220000;
      7332: inst = 32'h10408000;
      7333: inst = 32'hc405211;
      7334: inst = 32'h8220000;
      7335: inst = 32'h10408000;
      7336: inst = 32'hc405212;
      7337: inst = 32'h8220000;
      7338: inst = 32'h10408000;
      7339: inst = 32'hc405213;
      7340: inst = 32'h8220000;
      7341: inst = 32'h10408000;
      7342: inst = 32'hc405214;
      7343: inst = 32'h8220000;
      7344: inst = 32'h10408000;
      7345: inst = 32'hc405215;
      7346: inst = 32'h8220000;
      7347: inst = 32'h10408000;
      7348: inst = 32'hc405223;
      7349: inst = 32'h8220000;
      7350: inst = 32'h10408000;
      7351: inst = 32'hc405224;
      7352: inst = 32'h8220000;
      7353: inst = 32'h10408000;
      7354: inst = 32'hc405225;
      7355: inst = 32'h8220000;
      7356: inst = 32'h10408000;
      7357: inst = 32'hc405226;
      7358: inst = 32'h8220000;
      7359: inst = 32'h10408000;
      7360: inst = 32'hc405227;
      7361: inst = 32'h8220000;
      7362: inst = 32'h10408000;
      7363: inst = 32'hc405228;
      7364: inst = 32'h8220000;
      7365: inst = 32'h10408000;
      7366: inst = 32'hc405229;
      7367: inst = 32'h8220000;
      7368: inst = 32'h10408000;
      7369: inst = 32'hc40522a;
      7370: inst = 32'h8220000;
      7371: inst = 32'h10408000;
      7372: inst = 32'hc40522b;
      7373: inst = 32'h8220000;
      7374: inst = 32'h10408000;
      7375: inst = 32'hc40522c;
      7376: inst = 32'h8220000;
      7377: inst = 32'h10408000;
      7378: inst = 32'hc40522d;
      7379: inst = 32'h8220000;
      7380: inst = 32'h10408000;
      7381: inst = 32'hc40522e;
      7382: inst = 32'h8220000;
      7383: inst = 32'h10408000;
      7384: inst = 32'hc405257;
      7385: inst = 32'h8220000;
      7386: inst = 32'h10408000;
      7387: inst = 32'hc405258;
      7388: inst = 32'h8220000;
      7389: inst = 32'h10408000;
      7390: inst = 32'hc405259;
      7391: inst = 32'h8220000;
      7392: inst = 32'h10408000;
      7393: inst = 32'hc40525a;
      7394: inst = 32'h8220000;
      7395: inst = 32'h10408000;
      7396: inst = 32'hc40525b;
      7397: inst = 32'h8220000;
      7398: inst = 32'h10408000;
      7399: inst = 32'hc40526a;
      7400: inst = 32'h8220000;
      7401: inst = 32'h10408000;
      7402: inst = 32'hc40526b;
      7403: inst = 32'h8220000;
      7404: inst = 32'h10408000;
      7405: inst = 32'hc40526c;
      7406: inst = 32'h8220000;
      7407: inst = 32'h10408000;
      7408: inst = 32'hc40526d;
      7409: inst = 32'h8220000;
      7410: inst = 32'h10408000;
      7411: inst = 32'hc40526e;
      7412: inst = 32'h8220000;
      7413: inst = 32'h10408000;
      7414: inst = 32'hc40526f;
      7415: inst = 32'h8220000;
      7416: inst = 32'h10408000;
      7417: inst = 32'hc405270;
      7418: inst = 32'h8220000;
      7419: inst = 32'h10408000;
      7420: inst = 32'hc405271;
      7421: inst = 32'h8220000;
      7422: inst = 32'h10408000;
      7423: inst = 32'hc405272;
      7424: inst = 32'h8220000;
      7425: inst = 32'h10408000;
      7426: inst = 32'hc405273;
      7427: inst = 32'h8220000;
      7428: inst = 32'h10408000;
      7429: inst = 32'hc405274;
      7430: inst = 32'h8220000;
      7431: inst = 32'h10408000;
      7432: inst = 32'hc405275;
      7433: inst = 32'h8220000;
      7434: inst = 32'h10408000;
      7435: inst = 32'hc405284;
      7436: inst = 32'h8220000;
      7437: inst = 32'h10408000;
      7438: inst = 32'hc405285;
      7439: inst = 32'h8220000;
      7440: inst = 32'h10408000;
      7441: inst = 32'hc405286;
      7442: inst = 32'h8220000;
      7443: inst = 32'h10408000;
      7444: inst = 32'hc405287;
      7445: inst = 32'h8220000;
      7446: inst = 32'h10408000;
      7447: inst = 32'hc405288;
      7448: inst = 32'h8220000;
      7449: inst = 32'h10408000;
      7450: inst = 32'hc405289;
      7451: inst = 32'h8220000;
      7452: inst = 32'h10408000;
      7453: inst = 32'hc40528a;
      7454: inst = 32'h8220000;
      7455: inst = 32'h10408000;
      7456: inst = 32'hc40528b;
      7457: inst = 32'h8220000;
      7458: inst = 32'h10408000;
      7459: inst = 32'hc40528c;
      7460: inst = 32'h8220000;
      7461: inst = 32'h10408000;
      7462: inst = 32'hc40528d;
      7463: inst = 32'h8220000;
      7464: inst = 32'h10408000;
      7465: inst = 32'hc40528e;
      7466: inst = 32'h8220000;
      7467: inst = 32'h10408000;
      7468: inst = 32'hc4052b7;
      7469: inst = 32'h8220000;
      7470: inst = 32'h10408000;
      7471: inst = 32'hc4052b8;
      7472: inst = 32'h8220000;
      7473: inst = 32'h10408000;
      7474: inst = 32'hc4052b9;
      7475: inst = 32'h8220000;
      7476: inst = 32'h10408000;
      7477: inst = 32'hc4052ba;
      7478: inst = 32'h8220000;
      7479: inst = 32'h10408000;
      7480: inst = 32'hc4052bb;
      7481: inst = 32'h8220000;
      7482: inst = 32'h10408000;
      7483: inst = 32'hc4052ca;
      7484: inst = 32'h8220000;
      7485: inst = 32'h10408000;
      7486: inst = 32'hc4052cb;
      7487: inst = 32'h8220000;
      7488: inst = 32'h10408000;
      7489: inst = 32'hc4052cc;
      7490: inst = 32'h8220000;
      7491: inst = 32'h10408000;
      7492: inst = 32'hc4052cd;
      7493: inst = 32'h8220000;
      7494: inst = 32'h10408000;
      7495: inst = 32'hc4052ce;
      7496: inst = 32'h8220000;
      7497: inst = 32'h10408000;
      7498: inst = 32'hc4052cf;
      7499: inst = 32'h8220000;
      7500: inst = 32'h10408000;
      7501: inst = 32'hc4052d0;
      7502: inst = 32'h8220000;
      7503: inst = 32'h10408000;
      7504: inst = 32'hc4052d1;
      7505: inst = 32'h8220000;
      7506: inst = 32'h10408000;
      7507: inst = 32'hc4052d2;
      7508: inst = 32'h8220000;
      7509: inst = 32'h10408000;
      7510: inst = 32'hc4052d3;
      7511: inst = 32'h8220000;
      7512: inst = 32'h10408000;
      7513: inst = 32'hc4052d4;
      7514: inst = 32'h8220000;
      7515: inst = 32'h10408000;
      7516: inst = 32'hc4052d5;
      7517: inst = 32'h8220000;
      7518: inst = 32'h10408000;
      7519: inst = 32'hc4052e4;
      7520: inst = 32'h8220000;
      7521: inst = 32'h10408000;
      7522: inst = 32'hc4052e5;
      7523: inst = 32'h8220000;
      7524: inst = 32'h10408000;
      7525: inst = 32'hc4052e6;
      7526: inst = 32'h8220000;
      7527: inst = 32'h10408000;
      7528: inst = 32'hc4052e7;
      7529: inst = 32'h8220000;
      7530: inst = 32'h10408000;
      7531: inst = 32'hc4052e8;
      7532: inst = 32'h8220000;
      7533: inst = 32'h10408000;
      7534: inst = 32'hc4052e9;
      7535: inst = 32'h8220000;
      7536: inst = 32'h10408000;
      7537: inst = 32'hc4052ea;
      7538: inst = 32'h8220000;
      7539: inst = 32'h10408000;
      7540: inst = 32'hc4052eb;
      7541: inst = 32'h8220000;
      7542: inst = 32'h10408000;
      7543: inst = 32'hc4052ec;
      7544: inst = 32'h8220000;
      7545: inst = 32'h10408000;
      7546: inst = 32'hc4052ed;
      7547: inst = 32'h8220000;
      7548: inst = 32'h10408000;
      7549: inst = 32'hc4052ee;
      7550: inst = 32'h8220000;
      7551: inst = 32'hc2094b2;
      7552: inst = 32'h10408000;
      7553: inst = 32'hc403feb;
      7554: inst = 32'h8220000;
      7555: inst = 32'h10408000;
      7556: inst = 32'hc40404b;
      7557: inst = 32'h8220000;
      7558: inst = 32'h10408000;
      7559: inst = 32'hc4040ab;
      7560: inst = 32'h8220000;
      7561: inst = 32'h10408000;
      7562: inst = 32'hc40410b;
      7563: inst = 32'h8220000;
      7564: inst = 32'h10408000;
      7565: inst = 32'hc40416b;
      7566: inst = 32'h8220000;
      7567: inst = 32'h10408000;
      7568: inst = 32'hc4041cb;
      7569: inst = 32'h8220000;
      7570: inst = 32'h10408000;
      7571: inst = 32'hc40422b;
      7572: inst = 32'h8220000;
      7573: inst = 32'h10408000;
      7574: inst = 32'hc40428b;
      7575: inst = 32'h8220000;
      7576: inst = 32'hc20b596;
      7577: inst = 32'h10408000;
      7578: inst = 32'hc4041da;
      7579: inst = 32'h8220000;
      7580: inst = 32'h10408000;
      7581: inst = 32'hc4041db;
      7582: inst = 32'h8220000;
      7583: inst = 32'h10408000;
      7584: inst = 32'hc4041dc;
      7585: inst = 32'h8220000;
      7586: inst = 32'h10408000;
      7587: inst = 32'hc4041dd;
      7588: inst = 32'h8220000;
      7589: inst = 32'h10408000;
      7590: inst = 32'hc4041de;
      7591: inst = 32'h8220000;
      7592: inst = 32'h10408000;
      7593: inst = 32'hc4041df;
      7594: inst = 32'h8220000;
      7595: inst = 32'h10408000;
      7596: inst = 32'hc4041e0;
      7597: inst = 32'h8220000;
      7598: inst = 32'h10408000;
      7599: inst = 32'hc4041e1;
      7600: inst = 32'h8220000;
      7601: inst = 32'h10408000;
      7602: inst = 32'hc4041e2;
      7603: inst = 32'h8220000;
      7604: inst = 32'h10408000;
      7605: inst = 32'hc4041e3;
      7606: inst = 32'h8220000;
      7607: inst = 32'h10408000;
      7608: inst = 32'hc4041e4;
      7609: inst = 32'h8220000;
      7610: inst = 32'h10408000;
      7611: inst = 32'hc4041e5;
      7612: inst = 32'h8220000;
      7613: inst = 32'h10408000;
      7614: inst = 32'hc4041e6;
      7615: inst = 32'h8220000;
      7616: inst = 32'h10408000;
      7617: inst = 32'hc4041e7;
      7618: inst = 32'h8220000;
      7619: inst = 32'h10408000;
      7620: inst = 32'hc4041e8;
      7621: inst = 32'h8220000;
      7622: inst = 32'h10408000;
      7623: inst = 32'hc4041e9;
      7624: inst = 32'h8220000;
      7625: inst = 32'h10408000;
      7626: inst = 32'hc4041ea;
      7627: inst = 32'h8220000;
      7628: inst = 32'h10408000;
      7629: inst = 32'hc4041eb;
      7630: inst = 32'h8220000;
      7631: inst = 32'h10408000;
      7632: inst = 32'hc4041ec;
      7633: inst = 32'h8220000;
      7634: inst = 32'h10408000;
      7635: inst = 32'hc4041ed;
      7636: inst = 32'h8220000;
      7637: inst = 32'h10408000;
      7638: inst = 32'hc4041ee;
      7639: inst = 32'h8220000;
      7640: inst = 32'h10408000;
      7641: inst = 32'hc4041ef;
      7642: inst = 32'h8220000;
      7643: inst = 32'h10408000;
      7644: inst = 32'hc4041f0;
      7645: inst = 32'h8220000;
      7646: inst = 32'h10408000;
      7647: inst = 32'hc4041f1;
      7648: inst = 32'h8220000;
      7649: inst = 32'h10408000;
      7650: inst = 32'hc4041f2;
      7651: inst = 32'h8220000;
      7652: inst = 32'h10408000;
      7653: inst = 32'hc4041f3;
      7654: inst = 32'h8220000;
      7655: inst = 32'h10408000;
      7656: inst = 32'hc4041f4;
      7657: inst = 32'h8220000;
      7658: inst = 32'h10408000;
      7659: inst = 32'hc4041f5;
      7660: inst = 32'h8220000;
      7661: inst = 32'h10408000;
      7662: inst = 32'hc4041f6;
      7663: inst = 32'h8220000;
      7664: inst = 32'h10408000;
      7665: inst = 32'hc4041f7;
      7666: inst = 32'h8220000;
      7667: inst = 32'h10408000;
      7668: inst = 32'hc4041f8;
      7669: inst = 32'h8220000;
      7670: inst = 32'h10408000;
      7671: inst = 32'hc4041f9;
      7672: inst = 32'h8220000;
      7673: inst = 32'h10408000;
      7674: inst = 32'hc4041fa;
      7675: inst = 32'h8220000;
      7676: inst = 32'h10408000;
      7677: inst = 32'hc4041fb;
      7678: inst = 32'h8220000;
      7679: inst = 32'h10408000;
      7680: inst = 32'hc4041fc;
      7681: inst = 32'h8220000;
      7682: inst = 32'h10408000;
      7683: inst = 32'hc4041fd;
      7684: inst = 32'h8220000;
      7685: inst = 32'h10408000;
      7686: inst = 32'hc4041fe;
      7687: inst = 32'h8220000;
      7688: inst = 32'h10408000;
      7689: inst = 32'hc4041ff;
      7690: inst = 32'h8220000;
      7691: inst = 32'h10408000;
      7692: inst = 32'hc404200;
      7693: inst = 32'h8220000;
      7694: inst = 32'h10408000;
      7695: inst = 32'hc404201;
      7696: inst = 32'h8220000;
      7697: inst = 32'h10408000;
      7698: inst = 32'hc404202;
      7699: inst = 32'h8220000;
      7700: inst = 32'h10408000;
      7701: inst = 32'hc404203;
      7702: inst = 32'h8220000;
      7703: inst = 32'h10408000;
      7704: inst = 32'hc404204;
      7705: inst = 32'h8220000;
      7706: inst = 32'h10408000;
      7707: inst = 32'hc404205;
      7708: inst = 32'h8220000;
      7709: inst = 32'h10408000;
      7710: inst = 32'hc404bfa;
      7711: inst = 32'h8220000;
      7712: inst = 32'h10408000;
      7713: inst = 32'hc404bfb;
      7714: inst = 32'h8220000;
      7715: inst = 32'h10408000;
      7716: inst = 32'hc404bfc;
      7717: inst = 32'h8220000;
      7718: inst = 32'h10408000;
      7719: inst = 32'hc404bfd;
      7720: inst = 32'h8220000;
      7721: inst = 32'h10408000;
      7722: inst = 32'hc404bfe;
      7723: inst = 32'h8220000;
      7724: inst = 32'h10408000;
      7725: inst = 32'hc404bff;
      7726: inst = 32'h8220000;
      7727: inst = 32'h10408000;
      7728: inst = 32'hc404c00;
      7729: inst = 32'h8220000;
      7730: inst = 32'h10408000;
      7731: inst = 32'hc404c01;
      7732: inst = 32'h8220000;
      7733: inst = 32'h10408000;
      7734: inst = 32'hc404c02;
      7735: inst = 32'h8220000;
      7736: inst = 32'h10408000;
      7737: inst = 32'hc404c03;
      7738: inst = 32'h8220000;
      7739: inst = 32'h10408000;
      7740: inst = 32'hc404c04;
      7741: inst = 32'h8220000;
      7742: inst = 32'h10408000;
      7743: inst = 32'hc404c05;
      7744: inst = 32'h8220000;
      7745: inst = 32'h10408000;
      7746: inst = 32'hc404c06;
      7747: inst = 32'h8220000;
      7748: inst = 32'h10408000;
      7749: inst = 32'hc404c07;
      7750: inst = 32'h8220000;
      7751: inst = 32'h10408000;
      7752: inst = 32'hc404c08;
      7753: inst = 32'h8220000;
      7754: inst = 32'h10408000;
      7755: inst = 32'hc404c09;
      7756: inst = 32'h8220000;
      7757: inst = 32'h10408000;
      7758: inst = 32'hc404c0a;
      7759: inst = 32'h8220000;
      7760: inst = 32'h10408000;
      7761: inst = 32'hc404c0b;
      7762: inst = 32'h8220000;
      7763: inst = 32'h10408000;
      7764: inst = 32'hc404c0c;
      7765: inst = 32'h8220000;
      7766: inst = 32'h10408000;
      7767: inst = 32'hc404c0d;
      7768: inst = 32'h8220000;
      7769: inst = 32'h10408000;
      7770: inst = 32'hc404c0e;
      7771: inst = 32'h8220000;
      7772: inst = 32'h10408000;
      7773: inst = 32'hc404c0f;
      7774: inst = 32'h8220000;
      7775: inst = 32'h10408000;
      7776: inst = 32'hc404c10;
      7777: inst = 32'h8220000;
      7778: inst = 32'h10408000;
      7779: inst = 32'hc404c11;
      7780: inst = 32'h8220000;
      7781: inst = 32'h10408000;
      7782: inst = 32'hc404c12;
      7783: inst = 32'h8220000;
      7784: inst = 32'h10408000;
      7785: inst = 32'hc404c13;
      7786: inst = 32'h8220000;
      7787: inst = 32'h10408000;
      7788: inst = 32'hc404c14;
      7789: inst = 32'h8220000;
      7790: inst = 32'h10408000;
      7791: inst = 32'hc404c15;
      7792: inst = 32'h8220000;
      7793: inst = 32'h10408000;
      7794: inst = 32'hc404c16;
      7795: inst = 32'h8220000;
      7796: inst = 32'h10408000;
      7797: inst = 32'hc404c17;
      7798: inst = 32'h8220000;
      7799: inst = 32'h10408000;
      7800: inst = 32'hc404c18;
      7801: inst = 32'h8220000;
      7802: inst = 32'h10408000;
      7803: inst = 32'hc404c19;
      7804: inst = 32'h8220000;
      7805: inst = 32'h10408000;
      7806: inst = 32'hc404c1a;
      7807: inst = 32'h8220000;
      7808: inst = 32'h10408000;
      7809: inst = 32'hc404c1b;
      7810: inst = 32'h8220000;
      7811: inst = 32'h10408000;
      7812: inst = 32'hc404c1c;
      7813: inst = 32'h8220000;
      7814: inst = 32'h10408000;
      7815: inst = 32'hc404c1d;
      7816: inst = 32'h8220000;
      7817: inst = 32'h10408000;
      7818: inst = 32'hc404c1e;
      7819: inst = 32'h8220000;
      7820: inst = 32'h10408000;
      7821: inst = 32'hc404c1f;
      7822: inst = 32'h8220000;
      7823: inst = 32'h10408000;
      7824: inst = 32'hc404c20;
      7825: inst = 32'h8220000;
      7826: inst = 32'h10408000;
      7827: inst = 32'hc404c21;
      7828: inst = 32'h8220000;
      7829: inst = 32'h10408000;
      7830: inst = 32'hc404c22;
      7831: inst = 32'h8220000;
      7832: inst = 32'h10408000;
      7833: inst = 32'hc404c23;
      7834: inst = 32'h8220000;
      7835: inst = 32'h10408000;
      7836: inst = 32'hc404c24;
      7837: inst = 32'h8220000;
      7838: inst = 32'h10408000;
      7839: inst = 32'hc404c25;
      7840: inst = 32'h8220000;
      7841: inst = 32'hc20ffff;
      7842: inst = 32'h10408000;
      7843: inst = 32'hc40423c;
      7844: inst = 32'h8220000;
      7845: inst = 32'h10408000;
      7846: inst = 32'hc40423d;
      7847: inst = 32'h8220000;
      7848: inst = 32'h10408000;
      7849: inst = 32'hc40423e;
      7850: inst = 32'h8220000;
      7851: inst = 32'h10408000;
      7852: inst = 32'hc40423f;
      7853: inst = 32'h8220000;
      7854: inst = 32'h10408000;
      7855: inst = 32'hc404240;
      7856: inst = 32'h8220000;
      7857: inst = 32'h10408000;
      7858: inst = 32'hc404241;
      7859: inst = 32'h8220000;
      7860: inst = 32'h10408000;
      7861: inst = 32'hc404242;
      7862: inst = 32'h8220000;
      7863: inst = 32'h10408000;
      7864: inst = 32'hc404243;
      7865: inst = 32'h8220000;
      7866: inst = 32'h10408000;
      7867: inst = 32'hc404244;
      7868: inst = 32'h8220000;
      7869: inst = 32'h10408000;
      7870: inst = 32'hc404245;
      7871: inst = 32'h8220000;
      7872: inst = 32'h10408000;
      7873: inst = 32'hc404246;
      7874: inst = 32'h8220000;
      7875: inst = 32'h10408000;
      7876: inst = 32'hc404247;
      7877: inst = 32'h8220000;
      7878: inst = 32'h10408000;
      7879: inst = 32'hc404248;
      7880: inst = 32'h8220000;
      7881: inst = 32'h10408000;
      7882: inst = 32'hc404249;
      7883: inst = 32'h8220000;
      7884: inst = 32'h10408000;
      7885: inst = 32'hc40424a;
      7886: inst = 32'h8220000;
      7887: inst = 32'h10408000;
      7888: inst = 32'hc40424b;
      7889: inst = 32'h8220000;
      7890: inst = 32'h10408000;
      7891: inst = 32'hc40424c;
      7892: inst = 32'h8220000;
      7893: inst = 32'h10408000;
      7894: inst = 32'hc40424d;
      7895: inst = 32'h8220000;
      7896: inst = 32'h10408000;
      7897: inst = 32'hc40424e;
      7898: inst = 32'h8220000;
      7899: inst = 32'h10408000;
      7900: inst = 32'hc40424f;
      7901: inst = 32'h8220000;
      7902: inst = 32'h10408000;
      7903: inst = 32'hc404250;
      7904: inst = 32'h8220000;
      7905: inst = 32'h10408000;
      7906: inst = 32'hc404251;
      7907: inst = 32'h8220000;
      7908: inst = 32'h10408000;
      7909: inst = 32'hc404252;
      7910: inst = 32'h8220000;
      7911: inst = 32'h10408000;
      7912: inst = 32'hc404253;
      7913: inst = 32'h8220000;
      7914: inst = 32'h10408000;
      7915: inst = 32'hc404254;
      7916: inst = 32'h8220000;
      7917: inst = 32'h10408000;
      7918: inst = 32'hc404255;
      7919: inst = 32'h8220000;
      7920: inst = 32'h10408000;
      7921: inst = 32'hc404256;
      7922: inst = 32'h8220000;
      7923: inst = 32'h10408000;
      7924: inst = 32'hc404257;
      7925: inst = 32'h8220000;
      7926: inst = 32'h10408000;
      7927: inst = 32'hc404258;
      7928: inst = 32'h8220000;
      7929: inst = 32'h10408000;
      7930: inst = 32'hc404259;
      7931: inst = 32'h8220000;
      7932: inst = 32'h10408000;
      7933: inst = 32'hc40425a;
      7934: inst = 32'h8220000;
      7935: inst = 32'h10408000;
      7936: inst = 32'hc40425b;
      7937: inst = 32'h8220000;
      7938: inst = 32'h10408000;
      7939: inst = 32'hc40425c;
      7940: inst = 32'h8220000;
      7941: inst = 32'h10408000;
      7942: inst = 32'hc40425d;
      7943: inst = 32'h8220000;
      7944: inst = 32'h10408000;
      7945: inst = 32'hc40425e;
      7946: inst = 32'h8220000;
      7947: inst = 32'h10408000;
      7948: inst = 32'hc40425f;
      7949: inst = 32'h8220000;
      7950: inst = 32'h10408000;
      7951: inst = 32'hc404260;
      7952: inst = 32'h8220000;
      7953: inst = 32'h10408000;
      7954: inst = 32'hc404261;
      7955: inst = 32'h8220000;
      7956: inst = 32'h10408000;
      7957: inst = 32'hc404262;
      7958: inst = 32'h8220000;
      7959: inst = 32'h10408000;
      7960: inst = 32'hc404263;
      7961: inst = 32'h8220000;
      7962: inst = 32'h10408000;
      7963: inst = 32'hc40429c;
      7964: inst = 32'h8220000;
      7965: inst = 32'h10408000;
      7966: inst = 32'hc40429d;
      7967: inst = 32'h8220000;
      7968: inst = 32'h10408000;
      7969: inst = 32'hc40429e;
      7970: inst = 32'h8220000;
      7971: inst = 32'h10408000;
      7972: inst = 32'hc40429f;
      7973: inst = 32'h8220000;
      7974: inst = 32'h10408000;
      7975: inst = 32'hc4042a0;
      7976: inst = 32'h8220000;
      7977: inst = 32'h10408000;
      7978: inst = 32'hc4042a1;
      7979: inst = 32'h8220000;
      7980: inst = 32'h10408000;
      7981: inst = 32'hc4042a2;
      7982: inst = 32'h8220000;
      7983: inst = 32'h10408000;
      7984: inst = 32'hc4042a3;
      7985: inst = 32'h8220000;
      7986: inst = 32'h10408000;
      7987: inst = 32'hc4042a4;
      7988: inst = 32'h8220000;
      7989: inst = 32'h10408000;
      7990: inst = 32'hc4042a5;
      7991: inst = 32'h8220000;
      7992: inst = 32'h10408000;
      7993: inst = 32'hc4042a6;
      7994: inst = 32'h8220000;
      7995: inst = 32'h10408000;
      7996: inst = 32'hc4042a7;
      7997: inst = 32'h8220000;
      7998: inst = 32'h10408000;
      7999: inst = 32'hc4042a8;
      8000: inst = 32'h8220000;
      8001: inst = 32'h10408000;
      8002: inst = 32'hc4042a9;
      8003: inst = 32'h8220000;
      8004: inst = 32'h10408000;
      8005: inst = 32'hc4042aa;
      8006: inst = 32'h8220000;
      8007: inst = 32'h10408000;
      8008: inst = 32'hc4042ab;
      8009: inst = 32'h8220000;
      8010: inst = 32'h10408000;
      8011: inst = 32'hc4042ac;
      8012: inst = 32'h8220000;
      8013: inst = 32'h10408000;
      8014: inst = 32'hc4042ad;
      8015: inst = 32'h8220000;
      8016: inst = 32'h10408000;
      8017: inst = 32'hc4042ae;
      8018: inst = 32'h8220000;
      8019: inst = 32'h10408000;
      8020: inst = 32'hc4042af;
      8021: inst = 32'h8220000;
      8022: inst = 32'h10408000;
      8023: inst = 32'hc4042b0;
      8024: inst = 32'h8220000;
      8025: inst = 32'h10408000;
      8026: inst = 32'hc4042b1;
      8027: inst = 32'h8220000;
      8028: inst = 32'h10408000;
      8029: inst = 32'hc4042b2;
      8030: inst = 32'h8220000;
      8031: inst = 32'h10408000;
      8032: inst = 32'hc4042b3;
      8033: inst = 32'h8220000;
      8034: inst = 32'h10408000;
      8035: inst = 32'hc4042b4;
      8036: inst = 32'h8220000;
      8037: inst = 32'h10408000;
      8038: inst = 32'hc4042b5;
      8039: inst = 32'h8220000;
      8040: inst = 32'h10408000;
      8041: inst = 32'hc4042b6;
      8042: inst = 32'h8220000;
      8043: inst = 32'h10408000;
      8044: inst = 32'hc4042b7;
      8045: inst = 32'h8220000;
      8046: inst = 32'h10408000;
      8047: inst = 32'hc4042b8;
      8048: inst = 32'h8220000;
      8049: inst = 32'h10408000;
      8050: inst = 32'hc4042b9;
      8051: inst = 32'h8220000;
      8052: inst = 32'h10408000;
      8053: inst = 32'hc4042ba;
      8054: inst = 32'h8220000;
      8055: inst = 32'h10408000;
      8056: inst = 32'hc4042bb;
      8057: inst = 32'h8220000;
      8058: inst = 32'h10408000;
      8059: inst = 32'hc4042bc;
      8060: inst = 32'h8220000;
      8061: inst = 32'h10408000;
      8062: inst = 32'hc4042bd;
      8063: inst = 32'h8220000;
      8064: inst = 32'h10408000;
      8065: inst = 32'hc4042be;
      8066: inst = 32'h8220000;
      8067: inst = 32'h10408000;
      8068: inst = 32'hc4042bf;
      8069: inst = 32'h8220000;
      8070: inst = 32'h10408000;
      8071: inst = 32'hc4042c0;
      8072: inst = 32'h8220000;
      8073: inst = 32'h10408000;
      8074: inst = 32'hc4042c1;
      8075: inst = 32'h8220000;
      8076: inst = 32'h10408000;
      8077: inst = 32'hc4042c2;
      8078: inst = 32'h8220000;
      8079: inst = 32'h10408000;
      8080: inst = 32'hc4042c3;
      8081: inst = 32'h8220000;
      8082: inst = 32'h10408000;
      8083: inst = 32'hc4042fc;
      8084: inst = 32'h8220000;
      8085: inst = 32'h10408000;
      8086: inst = 32'hc4042fd;
      8087: inst = 32'h8220000;
      8088: inst = 32'h10408000;
      8089: inst = 32'hc4042fe;
      8090: inst = 32'h8220000;
      8091: inst = 32'h10408000;
      8092: inst = 32'hc4042ff;
      8093: inst = 32'h8220000;
      8094: inst = 32'h10408000;
      8095: inst = 32'hc404300;
      8096: inst = 32'h8220000;
      8097: inst = 32'h10408000;
      8098: inst = 32'hc404301;
      8099: inst = 32'h8220000;
      8100: inst = 32'h10408000;
      8101: inst = 32'hc404302;
      8102: inst = 32'h8220000;
      8103: inst = 32'h10408000;
      8104: inst = 32'hc404303;
      8105: inst = 32'h8220000;
      8106: inst = 32'h10408000;
      8107: inst = 32'hc404304;
      8108: inst = 32'h8220000;
      8109: inst = 32'h10408000;
      8110: inst = 32'hc404305;
      8111: inst = 32'h8220000;
      8112: inst = 32'h10408000;
      8113: inst = 32'hc404306;
      8114: inst = 32'h8220000;
      8115: inst = 32'h10408000;
      8116: inst = 32'hc404307;
      8117: inst = 32'h8220000;
      8118: inst = 32'h10408000;
      8119: inst = 32'hc404308;
      8120: inst = 32'h8220000;
      8121: inst = 32'h10408000;
      8122: inst = 32'hc404309;
      8123: inst = 32'h8220000;
      8124: inst = 32'h10408000;
      8125: inst = 32'hc40430a;
      8126: inst = 32'h8220000;
      8127: inst = 32'h10408000;
      8128: inst = 32'hc40430b;
      8129: inst = 32'h8220000;
      8130: inst = 32'h10408000;
      8131: inst = 32'hc40430c;
      8132: inst = 32'h8220000;
      8133: inst = 32'h10408000;
      8134: inst = 32'hc40430d;
      8135: inst = 32'h8220000;
      8136: inst = 32'h10408000;
      8137: inst = 32'hc40430e;
      8138: inst = 32'h8220000;
      8139: inst = 32'h10408000;
      8140: inst = 32'hc40430f;
      8141: inst = 32'h8220000;
      8142: inst = 32'h10408000;
      8143: inst = 32'hc404310;
      8144: inst = 32'h8220000;
      8145: inst = 32'h10408000;
      8146: inst = 32'hc404311;
      8147: inst = 32'h8220000;
      8148: inst = 32'h10408000;
      8149: inst = 32'hc404312;
      8150: inst = 32'h8220000;
      8151: inst = 32'h10408000;
      8152: inst = 32'hc404313;
      8153: inst = 32'h8220000;
      8154: inst = 32'h10408000;
      8155: inst = 32'hc404314;
      8156: inst = 32'h8220000;
      8157: inst = 32'h10408000;
      8158: inst = 32'hc404315;
      8159: inst = 32'h8220000;
      8160: inst = 32'h10408000;
      8161: inst = 32'hc404316;
      8162: inst = 32'h8220000;
      8163: inst = 32'h10408000;
      8164: inst = 32'hc404317;
      8165: inst = 32'h8220000;
      8166: inst = 32'h10408000;
      8167: inst = 32'hc404318;
      8168: inst = 32'h8220000;
      8169: inst = 32'h10408000;
      8170: inst = 32'hc404319;
      8171: inst = 32'h8220000;
      8172: inst = 32'h10408000;
      8173: inst = 32'hc40431a;
      8174: inst = 32'h8220000;
      8175: inst = 32'h10408000;
      8176: inst = 32'hc40431b;
      8177: inst = 32'h8220000;
      8178: inst = 32'h10408000;
      8179: inst = 32'hc40431c;
      8180: inst = 32'h8220000;
      8181: inst = 32'h10408000;
      8182: inst = 32'hc40431d;
      8183: inst = 32'h8220000;
      8184: inst = 32'h10408000;
      8185: inst = 32'hc40431e;
      8186: inst = 32'h8220000;
      8187: inst = 32'h10408000;
      8188: inst = 32'hc40431f;
      8189: inst = 32'h8220000;
      8190: inst = 32'h10408000;
      8191: inst = 32'hc404320;
      8192: inst = 32'h8220000;
      8193: inst = 32'h10408000;
      8194: inst = 32'hc404321;
      8195: inst = 32'h8220000;
      8196: inst = 32'h10408000;
      8197: inst = 32'hc404322;
      8198: inst = 32'h8220000;
      8199: inst = 32'h10408000;
      8200: inst = 32'hc404323;
      8201: inst = 32'h8220000;
      8202: inst = 32'h10408000;
      8203: inst = 32'hc40435c;
      8204: inst = 32'h8220000;
      8205: inst = 32'h10408000;
      8206: inst = 32'hc40435d;
      8207: inst = 32'h8220000;
      8208: inst = 32'h10408000;
      8209: inst = 32'hc40435e;
      8210: inst = 32'h8220000;
      8211: inst = 32'h10408000;
      8212: inst = 32'hc40435f;
      8213: inst = 32'h8220000;
      8214: inst = 32'h10408000;
      8215: inst = 32'hc404360;
      8216: inst = 32'h8220000;
      8217: inst = 32'h10408000;
      8218: inst = 32'hc404361;
      8219: inst = 32'h8220000;
      8220: inst = 32'h10408000;
      8221: inst = 32'hc404362;
      8222: inst = 32'h8220000;
      8223: inst = 32'h10408000;
      8224: inst = 32'hc404363;
      8225: inst = 32'h8220000;
      8226: inst = 32'h10408000;
      8227: inst = 32'hc404364;
      8228: inst = 32'h8220000;
      8229: inst = 32'h10408000;
      8230: inst = 32'hc404365;
      8231: inst = 32'h8220000;
      8232: inst = 32'h10408000;
      8233: inst = 32'hc404366;
      8234: inst = 32'h8220000;
      8235: inst = 32'h10408000;
      8236: inst = 32'hc404367;
      8237: inst = 32'h8220000;
      8238: inst = 32'h10408000;
      8239: inst = 32'hc404368;
      8240: inst = 32'h8220000;
      8241: inst = 32'h10408000;
      8242: inst = 32'hc404369;
      8243: inst = 32'h8220000;
      8244: inst = 32'h10408000;
      8245: inst = 32'hc40436a;
      8246: inst = 32'h8220000;
      8247: inst = 32'h10408000;
      8248: inst = 32'hc40436b;
      8249: inst = 32'h8220000;
      8250: inst = 32'h10408000;
      8251: inst = 32'hc40436c;
      8252: inst = 32'h8220000;
      8253: inst = 32'h10408000;
      8254: inst = 32'hc40436d;
      8255: inst = 32'h8220000;
      8256: inst = 32'h10408000;
      8257: inst = 32'hc40436e;
      8258: inst = 32'h8220000;
      8259: inst = 32'h10408000;
      8260: inst = 32'hc40436f;
      8261: inst = 32'h8220000;
      8262: inst = 32'h10408000;
      8263: inst = 32'hc404370;
      8264: inst = 32'h8220000;
      8265: inst = 32'h10408000;
      8266: inst = 32'hc404371;
      8267: inst = 32'h8220000;
      8268: inst = 32'h10408000;
      8269: inst = 32'hc404372;
      8270: inst = 32'h8220000;
      8271: inst = 32'h10408000;
      8272: inst = 32'hc404373;
      8273: inst = 32'h8220000;
      8274: inst = 32'h10408000;
      8275: inst = 32'hc404374;
      8276: inst = 32'h8220000;
      8277: inst = 32'h10408000;
      8278: inst = 32'hc404375;
      8279: inst = 32'h8220000;
      8280: inst = 32'h10408000;
      8281: inst = 32'hc404376;
      8282: inst = 32'h8220000;
      8283: inst = 32'h10408000;
      8284: inst = 32'hc404377;
      8285: inst = 32'h8220000;
      8286: inst = 32'h10408000;
      8287: inst = 32'hc404378;
      8288: inst = 32'h8220000;
      8289: inst = 32'h10408000;
      8290: inst = 32'hc404379;
      8291: inst = 32'h8220000;
      8292: inst = 32'h10408000;
      8293: inst = 32'hc40437a;
      8294: inst = 32'h8220000;
      8295: inst = 32'h10408000;
      8296: inst = 32'hc40437b;
      8297: inst = 32'h8220000;
      8298: inst = 32'h10408000;
      8299: inst = 32'hc40437c;
      8300: inst = 32'h8220000;
      8301: inst = 32'h10408000;
      8302: inst = 32'hc40437d;
      8303: inst = 32'h8220000;
      8304: inst = 32'h10408000;
      8305: inst = 32'hc40437e;
      8306: inst = 32'h8220000;
      8307: inst = 32'h10408000;
      8308: inst = 32'hc40437f;
      8309: inst = 32'h8220000;
      8310: inst = 32'h10408000;
      8311: inst = 32'hc404380;
      8312: inst = 32'h8220000;
      8313: inst = 32'h10408000;
      8314: inst = 32'hc404381;
      8315: inst = 32'h8220000;
      8316: inst = 32'h10408000;
      8317: inst = 32'hc404382;
      8318: inst = 32'h8220000;
      8319: inst = 32'h10408000;
      8320: inst = 32'hc404383;
      8321: inst = 32'h8220000;
      8322: inst = 32'h10408000;
      8323: inst = 32'hc4043bc;
      8324: inst = 32'h8220000;
      8325: inst = 32'h10408000;
      8326: inst = 32'hc4043bd;
      8327: inst = 32'h8220000;
      8328: inst = 32'h10408000;
      8329: inst = 32'hc4043be;
      8330: inst = 32'h8220000;
      8331: inst = 32'h10408000;
      8332: inst = 32'hc4043bf;
      8333: inst = 32'h8220000;
      8334: inst = 32'h10408000;
      8335: inst = 32'hc4043c0;
      8336: inst = 32'h8220000;
      8337: inst = 32'h10408000;
      8338: inst = 32'hc4043c1;
      8339: inst = 32'h8220000;
      8340: inst = 32'h10408000;
      8341: inst = 32'hc4043c2;
      8342: inst = 32'h8220000;
      8343: inst = 32'h10408000;
      8344: inst = 32'hc4043c3;
      8345: inst = 32'h8220000;
      8346: inst = 32'h10408000;
      8347: inst = 32'hc4043c4;
      8348: inst = 32'h8220000;
      8349: inst = 32'h10408000;
      8350: inst = 32'hc4043c5;
      8351: inst = 32'h8220000;
      8352: inst = 32'h10408000;
      8353: inst = 32'hc4043c6;
      8354: inst = 32'h8220000;
      8355: inst = 32'h10408000;
      8356: inst = 32'hc4043c7;
      8357: inst = 32'h8220000;
      8358: inst = 32'h10408000;
      8359: inst = 32'hc4043c8;
      8360: inst = 32'h8220000;
      8361: inst = 32'h10408000;
      8362: inst = 32'hc4043c9;
      8363: inst = 32'h8220000;
      8364: inst = 32'h10408000;
      8365: inst = 32'hc4043ca;
      8366: inst = 32'h8220000;
      8367: inst = 32'h10408000;
      8368: inst = 32'hc4043cb;
      8369: inst = 32'h8220000;
      8370: inst = 32'h10408000;
      8371: inst = 32'hc4043cc;
      8372: inst = 32'h8220000;
      8373: inst = 32'h10408000;
      8374: inst = 32'hc4043cd;
      8375: inst = 32'h8220000;
      8376: inst = 32'h10408000;
      8377: inst = 32'hc4043ce;
      8378: inst = 32'h8220000;
      8379: inst = 32'h10408000;
      8380: inst = 32'hc4043cf;
      8381: inst = 32'h8220000;
      8382: inst = 32'h10408000;
      8383: inst = 32'hc4043d0;
      8384: inst = 32'h8220000;
      8385: inst = 32'h10408000;
      8386: inst = 32'hc4043d1;
      8387: inst = 32'h8220000;
      8388: inst = 32'h10408000;
      8389: inst = 32'hc4043d2;
      8390: inst = 32'h8220000;
      8391: inst = 32'h10408000;
      8392: inst = 32'hc4043d3;
      8393: inst = 32'h8220000;
      8394: inst = 32'h10408000;
      8395: inst = 32'hc4043d4;
      8396: inst = 32'h8220000;
      8397: inst = 32'h10408000;
      8398: inst = 32'hc4043d5;
      8399: inst = 32'h8220000;
      8400: inst = 32'h10408000;
      8401: inst = 32'hc4043d6;
      8402: inst = 32'h8220000;
      8403: inst = 32'h10408000;
      8404: inst = 32'hc4043d7;
      8405: inst = 32'h8220000;
      8406: inst = 32'h10408000;
      8407: inst = 32'hc4043d8;
      8408: inst = 32'h8220000;
      8409: inst = 32'h10408000;
      8410: inst = 32'hc4043d9;
      8411: inst = 32'h8220000;
      8412: inst = 32'h10408000;
      8413: inst = 32'hc4043da;
      8414: inst = 32'h8220000;
      8415: inst = 32'h10408000;
      8416: inst = 32'hc4043db;
      8417: inst = 32'h8220000;
      8418: inst = 32'h10408000;
      8419: inst = 32'hc4043dc;
      8420: inst = 32'h8220000;
      8421: inst = 32'h10408000;
      8422: inst = 32'hc4043dd;
      8423: inst = 32'h8220000;
      8424: inst = 32'h10408000;
      8425: inst = 32'hc4043de;
      8426: inst = 32'h8220000;
      8427: inst = 32'h10408000;
      8428: inst = 32'hc4043df;
      8429: inst = 32'h8220000;
      8430: inst = 32'h10408000;
      8431: inst = 32'hc4043e0;
      8432: inst = 32'h8220000;
      8433: inst = 32'h10408000;
      8434: inst = 32'hc4043e1;
      8435: inst = 32'h8220000;
      8436: inst = 32'h10408000;
      8437: inst = 32'hc4043e2;
      8438: inst = 32'h8220000;
      8439: inst = 32'h10408000;
      8440: inst = 32'hc4043e3;
      8441: inst = 32'h8220000;
      8442: inst = 32'h10408000;
      8443: inst = 32'hc40441c;
      8444: inst = 32'h8220000;
      8445: inst = 32'h10408000;
      8446: inst = 32'hc40441d;
      8447: inst = 32'h8220000;
      8448: inst = 32'h10408000;
      8449: inst = 32'hc40441e;
      8450: inst = 32'h8220000;
      8451: inst = 32'h10408000;
      8452: inst = 32'hc40441f;
      8453: inst = 32'h8220000;
      8454: inst = 32'h10408000;
      8455: inst = 32'hc404420;
      8456: inst = 32'h8220000;
      8457: inst = 32'h10408000;
      8458: inst = 32'hc404421;
      8459: inst = 32'h8220000;
      8460: inst = 32'h10408000;
      8461: inst = 32'hc404422;
      8462: inst = 32'h8220000;
      8463: inst = 32'h10408000;
      8464: inst = 32'hc404423;
      8465: inst = 32'h8220000;
      8466: inst = 32'h10408000;
      8467: inst = 32'hc404424;
      8468: inst = 32'h8220000;
      8469: inst = 32'h10408000;
      8470: inst = 32'hc404425;
      8471: inst = 32'h8220000;
      8472: inst = 32'h10408000;
      8473: inst = 32'hc404426;
      8474: inst = 32'h8220000;
      8475: inst = 32'h10408000;
      8476: inst = 32'hc404427;
      8477: inst = 32'h8220000;
      8478: inst = 32'h10408000;
      8479: inst = 32'hc404428;
      8480: inst = 32'h8220000;
      8481: inst = 32'h10408000;
      8482: inst = 32'hc404429;
      8483: inst = 32'h8220000;
      8484: inst = 32'h10408000;
      8485: inst = 32'hc40442a;
      8486: inst = 32'h8220000;
      8487: inst = 32'h10408000;
      8488: inst = 32'hc40442b;
      8489: inst = 32'h8220000;
      8490: inst = 32'h10408000;
      8491: inst = 32'hc40442c;
      8492: inst = 32'h8220000;
      8493: inst = 32'h10408000;
      8494: inst = 32'hc40442d;
      8495: inst = 32'h8220000;
      8496: inst = 32'h10408000;
      8497: inst = 32'hc40442e;
      8498: inst = 32'h8220000;
      8499: inst = 32'h10408000;
      8500: inst = 32'hc40442f;
      8501: inst = 32'h8220000;
      8502: inst = 32'h10408000;
      8503: inst = 32'hc404430;
      8504: inst = 32'h8220000;
      8505: inst = 32'h10408000;
      8506: inst = 32'hc404431;
      8507: inst = 32'h8220000;
      8508: inst = 32'h10408000;
      8509: inst = 32'hc404432;
      8510: inst = 32'h8220000;
      8511: inst = 32'h10408000;
      8512: inst = 32'hc404433;
      8513: inst = 32'h8220000;
      8514: inst = 32'h10408000;
      8515: inst = 32'hc404434;
      8516: inst = 32'h8220000;
      8517: inst = 32'h10408000;
      8518: inst = 32'hc404435;
      8519: inst = 32'h8220000;
      8520: inst = 32'h10408000;
      8521: inst = 32'hc404436;
      8522: inst = 32'h8220000;
      8523: inst = 32'h10408000;
      8524: inst = 32'hc404437;
      8525: inst = 32'h8220000;
      8526: inst = 32'h10408000;
      8527: inst = 32'hc404438;
      8528: inst = 32'h8220000;
      8529: inst = 32'h10408000;
      8530: inst = 32'hc404439;
      8531: inst = 32'h8220000;
      8532: inst = 32'h10408000;
      8533: inst = 32'hc40443a;
      8534: inst = 32'h8220000;
      8535: inst = 32'h10408000;
      8536: inst = 32'hc40443b;
      8537: inst = 32'h8220000;
      8538: inst = 32'h10408000;
      8539: inst = 32'hc40443c;
      8540: inst = 32'h8220000;
      8541: inst = 32'h10408000;
      8542: inst = 32'hc40443d;
      8543: inst = 32'h8220000;
      8544: inst = 32'h10408000;
      8545: inst = 32'hc40443e;
      8546: inst = 32'h8220000;
      8547: inst = 32'h10408000;
      8548: inst = 32'hc40443f;
      8549: inst = 32'h8220000;
      8550: inst = 32'h10408000;
      8551: inst = 32'hc404440;
      8552: inst = 32'h8220000;
      8553: inst = 32'h10408000;
      8554: inst = 32'hc404441;
      8555: inst = 32'h8220000;
      8556: inst = 32'h10408000;
      8557: inst = 32'hc404442;
      8558: inst = 32'h8220000;
      8559: inst = 32'h10408000;
      8560: inst = 32'hc404443;
      8561: inst = 32'h8220000;
      8562: inst = 32'h10408000;
      8563: inst = 32'hc40447c;
      8564: inst = 32'h8220000;
      8565: inst = 32'h10408000;
      8566: inst = 32'hc40447d;
      8567: inst = 32'h8220000;
      8568: inst = 32'h10408000;
      8569: inst = 32'hc40447e;
      8570: inst = 32'h8220000;
      8571: inst = 32'h10408000;
      8572: inst = 32'hc40447f;
      8573: inst = 32'h8220000;
      8574: inst = 32'h10408000;
      8575: inst = 32'hc404480;
      8576: inst = 32'h8220000;
      8577: inst = 32'h10408000;
      8578: inst = 32'hc404481;
      8579: inst = 32'h8220000;
      8580: inst = 32'h10408000;
      8581: inst = 32'hc404482;
      8582: inst = 32'h8220000;
      8583: inst = 32'h10408000;
      8584: inst = 32'hc404483;
      8585: inst = 32'h8220000;
      8586: inst = 32'h10408000;
      8587: inst = 32'hc404484;
      8588: inst = 32'h8220000;
      8589: inst = 32'h10408000;
      8590: inst = 32'hc404485;
      8591: inst = 32'h8220000;
      8592: inst = 32'h10408000;
      8593: inst = 32'hc404486;
      8594: inst = 32'h8220000;
      8595: inst = 32'h10408000;
      8596: inst = 32'hc404487;
      8597: inst = 32'h8220000;
      8598: inst = 32'h10408000;
      8599: inst = 32'hc404488;
      8600: inst = 32'h8220000;
      8601: inst = 32'h10408000;
      8602: inst = 32'hc404489;
      8603: inst = 32'h8220000;
      8604: inst = 32'h10408000;
      8605: inst = 32'hc40448a;
      8606: inst = 32'h8220000;
      8607: inst = 32'h10408000;
      8608: inst = 32'hc40448b;
      8609: inst = 32'h8220000;
      8610: inst = 32'h10408000;
      8611: inst = 32'hc40448c;
      8612: inst = 32'h8220000;
      8613: inst = 32'h10408000;
      8614: inst = 32'hc40448d;
      8615: inst = 32'h8220000;
      8616: inst = 32'h10408000;
      8617: inst = 32'hc40448e;
      8618: inst = 32'h8220000;
      8619: inst = 32'h10408000;
      8620: inst = 32'hc40448f;
      8621: inst = 32'h8220000;
      8622: inst = 32'h10408000;
      8623: inst = 32'hc404490;
      8624: inst = 32'h8220000;
      8625: inst = 32'h10408000;
      8626: inst = 32'hc404491;
      8627: inst = 32'h8220000;
      8628: inst = 32'h10408000;
      8629: inst = 32'hc404492;
      8630: inst = 32'h8220000;
      8631: inst = 32'h10408000;
      8632: inst = 32'hc404493;
      8633: inst = 32'h8220000;
      8634: inst = 32'h10408000;
      8635: inst = 32'hc404494;
      8636: inst = 32'h8220000;
      8637: inst = 32'h10408000;
      8638: inst = 32'hc404495;
      8639: inst = 32'h8220000;
      8640: inst = 32'h10408000;
      8641: inst = 32'hc404496;
      8642: inst = 32'h8220000;
      8643: inst = 32'h10408000;
      8644: inst = 32'hc404497;
      8645: inst = 32'h8220000;
      8646: inst = 32'h10408000;
      8647: inst = 32'hc404498;
      8648: inst = 32'h8220000;
      8649: inst = 32'h10408000;
      8650: inst = 32'hc404499;
      8651: inst = 32'h8220000;
      8652: inst = 32'h10408000;
      8653: inst = 32'hc40449a;
      8654: inst = 32'h8220000;
      8655: inst = 32'h10408000;
      8656: inst = 32'hc40449b;
      8657: inst = 32'h8220000;
      8658: inst = 32'h10408000;
      8659: inst = 32'hc40449c;
      8660: inst = 32'h8220000;
      8661: inst = 32'h10408000;
      8662: inst = 32'hc40449d;
      8663: inst = 32'h8220000;
      8664: inst = 32'h10408000;
      8665: inst = 32'hc40449e;
      8666: inst = 32'h8220000;
      8667: inst = 32'h10408000;
      8668: inst = 32'hc40449f;
      8669: inst = 32'h8220000;
      8670: inst = 32'h10408000;
      8671: inst = 32'hc4044a0;
      8672: inst = 32'h8220000;
      8673: inst = 32'h10408000;
      8674: inst = 32'hc4044a1;
      8675: inst = 32'h8220000;
      8676: inst = 32'h10408000;
      8677: inst = 32'hc4044a2;
      8678: inst = 32'h8220000;
      8679: inst = 32'h10408000;
      8680: inst = 32'hc4044a3;
      8681: inst = 32'h8220000;
      8682: inst = 32'h10408000;
      8683: inst = 32'hc4044dc;
      8684: inst = 32'h8220000;
      8685: inst = 32'h10408000;
      8686: inst = 32'hc4044dd;
      8687: inst = 32'h8220000;
      8688: inst = 32'h10408000;
      8689: inst = 32'hc4044de;
      8690: inst = 32'h8220000;
      8691: inst = 32'h10408000;
      8692: inst = 32'hc4044df;
      8693: inst = 32'h8220000;
      8694: inst = 32'h10408000;
      8695: inst = 32'hc4044e0;
      8696: inst = 32'h8220000;
      8697: inst = 32'h10408000;
      8698: inst = 32'hc4044e1;
      8699: inst = 32'h8220000;
      8700: inst = 32'h10408000;
      8701: inst = 32'hc4044e2;
      8702: inst = 32'h8220000;
      8703: inst = 32'h10408000;
      8704: inst = 32'hc4044e3;
      8705: inst = 32'h8220000;
      8706: inst = 32'h10408000;
      8707: inst = 32'hc4044e4;
      8708: inst = 32'h8220000;
      8709: inst = 32'h10408000;
      8710: inst = 32'hc4044e5;
      8711: inst = 32'h8220000;
      8712: inst = 32'h10408000;
      8713: inst = 32'hc4044e6;
      8714: inst = 32'h8220000;
      8715: inst = 32'h10408000;
      8716: inst = 32'hc4044e7;
      8717: inst = 32'h8220000;
      8718: inst = 32'h10408000;
      8719: inst = 32'hc4044e8;
      8720: inst = 32'h8220000;
      8721: inst = 32'h10408000;
      8722: inst = 32'hc4044e9;
      8723: inst = 32'h8220000;
      8724: inst = 32'h10408000;
      8725: inst = 32'hc4044ea;
      8726: inst = 32'h8220000;
      8727: inst = 32'h10408000;
      8728: inst = 32'hc4044eb;
      8729: inst = 32'h8220000;
      8730: inst = 32'h10408000;
      8731: inst = 32'hc4044ec;
      8732: inst = 32'h8220000;
      8733: inst = 32'h10408000;
      8734: inst = 32'hc4044ed;
      8735: inst = 32'h8220000;
      8736: inst = 32'h10408000;
      8737: inst = 32'hc4044ee;
      8738: inst = 32'h8220000;
      8739: inst = 32'h10408000;
      8740: inst = 32'hc4044ef;
      8741: inst = 32'h8220000;
      8742: inst = 32'h10408000;
      8743: inst = 32'hc4044f0;
      8744: inst = 32'h8220000;
      8745: inst = 32'h10408000;
      8746: inst = 32'hc4044f1;
      8747: inst = 32'h8220000;
      8748: inst = 32'h10408000;
      8749: inst = 32'hc4044f2;
      8750: inst = 32'h8220000;
      8751: inst = 32'h10408000;
      8752: inst = 32'hc4044f3;
      8753: inst = 32'h8220000;
      8754: inst = 32'h10408000;
      8755: inst = 32'hc4044f4;
      8756: inst = 32'h8220000;
      8757: inst = 32'h10408000;
      8758: inst = 32'hc4044f5;
      8759: inst = 32'h8220000;
      8760: inst = 32'h10408000;
      8761: inst = 32'hc4044f6;
      8762: inst = 32'h8220000;
      8763: inst = 32'h10408000;
      8764: inst = 32'hc4044f7;
      8765: inst = 32'h8220000;
      8766: inst = 32'h10408000;
      8767: inst = 32'hc4044f8;
      8768: inst = 32'h8220000;
      8769: inst = 32'h10408000;
      8770: inst = 32'hc4044f9;
      8771: inst = 32'h8220000;
      8772: inst = 32'h10408000;
      8773: inst = 32'hc4044fa;
      8774: inst = 32'h8220000;
      8775: inst = 32'h10408000;
      8776: inst = 32'hc4044fb;
      8777: inst = 32'h8220000;
      8778: inst = 32'h10408000;
      8779: inst = 32'hc4044fc;
      8780: inst = 32'h8220000;
      8781: inst = 32'h10408000;
      8782: inst = 32'hc4044fd;
      8783: inst = 32'h8220000;
      8784: inst = 32'h10408000;
      8785: inst = 32'hc4044fe;
      8786: inst = 32'h8220000;
      8787: inst = 32'h10408000;
      8788: inst = 32'hc4044ff;
      8789: inst = 32'h8220000;
      8790: inst = 32'h10408000;
      8791: inst = 32'hc404500;
      8792: inst = 32'h8220000;
      8793: inst = 32'h10408000;
      8794: inst = 32'hc404501;
      8795: inst = 32'h8220000;
      8796: inst = 32'h10408000;
      8797: inst = 32'hc404502;
      8798: inst = 32'h8220000;
      8799: inst = 32'h10408000;
      8800: inst = 32'hc404503;
      8801: inst = 32'h8220000;
      8802: inst = 32'h10408000;
      8803: inst = 32'hc40453c;
      8804: inst = 32'h8220000;
      8805: inst = 32'h10408000;
      8806: inst = 32'hc40453d;
      8807: inst = 32'h8220000;
      8808: inst = 32'h10408000;
      8809: inst = 32'hc40453e;
      8810: inst = 32'h8220000;
      8811: inst = 32'h10408000;
      8812: inst = 32'hc40453f;
      8813: inst = 32'h8220000;
      8814: inst = 32'h10408000;
      8815: inst = 32'hc404540;
      8816: inst = 32'h8220000;
      8817: inst = 32'h10408000;
      8818: inst = 32'hc404541;
      8819: inst = 32'h8220000;
      8820: inst = 32'h10408000;
      8821: inst = 32'hc404542;
      8822: inst = 32'h8220000;
      8823: inst = 32'h10408000;
      8824: inst = 32'hc404543;
      8825: inst = 32'h8220000;
      8826: inst = 32'h10408000;
      8827: inst = 32'hc404544;
      8828: inst = 32'h8220000;
      8829: inst = 32'h10408000;
      8830: inst = 32'hc404545;
      8831: inst = 32'h8220000;
      8832: inst = 32'h10408000;
      8833: inst = 32'hc404546;
      8834: inst = 32'h8220000;
      8835: inst = 32'h10408000;
      8836: inst = 32'hc404547;
      8837: inst = 32'h8220000;
      8838: inst = 32'h10408000;
      8839: inst = 32'hc404548;
      8840: inst = 32'h8220000;
      8841: inst = 32'h10408000;
      8842: inst = 32'hc404549;
      8843: inst = 32'h8220000;
      8844: inst = 32'h10408000;
      8845: inst = 32'hc40454a;
      8846: inst = 32'h8220000;
      8847: inst = 32'h10408000;
      8848: inst = 32'hc40454b;
      8849: inst = 32'h8220000;
      8850: inst = 32'h10408000;
      8851: inst = 32'hc40454c;
      8852: inst = 32'h8220000;
      8853: inst = 32'h10408000;
      8854: inst = 32'hc40454d;
      8855: inst = 32'h8220000;
      8856: inst = 32'h10408000;
      8857: inst = 32'hc40454e;
      8858: inst = 32'h8220000;
      8859: inst = 32'h10408000;
      8860: inst = 32'hc40454f;
      8861: inst = 32'h8220000;
      8862: inst = 32'h10408000;
      8863: inst = 32'hc404550;
      8864: inst = 32'h8220000;
      8865: inst = 32'h10408000;
      8866: inst = 32'hc404551;
      8867: inst = 32'h8220000;
      8868: inst = 32'h10408000;
      8869: inst = 32'hc404552;
      8870: inst = 32'h8220000;
      8871: inst = 32'h10408000;
      8872: inst = 32'hc404553;
      8873: inst = 32'h8220000;
      8874: inst = 32'h10408000;
      8875: inst = 32'hc404554;
      8876: inst = 32'h8220000;
      8877: inst = 32'h10408000;
      8878: inst = 32'hc404555;
      8879: inst = 32'h8220000;
      8880: inst = 32'h10408000;
      8881: inst = 32'hc404556;
      8882: inst = 32'h8220000;
      8883: inst = 32'h10408000;
      8884: inst = 32'hc404557;
      8885: inst = 32'h8220000;
      8886: inst = 32'h10408000;
      8887: inst = 32'hc404558;
      8888: inst = 32'h8220000;
      8889: inst = 32'h10408000;
      8890: inst = 32'hc404559;
      8891: inst = 32'h8220000;
      8892: inst = 32'h10408000;
      8893: inst = 32'hc40455a;
      8894: inst = 32'h8220000;
      8895: inst = 32'h10408000;
      8896: inst = 32'hc40455b;
      8897: inst = 32'h8220000;
      8898: inst = 32'h10408000;
      8899: inst = 32'hc40455c;
      8900: inst = 32'h8220000;
      8901: inst = 32'h10408000;
      8902: inst = 32'hc40455d;
      8903: inst = 32'h8220000;
      8904: inst = 32'h10408000;
      8905: inst = 32'hc40455e;
      8906: inst = 32'h8220000;
      8907: inst = 32'h10408000;
      8908: inst = 32'hc40455f;
      8909: inst = 32'h8220000;
      8910: inst = 32'h10408000;
      8911: inst = 32'hc404560;
      8912: inst = 32'h8220000;
      8913: inst = 32'h10408000;
      8914: inst = 32'hc404561;
      8915: inst = 32'h8220000;
      8916: inst = 32'h10408000;
      8917: inst = 32'hc404562;
      8918: inst = 32'h8220000;
      8919: inst = 32'h10408000;
      8920: inst = 32'hc404563;
      8921: inst = 32'h8220000;
      8922: inst = 32'h10408000;
      8923: inst = 32'hc40459c;
      8924: inst = 32'h8220000;
      8925: inst = 32'h10408000;
      8926: inst = 32'hc40459d;
      8927: inst = 32'h8220000;
      8928: inst = 32'h10408000;
      8929: inst = 32'hc40459e;
      8930: inst = 32'h8220000;
      8931: inst = 32'h10408000;
      8932: inst = 32'hc40459f;
      8933: inst = 32'h8220000;
      8934: inst = 32'h10408000;
      8935: inst = 32'hc4045a0;
      8936: inst = 32'h8220000;
      8937: inst = 32'h10408000;
      8938: inst = 32'hc4045a1;
      8939: inst = 32'h8220000;
      8940: inst = 32'h10408000;
      8941: inst = 32'hc4045a2;
      8942: inst = 32'h8220000;
      8943: inst = 32'h10408000;
      8944: inst = 32'hc4045a3;
      8945: inst = 32'h8220000;
      8946: inst = 32'h10408000;
      8947: inst = 32'hc4045a4;
      8948: inst = 32'h8220000;
      8949: inst = 32'h10408000;
      8950: inst = 32'hc4045a5;
      8951: inst = 32'h8220000;
      8952: inst = 32'h10408000;
      8953: inst = 32'hc4045a6;
      8954: inst = 32'h8220000;
      8955: inst = 32'h10408000;
      8956: inst = 32'hc4045a7;
      8957: inst = 32'h8220000;
      8958: inst = 32'h10408000;
      8959: inst = 32'hc4045a8;
      8960: inst = 32'h8220000;
      8961: inst = 32'h10408000;
      8962: inst = 32'hc4045a9;
      8963: inst = 32'h8220000;
      8964: inst = 32'h10408000;
      8965: inst = 32'hc4045aa;
      8966: inst = 32'h8220000;
      8967: inst = 32'h10408000;
      8968: inst = 32'hc4045ab;
      8969: inst = 32'h8220000;
      8970: inst = 32'h10408000;
      8971: inst = 32'hc4045ac;
      8972: inst = 32'h8220000;
      8973: inst = 32'h10408000;
      8974: inst = 32'hc4045ad;
      8975: inst = 32'h8220000;
      8976: inst = 32'h10408000;
      8977: inst = 32'hc4045ae;
      8978: inst = 32'h8220000;
      8979: inst = 32'h10408000;
      8980: inst = 32'hc4045af;
      8981: inst = 32'h8220000;
      8982: inst = 32'h10408000;
      8983: inst = 32'hc4045b0;
      8984: inst = 32'h8220000;
      8985: inst = 32'h10408000;
      8986: inst = 32'hc4045b1;
      8987: inst = 32'h8220000;
      8988: inst = 32'h10408000;
      8989: inst = 32'hc4045b2;
      8990: inst = 32'h8220000;
      8991: inst = 32'h10408000;
      8992: inst = 32'hc4045b3;
      8993: inst = 32'h8220000;
      8994: inst = 32'h10408000;
      8995: inst = 32'hc4045b4;
      8996: inst = 32'h8220000;
      8997: inst = 32'h10408000;
      8998: inst = 32'hc4045b5;
      8999: inst = 32'h8220000;
      9000: inst = 32'h10408000;
      9001: inst = 32'hc4045b6;
      9002: inst = 32'h8220000;
      9003: inst = 32'h10408000;
      9004: inst = 32'hc4045b7;
      9005: inst = 32'h8220000;
      9006: inst = 32'h10408000;
      9007: inst = 32'hc4045b8;
      9008: inst = 32'h8220000;
      9009: inst = 32'h10408000;
      9010: inst = 32'hc4045b9;
      9011: inst = 32'h8220000;
      9012: inst = 32'h10408000;
      9013: inst = 32'hc4045ba;
      9014: inst = 32'h8220000;
      9015: inst = 32'h10408000;
      9016: inst = 32'hc4045bb;
      9017: inst = 32'h8220000;
      9018: inst = 32'h10408000;
      9019: inst = 32'hc4045bc;
      9020: inst = 32'h8220000;
      9021: inst = 32'h10408000;
      9022: inst = 32'hc4045bd;
      9023: inst = 32'h8220000;
      9024: inst = 32'h10408000;
      9025: inst = 32'hc4045be;
      9026: inst = 32'h8220000;
      9027: inst = 32'h10408000;
      9028: inst = 32'hc4045bf;
      9029: inst = 32'h8220000;
      9030: inst = 32'h10408000;
      9031: inst = 32'hc4045c0;
      9032: inst = 32'h8220000;
      9033: inst = 32'h10408000;
      9034: inst = 32'hc4045c1;
      9035: inst = 32'h8220000;
      9036: inst = 32'h10408000;
      9037: inst = 32'hc4045c2;
      9038: inst = 32'h8220000;
      9039: inst = 32'h10408000;
      9040: inst = 32'hc4045c3;
      9041: inst = 32'h8220000;
      9042: inst = 32'h10408000;
      9043: inst = 32'hc4045fc;
      9044: inst = 32'h8220000;
      9045: inst = 32'h10408000;
      9046: inst = 32'hc4045fd;
      9047: inst = 32'h8220000;
      9048: inst = 32'h10408000;
      9049: inst = 32'hc4045fe;
      9050: inst = 32'h8220000;
      9051: inst = 32'h10408000;
      9052: inst = 32'hc4045ff;
      9053: inst = 32'h8220000;
      9054: inst = 32'h10408000;
      9055: inst = 32'hc404600;
      9056: inst = 32'h8220000;
      9057: inst = 32'h10408000;
      9058: inst = 32'hc404601;
      9059: inst = 32'h8220000;
      9060: inst = 32'h10408000;
      9061: inst = 32'hc404602;
      9062: inst = 32'h8220000;
      9063: inst = 32'h10408000;
      9064: inst = 32'hc404603;
      9065: inst = 32'h8220000;
      9066: inst = 32'h10408000;
      9067: inst = 32'hc404604;
      9068: inst = 32'h8220000;
      9069: inst = 32'h10408000;
      9070: inst = 32'hc404605;
      9071: inst = 32'h8220000;
      9072: inst = 32'h10408000;
      9073: inst = 32'hc404606;
      9074: inst = 32'h8220000;
      9075: inst = 32'h10408000;
      9076: inst = 32'hc404607;
      9077: inst = 32'h8220000;
      9078: inst = 32'h10408000;
      9079: inst = 32'hc404608;
      9080: inst = 32'h8220000;
      9081: inst = 32'h10408000;
      9082: inst = 32'hc404609;
      9083: inst = 32'h8220000;
      9084: inst = 32'h10408000;
      9085: inst = 32'hc40460a;
      9086: inst = 32'h8220000;
      9087: inst = 32'h10408000;
      9088: inst = 32'hc40460b;
      9089: inst = 32'h8220000;
      9090: inst = 32'h10408000;
      9091: inst = 32'hc40460c;
      9092: inst = 32'h8220000;
      9093: inst = 32'h10408000;
      9094: inst = 32'hc40460d;
      9095: inst = 32'h8220000;
      9096: inst = 32'h10408000;
      9097: inst = 32'hc40460e;
      9098: inst = 32'h8220000;
      9099: inst = 32'h10408000;
      9100: inst = 32'hc40460f;
      9101: inst = 32'h8220000;
      9102: inst = 32'h10408000;
      9103: inst = 32'hc404610;
      9104: inst = 32'h8220000;
      9105: inst = 32'h10408000;
      9106: inst = 32'hc404611;
      9107: inst = 32'h8220000;
      9108: inst = 32'h10408000;
      9109: inst = 32'hc404612;
      9110: inst = 32'h8220000;
      9111: inst = 32'h10408000;
      9112: inst = 32'hc404613;
      9113: inst = 32'h8220000;
      9114: inst = 32'h10408000;
      9115: inst = 32'hc404614;
      9116: inst = 32'h8220000;
      9117: inst = 32'h10408000;
      9118: inst = 32'hc404615;
      9119: inst = 32'h8220000;
      9120: inst = 32'h10408000;
      9121: inst = 32'hc404616;
      9122: inst = 32'h8220000;
      9123: inst = 32'h10408000;
      9124: inst = 32'hc404617;
      9125: inst = 32'h8220000;
      9126: inst = 32'h10408000;
      9127: inst = 32'hc404618;
      9128: inst = 32'h8220000;
      9129: inst = 32'h10408000;
      9130: inst = 32'hc404619;
      9131: inst = 32'h8220000;
      9132: inst = 32'h10408000;
      9133: inst = 32'hc40461a;
      9134: inst = 32'h8220000;
      9135: inst = 32'h10408000;
      9136: inst = 32'hc40461b;
      9137: inst = 32'h8220000;
      9138: inst = 32'h10408000;
      9139: inst = 32'hc40461c;
      9140: inst = 32'h8220000;
      9141: inst = 32'h10408000;
      9142: inst = 32'hc40461d;
      9143: inst = 32'h8220000;
      9144: inst = 32'h10408000;
      9145: inst = 32'hc40461e;
      9146: inst = 32'h8220000;
      9147: inst = 32'h10408000;
      9148: inst = 32'hc40461f;
      9149: inst = 32'h8220000;
      9150: inst = 32'h10408000;
      9151: inst = 32'hc404620;
      9152: inst = 32'h8220000;
      9153: inst = 32'h10408000;
      9154: inst = 32'hc404621;
      9155: inst = 32'h8220000;
      9156: inst = 32'h10408000;
      9157: inst = 32'hc404622;
      9158: inst = 32'h8220000;
      9159: inst = 32'h10408000;
      9160: inst = 32'hc404623;
      9161: inst = 32'h8220000;
      9162: inst = 32'h10408000;
      9163: inst = 32'hc40465c;
      9164: inst = 32'h8220000;
      9165: inst = 32'h10408000;
      9166: inst = 32'hc40465d;
      9167: inst = 32'h8220000;
      9168: inst = 32'h10408000;
      9169: inst = 32'hc40465e;
      9170: inst = 32'h8220000;
      9171: inst = 32'h10408000;
      9172: inst = 32'hc40465f;
      9173: inst = 32'h8220000;
      9174: inst = 32'h10408000;
      9175: inst = 32'hc404660;
      9176: inst = 32'h8220000;
      9177: inst = 32'h10408000;
      9178: inst = 32'hc404661;
      9179: inst = 32'h8220000;
      9180: inst = 32'h10408000;
      9181: inst = 32'hc404662;
      9182: inst = 32'h8220000;
      9183: inst = 32'h10408000;
      9184: inst = 32'hc404663;
      9185: inst = 32'h8220000;
      9186: inst = 32'h10408000;
      9187: inst = 32'hc404664;
      9188: inst = 32'h8220000;
      9189: inst = 32'h10408000;
      9190: inst = 32'hc404665;
      9191: inst = 32'h8220000;
      9192: inst = 32'h10408000;
      9193: inst = 32'hc404666;
      9194: inst = 32'h8220000;
      9195: inst = 32'h10408000;
      9196: inst = 32'hc404667;
      9197: inst = 32'h8220000;
      9198: inst = 32'h10408000;
      9199: inst = 32'hc404668;
      9200: inst = 32'h8220000;
      9201: inst = 32'h10408000;
      9202: inst = 32'hc404669;
      9203: inst = 32'h8220000;
      9204: inst = 32'h10408000;
      9205: inst = 32'hc40466a;
      9206: inst = 32'h8220000;
      9207: inst = 32'h10408000;
      9208: inst = 32'hc40466b;
      9209: inst = 32'h8220000;
      9210: inst = 32'h10408000;
      9211: inst = 32'hc40466c;
      9212: inst = 32'h8220000;
      9213: inst = 32'h10408000;
      9214: inst = 32'hc40466d;
      9215: inst = 32'h8220000;
      9216: inst = 32'h10408000;
      9217: inst = 32'hc40466e;
      9218: inst = 32'h8220000;
      9219: inst = 32'h10408000;
      9220: inst = 32'hc40466f;
      9221: inst = 32'h8220000;
      9222: inst = 32'h10408000;
      9223: inst = 32'hc404670;
      9224: inst = 32'h8220000;
      9225: inst = 32'h10408000;
      9226: inst = 32'hc404671;
      9227: inst = 32'h8220000;
      9228: inst = 32'h10408000;
      9229: inst = 32'hc404672;
      9230: inst = 32'h8220000;
      9231: inst = 32'h10408000;
      9232: inst = 32'hc404673;
      9233: inst = 32'h8220000;
      9234: inst = 32'h10408000;
      9235: inst = 32'hc404674;
      9236: inst = 32'h8220000;
      9237: inst = 32'h10408000;
      9238: inst = 32'hc404675;
      9239: inst = 32'h8220000;
      9240: inst = 32'h10408000;
      9241: inst = 32'hc404676;
      9242: inst = 32'h8220000;
      9243: inst = 32'h10408000;
      9244: inst = 32'hc404677;
      9245: inst = 32'h8220000;
      9246: inst = 32'h10408000;
      9247: inst = 32'hc404678;
      9248: inst = 32'h8220000;
      9249: inst = 32'h10408000;
      9250: inst = 32'hc404679;
      9251: inst = 32'h8220000;
      9252: inst = 32'h10408000;
      9253: inst = 32'hc40467a;
      9254: inst = 32'h8220000;
      9255: inst = 32'h10408000;
      9256: inst = 32'hc40467b;
      9257: inst = 32'h8220000;
      9258: inst = 32'h10408000;
      9259: inst = 32'hc40467c;
      9260: inst = 32'h8220000;
      9261: inst = 32'h10408000;
      9262: inst = 32'hc40467d;
      9263: inst = 32'h8220000;
      9264: inst = 32'h10408000;
      9265: inst = 32'hc40467e;
      9266: inst = 32'h8220000;
      9267: inst = 32'h10408000;
      9268: inst = 32'hc40467f;
      9269: inst = 32'h8220000;
      9270: inst = 32'h10408000;
      9271: inst = 32'hc404680;
      9272: inst = 32'h8220000;
      9273: inst = 32'h10408000;
      9274: inst = 32'hc404681;
      9275: inst = 32'h8220000;
      9276: inst = 32'h10408000;
      9277: inst = 32'hc404682;
      9278: inst = 32'h8220000;
      9279: inst = 32'h10408000;
      9280: inst = 32'hc404683;
      9281: inst = 32'h8220000;
      9282: inst = 32'h10408000;
      9283: inst = 32'hc4046bc;
      9284: inst = 32'h8220000;
      9285: inst = 32'h10408000;
      9286: inst = 32'hc4046bd;
      9287: inst = 32'h8220000;
      9288: inst = 32'h10408000;
      9289: inst = 32'hc4046be;
      9290: inst = 32'h8220000;
      9291: inst = 32'h10408000;
      9292: inst = 32'hc4046bf;
      9293: inst = 32'h8220000;
      9294: inst = 32'h10408000;
      9295: inst = 32'hc4046c0;
      9296: inst = 32'h8220000;
      9297: inst = 32'h10408000;
      9298: inst = 32'hc4046c1;
      9299: inst = 32'h8220000;
      9300: inst = 32'h10408000;
      9301: inst = 32'hc4046c2;
      9302: inst = 32'h8220000;
      9303: inst = 32'h10408000;
      9304: inst = 32'hc4046c3;
      9305: inst = 32'h8220000;
      9306: inst = 32'h10408000;
      9307: inst = 32'hc4046c4;
      9308: inst = 32'h8220000;
      9309: inst = 32'h10408000;
      9310: inst = 32'hc4046c5;
      9311: inst = 32'h8220000;
      9312: inst = 32'h10408000;
      9313: inst = 32'hc4046c6;
      9314: inst = 32'h8220000;
      9315: inst = 32'h10408000;
      9316: inst = 32'hc4046c7;
      9317: inst = 32'h8220000;
      9318: inst = 32'h10408000;
      9319: inst = 32'hc4046c8;
      9320: inst = 32'h8220000;
      9321: inst = 32'h10408000;
      9322: inst = 32'hc4046c9;
      9323: inst = 32'h8220000;
      9324: inst = 32'h10408000;
      9325: inst = 32'hc4046ca;
      9326: inst = 32'h8220000;
      9327: inst = 32'h10408000;
      9328: inst = 32'hc4046cb;
      9329: inst = 32'h8220000;
      9330: inst = 32'h10408000;
      9331: inst = 32'hc4046cc;
      9332: inst = 32'h8220000;
      9333: inst = 32'h10408000;
      9334: inst = 32'hc4046cd;
      9335: inst = 32'h8220000;
      9336: inst = 32'h10408000;
      9337: inst = 32'hc4046ce;
      9338: inst = 32'h8220000;
      9339: inst = 32'h10408000;
      9340: inst = 32'hc4046cf;
      9341: inst = 32'h8220000;
      9342: inst = 32'h10408000;
      9343: inst = 32'hc4046d0;
      9344: inst = 32'h8220000;
      9345: inst = 32'h10408000;
      9346: inst = 32'hc4046d1;
      9347: inst = 32'h8220000;
      9348: inst = 32'h10408000;
      9349: inst = 32'hc4046d2;
      9350: inst = 32'h8220000;
      9351: inst = 32'h10408000;
      9352: inst = 32'hc4046d3;
      9353: inst = 32'h8220000;
      9354: inst = 32'h10408000;
      9355: inst = 32'hc4046d4;
      9356: inst = 32'h8220000;
      9357: inst = 32'h10408000;
      9358: inst = 32'hc4046d5;
      9359: inst = 32'h8220000;
      9360: inst = 32'h10408000;
      9361: inst = 32'hc4046d6;
      9362: inst = 32'h8220000;
      9363: inst = 32'h10408000;
      9364: inst = 32'hc4046d7;
      9365: inst = 32'h8220000;
      9366: inst = 32'h10408000;
      9367: inst = 32'hc4046d8;
      9368: inst = 32'h8220000;
      9369: inst = 32'h10408000;
      9370: inst = 32'hc4046d9;
      9371: inst = 32'h8220000;
      9372: inst = 32'h10408000;
      9373: inst = 32'hc4046da;
      9374: inst = 32'h8220000;
      9375: inst = 32'h10408000;
      9376: inst = 32'hc4046db;
      9377: inst = 32'h8220000;
      9378: inst = 32'h10408000;
      9379: inst = 32'hc4046dc;
      9380: inst = 32'h8220000;
      9381: inst = 32'h10408000;
      9382: inst = 32'hc4046dd;
      9383: inst = 32'h8220000;
      9384: inst = 32'h10408000;
      9385: inst = 32'hc4046de;
      9386: inst = 32'h8220000;
      9387: inst = 32'h10408000;
      9388: inst = 32'hc4046df;
      9389: inst = 32'h8220000;
      9390: inst = 32'h10408000;
      9391: inst = 32'hc4046e0;
      9392: inst = 32'h8220000;
      9393: inst = 32'h10408000;
      9394: inst = 32'hc4046e1;
      9395: inst = 32'h8220000;
      9396: inst = 32'h10408000;
      9397: inst = 32'hc4046e2;
      9398: inst = 32'h8220000;
      9399: inst = 32'h10408000;
      9400: inst = 32'hc4046e3;
      9401: inst = 32'h8220000;
      9402: inst = 32'h10408000;
      9403: inst = 32'hc40471c;
      9404: inst = 32'h8220000;
      9405: inst = 32'h10408000;
      9406: inst = 32'hc40471d;
      9407: inst = 32'h8220000;
      9408: inst = 32'h10408000;
      9409: inst = 32'hc40471e;
      9410: inst = 32'h8220000;
      9411: inst = 32'h10408000;
      9412: inst = 32'hc40471f;
      9413: inst = 32'h8220000;
      9414: inst = 32'h10408000;
      9415: inst = 32'hc404720;
      9416: inst = 32'h8220000;
      9417: inst = 32'h10408000;
      9418: inst = 32'hc404721;
      9419: inst = 32'h8220000;
      9420: inst = 32'h10408000;
      9421: inst = 32'hc404722;
      9422: inst = 32'h8220000;
      9423: inst = 32'h10408000;
      9424: inst = 32'hc404723;
      9425: inst = 32'h8220000;
      9426: inst = 32'h10408000;
      9427: inst = 32'hc404724;
      9428: inst = 32'h8220000;
      9429: inst = 32'h10408000;
      9430: inst = 32'hc404725;
      9431: inst = 32'h8220000;
      9432: inst = 32'h10408000;
      9433: inst = 32'hc404726;
      9434: inst = 32'h8220000;
      9435: inst = 32'h10408000;
      9436: inst = 32'hc404727;
      9437: inst = 32'h8220000;
      9438: inst = 32'h10408000;
      9439: inst = 32'hc404728;
      9440: inst = 32'h8220000;
      9441: inst = 32'h10408000;
      9442: inst = 32'hc404729;
      9443: inst = 32'h8220000;
      9444: inst = 32'h10408000;
      9445: inst = 32'hc40472a;
      9446: inst = 32'h8220000;
      9447: inst = 32'h10408000;
      9448: inst = 32'hc40472b;
      9449: inst = 32'h8220000;
      9450: inst = 32'h10408000;
      9451: inst = 32'hc40472c;
      9452: inst = 32'h8220000;
      9453: inst = 32'h10408000;
      9454: inst = 32'hc40472d;
      9455: inst = 32'h8220000;
      9456: inst = 32'h10408000;
      9457: inst = 32'hc40472e;
      9458: inst = 32'h8220000;
      9459: inst = 32'h10408000;
      9460: inst = 32'hc40472f;
      9461: inst = 32'h8220000;
      9462: inst = 32'h10408000;
      9463: inst = 32'hc404730;
      9464: inst = 32'h8220000;
      9465: inst = 32'h10408000;
      9466: inst = 32'hc404731;
      9467: inst = 32'h8220000;
      9468: inst = 32'h10408000;
      9469: inst = 32'hc404732;
      9470: inst = 32'h8220000;
      9471: inst = 32'h10408000;
      9472: inst = 32'hc404733;
      9473: inst = 32'h8220000;
      9474: inst = 32'h10408000;
      9475: inst = 32'hc404734;
      9476: inst = 32'h8220000;
      9477: inst = 32'h10408000;
      9478: inst = 32'hc404735;
      9479: inst = 32'h8220000;
      9480: inst = 32'h10408000;
      9481: inst = 32'hc404736;
      9482: inst = 32'h8220000;
      9483: inst = 32'h10408000;
      9484: inst = 32'hc404737;
      9485: inst = 32'h8220000;
      9486: inst = 32'h10408000;
      9487: inst = 32'hc404738;
      9488: inst = 32'h8220000;
      9489: inst = 32'h10408000;
      9490: inst = 32'hc404739;
      9491: inst = 32'h8220000;
      9492: inst = 32'h10408000;
      9493: inst = 32'hc40473a;
      9494: inst = 32'h8220000;
      9495: inst = 32'h10408000;
      9496: inst = 32'hc40473b;
      9497: inst = 32'h8220000;
      9498: inst = 32'h10408000;
      9499: inst = 32'hc40473c;
      9500: inst = 32'h8220000;
      9501: inst = 32'h10408000;
      9502: inst = 32'hc40473d;
      9503: inst = 32'h8220000;
      9504: inst = 32'h10408000;
      9505: inst = 32'hc40473e;
      9506: inst = 32'h8220000;
      9507: inst = 32'h10408000;
      9508: inst = 32'hc40473f;
      9509: inst = 32'h8220000;
      9510: inst = 32'h10408000;
      9511: inst = 32'hc404740;
      9512: inst = 32'h8220000;
      9513: inst = 32'h10408000;
      9514: inst = 32'hc404741;
      9515: inst = 32'h8220000;
      9516: inst = 32'h10408000;
      9517: inst = 32'hc404742;
      9518: inst = 32'h8220000;
      9519: inst = 32'h10408000;
      9520: inst = 32'hc404743;
      9521: inst = 32'h8220000;
      9522: inst = 32'h10408000;
      9523: inst = 32'hc40477c;
      9524: inst = 32'h8220000;
      9525: inst = 32'h10408000;
      9526: inst = 32'hc40477d;
      9527: inst = 32'h8220000;
      9528: inst = 32'h10408000;
      9529: inst = 32'hc40477e;
      9530: inst = 32'h8220000;
      9531: inst = 32'h10408000;
      9532: inst = 32'hc40477f;
      9533: inst = 32'h8220000;
      9534: inst = 32'h10408000;
      9535: inst = 32'hc404780;
      9536: inst = 32'h8220000;
      9537: inst = 32'h10408000;
      9538: inst = 32'hc404781;
      9539: inst = 32'h8220000;
      9540: inst = 32'h10408000;
      9541: inst = 32'hc404782;
      9542: inst = 32'h8220000;
      9543: inst = 32'h10408000;
      9544: inst = 32'hc404783;
      9545: inst = 32'h8220000;
      9546: inst = 32'h10408000;
      9547: inst = 32'hc404784;
      9548: inst = 32'h8220000;
      9549: inst = 32'h10408000;
      9550: inst = 32'hc404785;
      9551: inst = 32'h8220000;
      9552: inst = 32'h10408000;
      9553: inst = 32'hc404786;
      9554: inst = 32'h8220000;
      9555: inst = 32'h10408000;
      9556: inst = 32'hc404787;
      9557: inst = 32'h8220000;
      9558: inst = 32'h10408000;
      9559: inst = 32'hc404788;
      9560: inst = 32'h8220000;
      9561: inst = 32'h10408000;
      9562: inst = 32'hc404789;
      9563: inst = 32'h8220000;
      9564: inst = 32'h10408000;
      9565: inst = 32'hc40478a;
      9566: inst = 32'h8220000;
      9567: inst = 32'h10408000;
      9568: inst = 32'hc40478b;
      9569: inst = 32'h8220000;
      9570: inst = 32'h10408000;
      9571: inst = 32'hc40478c;
      9572: inst = 32'h8220000;
      9573: inst = 32'h10408000;
      9574: inst = 32'hc40478d;
      9575: inst = 32'h8220000;
      9576: inst = 32'h10408000;
      9577: inst = 32'hc40478e;
      9578: inst = 32'h8220000;
      9579: inst = 32'h10408000;
      9580: inst = 32'hc40478f;
      9581: inst = 32'h8220000;
      9582: inst = 32'h10408000;
      9583: inst = 32'hc404790;
      9584: inst = 32'h8220000;
      9585: inst = 32'h10408000;
      9586: inst = 32'hc404791;
      9587: inst = 32'h8220000;
      9588: inst = 32'h10408000;
      9589: inst = 32'hc404792;
      9590: inst = 32'h8220000;
      9591: inst = 32'h10408000;
      9592: inst = 32'hc404793;
      9593: inst = 32'h8220000;
      9594: inst = 32'h10408000;
      9595: inst = 32'hc404794;
      9596: inst = 32'h8220000;
      9597: inst = 32'h10408000;
      9598: inst = 32'hc404795;
      9599: inst = 32'h8220000;
      9600: inst = 32'h10408000;
      9601: inst = 32'hc404796;
      9602: inst = 32'h8220000;
      9603: inst = 32'h10408000;
      9604: inst = 32'hc404797;
      9605: inst = 32'h8220000;
      9606: inst = 32'h10408000;
      9607: inst = 32'hc404798;
      9608: inst = 32'h8220000;
      9609: inst = 32'h10408000;
      9610: inst = 32'hc404799;
      9611: inst = 32'h8220000;
      9612: inst = 32'h10408000;
      9613: inst = 32'hc40479a;
      9614: inst = 32'h8220000;
      9615: inst = 32'h10408000;
      9616: inst = 32'hc40479b;
      9617: inst = 32'h8220000;
      9618: inst = 32'h10408000;
      9619: inst = 32'hc40479c;
      9620: inst = 32'h8220000;
      9621: inst = 32'h10408000;
      9622: inst = 32'hc40479d;
      9623: inst = 32'h8220000;
      9624: inst = 32'h10408000;
      9625: inst = 32'hc40479e;
      9626: inst = 32'h8220000;
      9627: inst = 32'h10408000;
      9628: inst = 32'hc40479f;
      9629: inst = 32'h8220000;
      9630: inst = 32'h10408000;
      9631: inst = 32'hc4047a0;
      9632: inst = 32'h8220000;
      9633: inst = 32'h10408000;
      9634: inst = 32'hc4047a1;
      9635: inst = 32'h8220000;
      9636: inst = 32'h10408000;
      9637: inst = 32'hc4047a2;
      9638: inst = 32'h8220000;
      9639: inst = 32'h10408000;
      9640: inst = 32'hc4047a3;
      9641: inst = 32'h8220000;
      9642: inst = 32'h10408000;
      9643: inst = 32'hc4047dc;
      9644: inst = 32'h8220000;
      9645: inst = 32'h10408000;
      9646: inst = 32'hc4047dd;
      9647: inst = 32'h8220000;
      9648: inst = 32'h10408000;
      9649: inst = 32'hc4047de;
      9650: inst = 32'h8220000;
      9651: inst = 32'h10408000;
      9652: inst = 32'hc4047df;
      9653: inst = 32'h8220000;
      9654: inst = 32'h10408000;
      9655: inst = 32'hc4047e0;
      9656: inst = 32'h8220000;
      9657: inst = 32'h10408000;
      9658: inst = 32'hc4047e1;
      9659: inst = 32'h8220000;
      9660: inst = 32'h10408000;
      9661: inst = 32'hc4047e2;
      9662: inst = 32'h8220000;
      9663: inst = 32'h10408000;
      9664: inst = 32'hc4047e3;
      9665: inst = 32'h8220000;
      9666: inst = 32'h10408000;
      9667: inst = 32'hc4047e4;
      9668: inst = 32'h8220000;
      9669: inst = 32'h10408000;
      9670: inst = 32'hc4047e5;
      9671: inst = 32'h8220000;
      9672: inst = 32'h10408000;
      9673: inst = 32'hc4047e6;
      9674: inst = 32'h8220000;
      9675: inst = 32'h10408000;
      9676: inst = 32'hc4047e7;
      9677: inst = 32'h8220000;
      9678: inst = 32'h10408000;
      9679: inst = 32'hc4047e8;
      9680: inst = 32'h8220000;
      9681: inst = 32'h10408000;
      9682: inst = 32'hc4047e9;
      9683: inst = 32'h8220000;
      9684: inst = 32'h10408000;
      9685: inst = 32'hc4047ea;
      9686: inst = 32'h8220000;
      9687: inst = 32'h10408000;
      9688: inst = 32'hc4047eb;
      9689: inst = 32'h8220000;
      9690: inst = 32'h10408000;
      9691: inst = 32'hc4047ec;
      9692: inst = 32'h8220000;
      9693: inst = 32'h10408000;
      9694: inst = 32'hc4047ed;
      9695: inst = 32'h8220000;
      9696: inst = 32'h10408000;
      9697: inst = 32'hc4047ee;
      9698: inst = 32'h8220000;
      9699: inst = 32'h10408000;
      9700: inst = 32'hc4047ef;
      9701: inst = 32'h8220000;
      9702: inst = 32'h10408000;
      9703: inst = 32'hc4047f0;
      9704: inst = 32'h8220000;
      9705: inst = 32'h10408000;
      9706: inst = 32'hc4047f1;
      9707: inst = 32'h8220000;
      9708: inst = 32'h10408000;
      9709: inst = 32'hc4047f2;
      9710: inst = 32'h8220000;
      9711: inst = 32'h10408000;
      9712: inst = 32'hc4047f3;
      9713: inst = 32'h8220000;
      9714: inst = 32'h10408000;
      9715: inst = 32'hc4047f4;
      9716: inst = 32'h8220000;
      9717: inst = 32'h10408000;
      9718: inst = 32'hc4047f5;
      9719: inst = 32'h8220000;
      9720: inst = 32'h10408000;
      9721: inst = 32'hc4047f6;
      9722: inst = 32'h8220000;
      9723: inst = 32'h10408000;
      9724: inst = 32'hc4047f7;
      9725: inst = 32'h8220000;
      9726: inst = 32'h10408000;
      9727: inst = 32'hc4047f8;
      9728: inst = 32'h8220000;
      9729: inst = 32'h10408000;
      9730: inst = 32'hc4047f9;
      9731: inst = 32'h8220000;
      9732: inst = 32'h10408000;
      9733: inst = 32'hc4047fa;
      9734: inst = 32'h8220000;
      9735: inst = 32'h10408000;
      9736: inst = 32'hc4047fb;
      9737: inst = 32'h8220000;
      9738: inst = 32'h10408000;
      9739: inst = 32'hc4047fc;
      9740: inst = 32'h8220000;
      9741: inst = 32'h10408000;
      9742: inst = 32'hc4047fd;
      9743: inst = 32'h8220000;
      9744: inst = 32'h10408000;
      9745: inst = 32'hc4047fe;
      9746: inst = 32'h8220000;
      9747: inst = 32'h10408000;
      9748: inst = 32'hc4047ff;
      9749: inst = 32'h8220000;
      9750: inst = 32'h10408000;
      9751: inst = 32'hc404800;
      9752: inst = 32'h8220000;
      9753: inst = 32'h10408000;
      9754: inst = 32'hc404801;
      9755: inst = 32'h8220000;
      9756: inst = 32'h10408000;
      9757: inst = 32'hc404802;
      9758: inst = 32'h8220000;
      9759: inst = 32'h10408000;
      9760: inst = 32'hc404803;
      9761: inst = 32'h8220000;
      9762: inst = 32'h10408000;
      9763: inst = 32'hc40483c;
      9764: inst = 32'h8220000;
      9765: inst = 32'h10408000;
      9766: inst = 32'hc40483d;
      9767: inst = 32'h8220000;
      9768: inst = 32'h10408000;
      9769: inst = 32'hc40483e;
      9770: inst = 32'h8220000;
      9771: inst = 32'h10408000;
      9772: inst = 32'hc40483f;
      9773: inst = 32'h8220000;
      9774: inst = 32'h10408000;
      9775: inst = 32'hc404840;
      9776: inst = 32'h8220000;
      9777: inst = 32'h10408000;
      9778: inst = 32'hc404841;
      9779: inst = 32'h8220000;
      9780: inst = 32'h10408000;
      9781: inst = 32'hc404842;
      9782: inst = 32'h8220000;
      9783: inst = 32'h10408000;
      9784: inst = 32'hc404843;
      9785: inst = 32'h8220000;
      9786: inst = 32'h10408000;
      9787: inst = 32'hc404844;
      9788: inst = 32'h8220000;
      9789: inst = 32'h10408000;
      9790: inst = 32'hc404845;
      9791: inst = 32'h8220000;
      9792: inst = 32'h10408000;
      9793: inst = 32'hc404846;
      9794: inst = 32'h8220000;
      9795: inst = 32'h10408000;
      9796: inst = 32'hc404847;
      9797: inst = 32'h8220000;
      9798: inst = 32'h10408000;
      9799: inst = 32'hc404848;
      9800: inst = 32'h8220000;
      9801: inst = 32'h10408000;
      9802: inst = 32'hc404849;
      9803: inst = 32'h8220000;
      9804: inst = 32'h10408000;
      9805: inst = 32'hc40484a;
      9806: inst = 32'h8220000;
      9807: inst = 32'h10408000;
      9808: inst = 32'hc40484b;
      9809: inst = 32'h8220000;
      9810: inst = 32'h10408000;
      9811: inst = 32'hc40484c;
      9812: inst = 32'h8220000;
      9813: inst = 32'h10408000;
      9814: inst = 32'hc40484d;
      9815: inst = 32'h8220000;
      9816: inst = 32'h10408000;
      9817: inst = 32'hc40484e;
      9818: inst = 32'h8220000;
      9819: inst = 32'h10408000;
      9820: inst = 32'hc40484f;
      9821: inst = 32'h8220000;
      9822: inst = 32'h10408000;
      9823: inst = 32'hc404850;
      9824: inst = 32'h8220000;
      9825: inst = 32'h10408000;
      9826: inst = 32'hc404851;
      9827: inst = 32'h8220000;
      9828: inst = 32'h10408000;
      9829: inst = 32'hc404852;
      9830: inst = 32'h8220000;
      9831: inst = 32'h10408000;
      9832: inst = 32'hc404853;
      9833: inst = 32'h8220000;
      9834: inst = 32'h10408000;
      9835: inst = 32'hc404854;
      9836: inst = 32'h8220000;
      9837: inst = 32'h10408000;
      9838: inst = 32'hc404855;
      9839: inst = 32'h8220000;
      9840: inst = 32'h10408000;
      9841: inst = 32'hc404856;
      9842: inst = 32'h8220000;
      9843: inst = 32'h10408000;
      9844: inst = 32'hc404857;
      9845: inst = 32'h8220000;
      9846: inst = 32'h10408000;
      9847: inst = 32'hc404858;
      9848: inst = 32'h8220000;
      9849: inst = 32'h10408000;
      9850: inst = 32'hc404859;
      9851: inst = 32'h8220000;
      9852: inst = 32'h10408000;
      9853: inst = 32'hc40485a;
      9854: inst = 32'h8220000;
      9855: inst = 32'h10408000;
      9856: inst = 32'hc40485b;
      9857: inst = 32'h8220000;
      9858: inst = 32'h10408000;
      9859: inst = 32'hc40485c;
      9860: inst = 32'h8220000;
      9861: inst = 32'h10408000;
      9862: inst = 32'hc40485d;
      9863: inst = 32'h8220000;
      9864: inst = 32'h10408000;
      9865: inst = 32'hc40485e;
      9866: inst = 32'h8220000;
      9867: inst = 32'h10408000;
      9868: inst = 32'hc40485f;
      9869: inst = 32'h8220000;
      9870: inst = 32'h10408000;
      9871: inst = 32'hc404860;
      9872: inst = 32'h8220000;
      9873: inst = 32'h10408000;
      9874: inst = 32'hc404861;
      9875: inst = 32'h8220000;
      9876: inst = 32'h10408000;
      9877: inst = 32'hc404862;
      9878: inst = 32'h8220000;
      9879: inst = 32'h10408000;
      9880: inst = 32'hc404863;
      9881: inst = 32'h8220000;
      9882: inst = 32'h10408000;
      9883: inst = 32'hc40489c;
      9884: inst = 32'h8220000;
      9885: inst = 32'h10408000;
      9886: inst = 32'hc40489d;
      9887: inst = 32'h8220000;
      9888: inst = 32'h10408000;
      9889: inst = 32'hc40489e;
      9890: inst = 32'h8220000;
      9891: inst = 32'h10408000;
      9892: inst = 32'hc40489f;
      9893: inst = 32'h8220000;
      9894: inst = 32'h10408000;
      9895: inst = 32'hc4048a0;
      9896: inst = 32'h8220000;
      9897: inst = 32'h10408000;
      9898: inst = 32'hc4048a1;
      9899: inst = 32'h8220000;
      9900: inst = 32'h10408000;
      9901: inst = 32'hc4048a2;
      9902: inst = 32'h8220000;
      9903: inst = 32'h10408000;
      9904: inst = 32'hc4048a3;
      9905: inst = 32'h8220000;
      9906: inst = 32'h10408000;
      9907: inst = 32'hc4048a4;
      9908: inst = 32'h8220000;
      9909: inst = 32'h10408000;
      9910: inst = 32'hc4048a5;
      9911: inst = 32'h8220000;
      9912: inst = 32'h10408000;
      9913: inst = 32'hc4048a6;
      9914: inst = 32'h8220000;
      9915: inst = 32'h10408000;
      9916: inst = 32'hc4048a7;
      9917: inst = 32'h8220000;
      9918: inst = 32'h10408000;
      9919: inst = 32'hc4048a8;
      9920: inst = 32'h8220000;
      9921: inst = 32'h10408000;
      9922: inst = 32'hc4048a9;
      9923: inst = 32'h8220000;
      9924: inst = 32'h10408000;
      9925: inst = 32'hc4048aa;
      9926: inst = 32'h8220000;
      9927: inst = 32'h10408000;
      9928: inst = 32'hc4048ab;
      9929: inst = 32'h8220000;
      9930: inst = 32'h10408000;
      9931: inst = 32'hc4048ac;
      9932: inst = 32'h8220000;
      9933: inst = 32'h10408000;
      9934: inst = 32'hc4048ad;
      9935: inst = 32'h8220000;
      9936: inst = 32'h10408000;
      9937: inst = 32'hc4048ae;
      9938: inst = 32'h8220000;
      9939: inst = 32'h10408000;
      9940: inst = 32'hc4048af;
      9941: inst = 32'h8220000;
      9942: inst = 32'h10408000;
      9943: inst = 32'hc4048b0;
      9944: inst = 32'h8220000;
      9945: inst = 32'h10408000;
      9946: inst = 32'hc4048b1;
      9947: inst = 32'h8220000;
      9948: inst = 32'h10408000;
      9949: inst = 32'hc4048b2;
      9950: inst = 32'h8220000;
      9951: inst = 32'h10408000;
      9952: inst = 32'hc4048b3;
      9953: inst = 32'h8220000;
      9954: inst = 32'h10408000;
      9955: inst = 32'hc4048b4;
      9956: inst = 32'h8220000;
      9957: inst = 32'h10408000;
      9958: inst = 32'hc4048b5;
      9959: inst = 32'h8220000;
      9960: inst = 32'h10408000;
      9961: inst = 32'hc4048b6;
      9962: inst = 32'h8220000;
      9963: inst = 32'h10408000;
      9964: inst = 32'hc4048b7;
      9965: inst = 32'h8220000;
      9966: inst = 32'h10408000;
      9967: inst = 32'hc4048b8;
      9968: inst = 32'h8220000;
      9969: inst = 32'h10408000;
      9970: inst = 32'hc4048b9;
      9971: inst = 32'h8220000;
      9972: inst = 32'h10408000;
      9973: inst = 32'hc4048ba;
      9974: inst = 32'h8220000;
      9975: inst = 32'h10408000;
      9976: inst = 32'hc4048bb;
      9977: inst = 32'h8220000;
      9978: inst = 32'h10408000;
      9979: inst = 32'hc4048bc;
      9980: inst = 32'h8220000;
      9981: inst = 32'h10408000;
      9982: inst = 32'hc4048bd;
      9983: inst = 32'h8220000;
      9984: inst = 32'h10408000;
      9985: inst = 32'hc4048be;
      9986: inst = 32'h8220000;
      9987: inst = 32'h10408000;
      9988: inst = 32'hc4048bf;
      9989: inst = 32'h8220000;
      9990: inst = 32'h10408000;
      9991: inst = 32'hc4048c0;
      9992: inst = 32'h8220000;
      9993: inst = 32'h10408000;
      9994: inst = 32'hc4048c1;
      9995: inst = 32'h8220000;
      9996: inst = 32'h10408000;
      9997: inst = 32'hc4048c2;
      9998: inst = 32'h8220000;
      9999: inst = 32'h10408000;
      10000: inst = 32'hc4048c3;
      10001: inst = 32'h8220000;
      10002: inst = 32'h10408000;
      10003: inst = 32'hc4048fc;
      10004: inst = 32'h8220000;
      10005: inst = 32'h10408000;
      10006: inst = 32'hc4048fd;
      10007: inst = 32'h8220000;
      10008: inst = 32'h10408000;
      10009: inst = 32'hc4048fe;
      10010: inst = 32'h8220000;
      10011: inst = 32'h10408000;
      10012: inst = 32'hc4048ff;
      10013: inst = 32'h8220000;
      10014: inst = 32'h10408000;
      10015: inst = 32'hc404900;
      10016: inst = 32'h8220000;
      10017: inst = 32'h10408000;
      10018: inst = 32'hc404901;
      10019: inst = 32'h8220000;
      10020: inst = 32'h10408000;
      10021: inst = 32'hc404902;
      10022: inst = 32'h8220000;
      10023: inst = 32'h10408000;
      10024: inst = 32'hc404903;
      10025: inst = 32'h8220000;
      10026: inst = 32'h10408000;
      10027: inst = 32'hc404904;
      10028: inst = 32'h8220000;
      10029: inst = 32'h10408000;
      10030: inst = 32'hc404905;
      10031: inst = 32'h8220000;
      10032: inst = 32'h10408000;
      10033: inst = 32'hc404906;
      10034: inst = 32'h8220000;
      10035: inst = 32'h10408000;
      10036: inst = 32'hc404907;
      10037: inst = 32'h8220000;
      10038: inst = 32'h10408000;
      10039: inst = 32'hc404908;
      10040: inst = 32'h8220000;
      10041: inst = 32'h10408000;
      10042: inst = 32'hc404909;
      10043: inst = 32'h8220000;
      10044: inst = 32'h10408000;
      10045: inst = 32'hc40490a;
      10046: inst = 32'h8220000;
      10047: inst = 32'h10408000;
      10048: inst = 32'hc40490b;
      10049: inst = 32'h8220000;
      10050: inst = 32'h10408000;
      10051: inst = 32'hc40490c;
      10052: inst = 32'h8220000;
      10053: inst = 32'h10408000;
      10054: inst = 32'hc40490d;
      10055: inst = 32'h8220000;
      10056: inst = 32'h10408000;
      10057: inst = 32'hc40490e;
      10058: inst = 32'h8220000;
      10059: inst = 32'h10408000;
      10060: inst = 32'hc40490f;
      10061: inst = 32'h8220000;
      10062: inst = 32'h10408000;
      10063: inst = 32'hc404910;
      10064: inst = 32'h8220000;
      10065: inst = 32'h10408000;
      10066: inst = 32'hc404911;
      10067: inst = 32'h8220000;
      10068: inst = 32'h10408000;
      10069: inst = 32'hc404912;
      10070: inst = 32'h8220000;
      10071: inst = 32'h10408000;
      10072: inst = 32'hc404913;
      10073: inst = 32'h8220000;
      10074: inst = 32'h10408000;
      10075: inst = 32'hc404914;
      10076: inst = 32'h8220000;
      10077: inst = 32'h10408000;
      10078: inst = 32'hc404915;
      10079: inst = 32'h8220000;
      10080: inst = 32'h10408000;
      10081: inst = 32'hc404916;
      10082: inst = 32'h8220000;
      10083: inst = 32'h10408000;
      10084: inst = 32'hc404917;
      10085: inst = 32'h8220000;
      10086: inst = 32'h10408000;
      10087: inst = 32'hc404918;
      10088: inst = 32'h8220000;
      10089: inst = 32'h10408000;
      10090: inst = 32'hc404919;
      10091: inst = 32'h8220000;
      10092: inst = 32'h10408000;
      10093: inst = 32'hc40491a;
      10094: inst = 32'h8220000;
      10095: inst = 32'h10408000;
      10096: inst = 32'hc40491b;
      10097: inst = 32'h8220000;
      10098: inst = 32'h10408000;
      10099: inst = 32'hc40491c;
      10100: inst = 32'h8220000;
      10101: inst = 32'h10408000;
      10102: inst = 32'hc40491d;
      10103: inst = 32'h8220000;
      10104: inst = 32'h10408000;
      10105: inst = 32'hc40491e;
      10106: inst = 32'h8220000;
      10107: inst = 32'h10408000;
      10108: inst = 32'hc40491f;
      10109: inst = 32'h8220000;
      10110: inst = 32'h10408000;
      10111: inst = 32'hc404920;
      10112: inst = 32'h8220000;
      10113: inst = 32'h10408000;
      10114: inst = 32'hc404921;
      10115: inst = 32'h8220000;
      10116: inst = 32'h10408000;
      10117: inst = 32'hc404922;
      10118: inst = 32'h8220000;
      10119: inst = 32'h10408000;
      10120: inst = 32'hc404923;
      10121: inst = 32'h8220000;
      10122: inst = 32'h10408000;
      10123: inst = 32'hc40495c;
      10124: inst = 32'h8220000;
      10125: inst = 32'h10408000;
      10126: inst = 32'hc40495d;
      10127: inst = 32'h8220000;
      10128: inst = 32'h10408000;
      10129: inst = 32'hc40495e;
      10130: inst = 32'h8220000;
      10131: inst = 32'h10408000;
      10132: inst = 32'hc40495f;
      10133: inst = 32'h8220000;
      10134: inst = 32'h10408000;
      10135: inst = 32'hc404960;
      10136: inst = 32'h8220000;
      10137: inst = 32'h10408000;
      10138: inst = 32'hc404961;
      10139: inst = 32'h8220000;
      10140: inst = 32'h10408000;
      10141: inst = 32'hc404962;
      10142: inst = 32'h8220000;
      10143: inst = 32'h10408000;
      10144: inst = 32'hc404963;
      10145: inst = 32'h8220000;
      10146: inst = 32'h10408000;
      10147: inst = 32'hc404964;
      10148: inst = 32'h8220000;
      10149: inst = 32'h10408000;
      10150: inst = 32'hc404965;
      10151: inst = 32'h8220000;
      10152: inst = 32'h10408000;
      10153: inst = 32'hc404966;
      10154: inst = 32'h8220000;
      10155: inst = 32'h10408000;
      10156: inst = 32'hc404967;
      10157: inst = 32'h8220000;
      10158: inst = 32'h10408000;
      10159: inst = 32'hc404968;
      10160: inst = 32'h8220000;
      10161: inst = 32'h10408000;
      10162: inst = 32'hc404969;
      10163: inst = 32'h8220000;
      10164: inst = 32'h10408000;
      10165: inst = 32'hc40496a;
      10166: inst = 32'h8220000;
      10167: inst = 32'h10408000;
      10168: inst = 32'hc40496b;
      10169: inst = 32'h8220000;
      10170: inst = 32'h10408000;
      10171: inst = 32'hc40496c;
      10172: inst = 32'h8220000;
      10173: inst = 32'h10408000;
      10174: inst = 32'hc40496d;
      10175: inst = 32'h8220000;
      10176: inst = 32'h10408000;
      10177: inst = 32'hc40496e;
      10178: inst = 32'h8220000;
      10179: inst = 32'h10408000;
      10180: inst = 32'hc40496f;
      10181: inst = 32'h8220000;
      10182: inst = 32'h10408000;
      10183: inst = 32'hc404970;
      10184: inst = 32'h8220000;
      10185: inst = 32'h10408000;
      10186: inst = 32'hc404971;
      10187: inst = 32'h8220000;
      10188: inst = 32'h10408000;
      10189: inst = 32'hc404972;
      10190: inst = 32'h8220000;
      10191: inst = 32'h10408000;
      10192: inst = 32'hc404973;
      10193: inst = 32'h8220000;
      10194: inst = 32'h10408000;
      10195: inst = 32'hc404974;
      10196: inst = 32'h8220000;
      10197: inst = 32'h10408000;
      10198: inst = 32'hc404975;
      10199: inst = 32'h8220000;
      10200: inst = 32'h10408000;
      10201: inst = 32'hc404976;
      10202: inst = 32'h8220000;
      10203: inst = 32'h10408000;
      10204: inst = 32'hc404977;
      10205: inst = 32'h8220000;
      10206: inst = 32'h10408000;
      10207: inst = 32'hc404978;
      10208: inst = 32'h8220000;
      10209: inst = 32'h10408000;
      10210: inst = 32'hc404979;
      10211: inst = 32'h8220000;
      10212: inst = 32'h10408000;
      10213: inst = 32'hc40497a;
      10214: inst = 32'h8220000;
      10215: inst = 32'h10408000;
      10216: inst = 32'hc40497b;
      10217: inst = 32'h8220000;
      10218: inst = 32'h10408000;
      10219: inst = 32'hc40497c;
      10220: inst = 32'h8220000;
      10221: inst = 32'h10408000;
      10222: inst = 32'hc40497d;
      10223: inst = 32'h8220000;
      10224: inst = 32'h10408000;
      10225: inst = 32'hc40497e;
      10226: inst = 32'h8220000;
      10227: inst = 32'h10408000;
      10228: inst = 32'hc40497f;
      10229: inst = 32'h8220000;
      10230: inst = 32'h10408000;
      10231: inst = 32'hc404980;
      10232: inst = 32'h8220000;
      10233: inst = 32'h10408000;
      10234: inst = 32'hc404981;
      10235: inst = 32'h8220000;
      10236: inst = 32'h10408000;
      10237: inst = 32'hc404982;
      10238: inst = 32'h8220000;
      10239: inst = 32'h10408000;
      10240: inst = 32'hc404983;
      10241: inst = 32'h8220000;
      10242: inst = 32'h10408000;
      10243: inst = 32'hc404992;
      10244: inst = 32'h8220000;
      10245: inst = 32'h10408000;
      10246: inst = 32'hc4049bc;
      10247: inst = 32'h8220000;
      10248: inst = 32'h10408000;
      10249: inst = 32'hc4049bd;
      10250: inst = 32'h8220000;
      10251: inst = 32'h10408000;
      10252: inst = 32'hc4049be;
      10253: inst = 32'h8220000;
      10254: inst = 32'h10408000;
      10255: inst = 32'hc4049bf;
      10256: inst = 32'h8220000;
      10257: inst = 32'h10408000;
      10258: inst = 32'hc4049c0;
      10259: inst = 32'h8220000;
      10260: inst = 32'h10408000;
      10261: inst = 32'hc4049c1;
      10262: inst = 32'h8220000;
      10263: inst = 32'h10408000;
      10264: inst = 32'hc4049c2;
      10265: inst = 32'h8220000;
      10266: inst = 32'h10408000;
      10267: inst = 32'hc4049c3;
      10268: inst = 32'h8220000;
      10269: inst = 32'h10408000;
      10270: inst = 32'hc4049c4;
      10271: inst = 32'h8220000;
      10272: inst = 32'h10408000;
      10273: inst = 32'hc4049c5;
      10274: inst = 32'h8220000;
      10275: inst = 32'h10408000;
      10276: inst = 32'hc4049c6;
      10277: inst = 32'h8220000;
      10278: inst = 32'h10408000;
      10279: inst = 32'hc4049c7;
      10280: inst = 32'h8220000;
      10281: inst = 32'h10408000;
      10282: inst = 32'hc4049c8;
      10283: inst = 32'h8220000;
      10284: inst = 32'h10408000;
      10285: inst = 32'hc4049c9;
      10286: inst = 32'h8220000;
      10287: inst = 32'h10408000;
      10288: inst = 32'hc4049ca;
      10289: inst = 32'h8220000;
      10290: inst = 32'h10408000;
      10291: inst = 32'hc4049cb;
      10292: inst = 32'h8220000;
      10293: inst = 32'h10408000;
      10294: inst = 32'hc4049cc;
      10295: inst = 32'h8220000;
      10296: inst = 32'h10408000;
      10297: inst = 32'hc4049cd;
      10298: inst = 32'h8220000;
      10299: inst = 32'h10408000;
      10300: inst = 32'hc4049ce;
      10301: inst = 32'h8220000;
      10302: inst = 32'h10408000;
      10303: inst = 32'hc4049cf;
      10304: inst = 32'h8220000;
      10305: inst = 32'h10408000;
      10306: inst = 32'hc4049d0;
      10307: inst = 32'h8220000;
      10308: inst = 32'h10408000;
      10309: inst = 32'hc4049d1;
      10310: inst = 32'h8220000;
      10311: inst = 32'h10408000;
      10312: inst = 32'hc4049d2;
      10313: inst = 32'h8220000;
      10314: inst = 32'h10408000;
      10315: inst = 32'hc4049d3;
      10316: inst = 32'h8220000;
      10317: inst = 32'h10408000;
      10318: inst = 32'hc4049d4;
      10319: inst = 32'h8220000;
      10320: inst = 32'h10408000;
      10321: inst = 32'hc4049d5;
      10322: inst = 32'h8220000;
      10323: inst = 32'h10408000;
      10324: inst = 32'hc4049d6;
      10325: inst = 32'h8220000;
      10326: inst = 32'h10408000;
      10327: inst = 32'hc4049d7;
      10328: inst = 32'h8220000;
      10329: inst = 32'h10408000;
      10330: inst = 32'hc4049d8;
      10331: inst = 32'h8220000;
      10332: inst = 32'h10408000;
      10333: inst = 32'hc4049d9;
      10334: inst = 32'h8220000;
      10335: inst = 32'h10408000;
      10336: inst = 32'hc4049da;
      10337: inst = 32'h8220000;
      10338: inst = 32'h10408000;
      10339: inst = 32'hc4049db;
      10340: inst = 32'h8220000;
      10341: inst = 32'h10408000;
      10342: inst = 32'hc4049dc;
      10343: inst = 32'h8220000;
      10344: inst = 32'h10408000;
      10345: inst = 32'hc4049dd;
      10346: inst = 32'h8220000;
      10347: inst = 32'h10408000;
      10348: inst = 32'hc4049de;
      10349: inst = 32'h8220000;
      10350: inst = 32'h10408000;
      10351: inst = 32'hc4049df;
      10352: inst = 32'h8220000;
      10353: inst = 32'h10408000;
      10354: inst = 32'hc4049e0;
      10355: inst = 32'h8220000;
      10356: inst = 32'h10408000;
      10357: inst = 32'hc4049e1;
      10358: inst = 32'h8220000;
      10359: inst = 32'h10408000;
      10360: inst = 32'hc4049e2;
      10361: inst = 32'h8220000;
      10362: inst = 32'h10408000;
      10363: inst = 32'hc4049e3;
      10364: inst = 32'h8220000;
      10365: inst = 32'h10408000;
      10366: inst = 32'hc4049f2;
      10367: inst = 32'h8220000;
      10368: inst = 32'h10408000;
      10369: inst = 32'hc404a1c;
      10370: inst = 32'h8220000;
      10371: inst = 32'h10408000;
      10372: inst = 32'hc404a1d;
      10373: inst = 32'h8220000;
      10374: inst = 32'h10408000;
      10375: inst = 32'hc404a1e;
      10376: inst = 32'h8220000;
      10377: inst = 32'h10408000;
      10378: inst = 32'hc404a1f;
      10379: inst = 32'h8220000;
      10380: inst = 32'h10408000;
      10381: inst = 32'hc404a20;
      10382: inst = 32'h8220000;
      10383: inst = 32'h10408000;
      10384: inst = 32'hc404a21;
      10385: inst = 32'h8220000;
      10386: inst = 32'h10408000;
      10387: inst = 32'hc404a22;
      10388: inst = 32'h8220000;
      10389: inst = 32'h10408000;
      10390: inst = 32'hc404a23;
      10391: inst = 32'h8220000;
      10392: inst = 32'h10408000;
      10393: inst = 32'hc404a24;
      10394: inst = 32'h8220000;
      10395: inst = 32'h10408000;
      10396: inst = 32'hc404a25;
      10397: inst = 32'h8220000;
      10398: inst = 32'h10408000;
      10399: inst = 32'hc404a26;
      10400: inst = 32'h8220000;
      10401: inst = 32'h10408000;
      10402: inst = 32'hc404a27;
      10403: inst = 32'h8220000;
      10404: inst = 32'h10408000;
      10405: inst = 32'hc404a28;
      10406: inst = 32'h8220000;
      10407: inst = 32'h10408000;
      10408: inst = 32'hc404a29;
      10409: inst = 32'h8220000;
      10410: inst = 32'h10408000;
      10411: inst = 32'hc404a2a;
      10412: inst = 32'h8220000;
      10413: inst = 32'h10408000;
      10414: inst = 32'hc404a2b;
      10415: inst = 32'h8220000;
      10416: inst = 32'h10408000;
      10417: inst = 32'hc404a2c;
      10418: inst = 32'h8220000;
      10419: inst = 32'h10408000;
      10420: inst = 32'hc404a2d;
      10421: inst = 32'h8220000;
      10422: inst = 32'h10408000;
      10423: inst = 32'hc404a2e;
      10424: inst = 32'h8220000;
      10425: inst = 32'h10408000;
      10426: inst = 32'hc404a2f;
      10427: inst = 32'h8220000;
      10428: inst = 32'h10408000;
      10429: inst = 32'hc404a30;
      10430: inst = 32'h8220000;
      10431: inst = 32'h10408000;
      10432: inst = 32'hc404a31;
      10433: inst = 32'h8220000;
      10434: inst = 32'h10408000;
      10435: inst = 32'hc404a32;
      10436: inst = 32'h8220000;
      10437: inst = 32'h10408000;
      10438: inst = 32'hc404a33;
      10439: inst = 32'h8220000;
      10440: inst = 32'h10408000;
      10441: inst = 32'hc404a34;
      10442: inst = 32'h8220000;
      10443: inst = 32'h10408000;
      10444: inst = 32'hc404a35;
      10445: inst = 32'h8220000;
      10446: inst = 32'h10408000;
      10447: inst = 32'hc404a36;
      10448: inst = 32'h8220000;
      10449: inst = 32'h10408000;
      10450: inst = 32'hc404a37;
      10451: inst = 32'h8220000;
      10452: inst = 32'h10408000;
      10453: inst = 32'hc404a38;
      10454: inst = 32'h8220000;
      10455: inst = 32'h10408000;
      10456: inst = 32'hc404a39;
      10457: inst = 32'h8220000;
      10458: inst = 32'h10408000;
      10459: inst = 32'hc404a3a;
      10460: inst = 32'h8220000;
      10461: inst = 32'h10408000;
      10462: inst = 32'hc404a3b;
      10463: inst = 32'h8220000;
      10464: inst = 32'h10408000;
      10465: inst = 32'hc404a3c;
      10466: inst = 32'h8220000;
      10467: inst = 32'h10408000;
      10468: inst = 32'hc404a3d;
      10469: inst = 32'h8220000;
      10470: inst = 32'h10408000;
      10471: inst = 32'hc404a3e;
      10472: inst = 32'h8220000;
      10473: inst = 32'h10408000;
      10474: inst = 32'hc404a3f;
      10475: inst = 32'h8220000;
      10476: inst = 32'h10408000;
      10477: inst = 32'hc404a40;
      10478: inst = 32'h8220000;
      10479: inst = 32'h10408000;
      10480: inst = 32'hc404a41;
      10481: inst = 32'h8220000;
      10482: inst = 32'h10408000;
      10483: inst = 32'hc404a42;
      10484: inst = 32'h8220000;
      10485: inst = 32'h10408000;
      10486: inst = 32'hc404a43;
      10487: inst = 32'h8220000;
      10488: inst = 32'h10408000;
      10489: inst = 32'hc404a52;
      10490: inst = 32'h8220000;
      10491: inst = 32'h10408000;
      10492: inst = 32'hc404a7c;
      10493: inst = 32'h8220000;
      10494: inst = 32'h10408000;
      10495: inst = 32'hc404a7d;
      10496: inst = 32'h8220000;
      10497: inst = 32'h10408000;
      10498: inst = 32'hc404a7e;
      10499: inst = 32'h8220000;
      10500: inst = 32'h10408000;
      10501: inst = 32'hc404a7f;
      10502: inst = 32'h8220000;
      10503: inst = 32'h10408000;
      10504: inst = 32'hc404a80;
      10505: inst = 32'h8220000;
      10506: inst = 32'h10408000;
      10507: inst = 32'hc404a81;
      10508: inst = 32'h8220000;
      10509: inst = 32'h10408000;
      10510: inst = 32'hc404a82;
      10511: inst = 32'h8220000;
      10512: inst = 32'h10408000;
      10513: inst = 32'hc404a83;
      10514: inst = 32'h8220000;
      10515: inst = 32'h10408000;
      10516: inst = 32'hc404a84;
      10517: inst = 32'h8220000;
      10518: inst = 32'h10408000;
      10519: inst = 32'hc404a85;
      10520: inst = 32'h8220000;
      10521: inst = 32'h10408000;
      10522: inst = 32'hc404a86;
      10523: inst = 32'h8220000;
      10524: inst = 32'h10408000;
      10525: inst = 32'hc404a87;
      10526: inst = 32'h8220000;
      10527: inst = 32'h10408000;
      10528: inst = 32'hc404a88;
      10529: inst = 32'h8220000;
      10530: inst = 32'h10408000;
      10531: inst = 32'hc404a89;
      10532: inst = 32'h8220000;
      10533: inst = 32'h10408000;
      10534: inst = 32'hc404a8a;
      10535: inst = 32'h8220000;
      10536: inst = 32'h10408000;
      10537: inst = 32'hc404a8b;
      10538: inst = 32'h8220000;
      10539: inst = 32'h10408000;
      10540: inst = 32'hc404a8c;
      10541: inst = 32'h8220000;
      10542: inst = 32'h10408000;
      10543: inst = 32'hc404a8d;
      10544: inst = 32'h8220000;
      10545: inst = 32'h10408000;
      10546: inst = 32'hc404a8e;
      10547: inst = 32'h8220000;
      10548: inst = 32'h10408000;
      10549: inst = 32'hc404a8f;
      10550: inst = 32'h8220000;
      10551: inst = 32'h10408000;
      10552: inst = 32'hc404a90;
      10553: inst = 32'h8220000;
      10554: inst = 32'h10408000;
      10555: inst = 32'hc404a91;
      10556: inst = 32'h8220000;
      10557: inst = 32'h10408000;
      10558: inst = 32'hc404a92;
      10559: inst = 32'h8220000;
      10560: inst = 32'h10408000;
      10561: inst = 32'hc404a93;
      10562: inst = 32'h8220000;
      10563: inst = 32'h10408000;
      10564: inst = 32'hc404a94;
      10565: inst = 32'h8220000;
      10566: inst = 32'h10408000;
      10567: inst = 32'hc404a95;
      10568: inst = 32'h8220000;
      10569: inst = 32'h10408000;
      10570: inst = 32'hc404a96;
      10571: inst = 32'h8220000;
      10572: inst = 32'h10408000;
      10573: inst = 32'hc404a97;
      10574: inst = 32'h8220000;
      10575: inst = 32'h10408000;
      10576: inst = 32'hc404a98;
      10577: inst = 32'h8220000;
      10578: inst = 32'h10408000;
      10579: inst = 32'hc404a99;
      10580: inst = 32'h8220000;
      10581: inst = 32'h10408000;
      10582: inst = 32'hc404a9a;
      10583: inst = 32'h8220000;
      10584: inst = 32'h10408000;
      10585: inst = 32'hc404a9b;
      10586: inst = 32'h8220000;
      10587: inst = 32'h10408000;
      10588: inst = 32'hc404a9c;
      10589: inst = 32'h8220000;
      10590: inst = 32'h10408000;
      10591: inst = 32'hc404a9d;
      10592: inst = 32'h8220000;
      10593: inst = 32'h10408000;
      10594: inst = 32'hc404a9e;
      10595: inst = 32'h8220000;
      10596: inst = 32'h10408000;
      10597: inst = 32'hc404a9f;
      10598: inst = 32'h8220000;
      10599: inst = 32'h10408000;
      10600: inst = 32'hc404aa0;
      10601: inst = 32'h8220000;
      10602: inst = 32'h10408000;
      10603: inst = 32'hc404aa1;
      10604: inst = 32'h8220000;
      10605: inst = 32'h10408000;
      10606: inst = 32'hc404aa2;
      10607: inst = 32'h8220000;
      10608: inst = 32'h10408000;
      10609: inst = 32'hc404aa3;
      10610: inst = 32'h8220000;
      10611: inst = 32'h10408000;
      10612: inst = 32'hc404ab4;
      10613: inst = 32'h8220000;
      10614: inst = 32'h10408000;
      10615: inst = 32'hc404adc;
      10616: inst = 32'h8220000;
      10617: inst = 32'h10408000;
      10618: inst = 32'hc404add;
      10619: inst = 32'h8220000;
      10620: inst = 32'h10408000;
      10621: inst = 32'hc404ade;
      10622: inst = 32'h8220000;
      10623: inst = 32'h10408000;
      10624: inst = 32'hc404adf;
      10625: inst = 32'h8220000;
      10626: inst = 32'h10408000;
      10627: inst = 32'hc404ae0;
      10628: inst = 32'h8220000;
      10629: inst = 32'h10408000;
      10630: inst = 32'hc404ae1;
      10631: inst = 32'h8220000;
      10632: inst = 32'h10408000;
      10633: inst = 32'hc404ae2;
      10634: inst = 32'h8220000;
      10635: inst = 32'h10408000;
      10636: inst = 32'hc404ae3;
      10637: inst = 32'h8220000;
      10638: inst = 32'h10408000;
      10639: inst = 32'hc404ae4;
      10640: inst = 32'h8220000;
      10641: inst = 32'h10408000;
      10642: inst = 32'hc404ae5;
      10643: inst = 32'h8220000;
      10644: inst = 32'h10408000;
      10645: inst = 32'hc404ae6;
      10646: inst = 32'h8220000;
      10647: inst = 32'h10408000;
      10648: inst = 32'hc404ae7;
      10649: inst = 32'h8220000;
      10650: inst = 32'h10408000;
      10651: inst = 32'hc404ae8;
      10652: inst = 32'h8220000;
      10653: inst = 32'h10408000;
      10654: inst = 32'hc404ae9;
      10655: inst = 32'h8220000;
      10656: inst = 32'h10408000;
      10657: inst = 32'hc404aea;
      10658: inst = 32'h8220000;
      10659: inst = 32'h10408000;
      10660: inst = 32'hc404aeb;
      10661: inst = 32'h8220000;
      10662: inst = 32'h10408000;
      10663: inst = 32'hc404aec;
      10664: inst = 32'h8220000;
      10665: inst = 32'h10408000;
      10666: inst = 32'hc404aed;
      10667: inst = 32'h8220000;
      10668: inst = 32'h10408000;
      10669: inst = 32'hc404aee;
      10670: inst = 32'h8220000;
      10671: inst = 32'h10408000;
      10672: inst = 32'hc404aef;
      10673: inst = 32'h8220000;
      10674: inst = 32'h10408000;
      10675: inst = 32'hc404af0;
      10676: inst = 32'h8220000;
      10677: inst = 32'h10408000;
      10678: inst = 32'hc404af1;
      10679: inst = 32'h8220000;
      10680: inst = 32'h10408000;
      10681: inst = 32'hc404af2;
      10682: inst = 32'h8220000;
      10683: inst = 32'h10408000;
      10684: inst = 32'hc404af3;
      10685: inst = 32'h8220000;
      10686: inst = 32'h10408000;
      10687: inst = 32'hc404af4;
      10688: inst = 32'h8220000;
      10689: inst = 32'h10408000;
      10690: inst = 32'hc404af5;
      10691: inst = 32'h8220000;
      10692: inst = 32'h10408000;
      10693: inst = 32'hc404af6;
      10694: inst = 32'h8220000;
      10695: inst = 32'h10408000;
      10696: inst = 32'hc404af7;
      10697: inst = 32'h8220000;
      10698: inst = 32'h10408000;
      10699: inst = 32'hc404af8;
      10700: inst = 32'h8220000;
      10701: inst = 32'h10408000;
      10702: inst = 32'hc404af9;
      10703: inst = 32'h8220000;
      10704: inst = 32'h10408000;
      10705: inst = 32'hc404afa;
      10706: inst = 32'h8220000;
      10707: inst = 32'h10408000;
      10708: inst = 32'hc404afb;
      10709: inst = 32'h8220000;
      10710: inst = 32'h10408000;
      10711: inst = 32'hc404afc;
      10712: inst = 32'h8220000;
      10713: inst = 32'h10408000;
      10714: inst = 32'hc404afd;
      10715: inst = 32'h8220000;
      10716: inst = 32'h10408000;
      10717: inst = 32'hc404afe;
      10718: inst = 32'h8220000;
      10719: inst = 32'h10408000;
      10720: inst = 32'hc404aff;
      10721: inst = 32'h8220000;
      10722: inst = 32'h10408000;
      10723: inst = 32'hc404b00;
      10724: inst = 32'h8220000;
      10725: inst = 32'h10408000;
      10726: inst = 32'hc404b01;
      10727: inst = 32'h8220000;
      10728: inst = 32'h10408000;
      10729: inst = 32'hc404b02;
      10730: inst = 32'h8220000;
      10731: inst = 32'h10408000;
      10732: inst = 32'hc404b03;
      10733: inst = 32'h8220000;
      10734: inst = 32'h10408000;
      10735: inst = 32'hc404b14;
      10736: inst = 32'h8220000;
      10737: inst = 32'h10408000;
      10738: inst = 32'hc404b3c;
      10739: inst = 32'h8220000;
      10740: inst = 32'h10408000;
      10741: inst = 32'hc404b3d;
      10742: inst = 32'h8220000;
      10743: inst = 32'h10408000;
      10744: inst = 32'hc404b3e;
      10745: inst = 32'h8220000;
      10746: inst = 32'h10408000;
      10747: inst = 32'hc404b3f;
      10748: inst = 32'h8220000;
      10749: inst = 32'h10408000;
      10750: inst = 32'hc404b40;
      10751: inst = 32'h8220000;
      10752: inst = 32'h10408000;
      10753: inst = 32'hc404b41;
      10754: inst = 32'h8220000;
      10755: inst = 32'h10408000;
      10756: inst = 32'hc404b42;
      10757: inst = 32'h8220000;
      10758: inst = 32'h10408000;
      10759: inst = 32'hc404b43;
      10760: inst = 32'h8220000;
      10761: inst = 32'h10408000;
      10762: inst = 32'hc404b44;
      10763: inst = 32'h8220000;
      10764: inst = 32'h10408000;
      10765: inst = 32'hc404b45;
      10766: inst = 32'h8220000;
      10767: inst = 32'h10408000;
      10768: inst = 32'hc404b46;
      10769: inst = 32'h8220000;
      10770: inst = 32'h10408000;
      10771: inst = 32'hc404b47;
      10772: inst = 32'h8220000;
      10773: inst = 32'h10408000;
      10774: inst = 32'hc404b48;
      10775: inst = 32'h8220000;
      10776: inst = 32'h10408000;
      10777: inst = 32'hc404b49;
      10778: inst = 32'h8220000;
      10779: inst = 32'h10408000;
      10780: inst = 32'hc404b4a;
      10781: inst = 32'h8220000;
      10782: inst = 32'h10408000;
      10783: inst = 32'hc404b4b;
      10784: inst = 32'h8220000;
      10785: inst = 32'h10408000;
      10786: inst = 32'hc404b4c;
      10787: inst = 32'h8220000;
      10788: inst = 32'h10408000;
      10789: inst = 32'hc404b4d;
      10790: inst = 32'h8220000;
      10791: inst = 32'h10408000;
      10792: inst = 32'hc404b4e;
      10793: inst = 32'h8220000;
      10794: inst = 32'h10408000;
      10795: inst = 32'hc404b4f;
      10796: inst = 32'h8220000;
      10797: inst = 32'h10408000;
      10798: inst = 32'hc404b50;
      10799: inst = 32'h8220000;
      10800: inst = 32'h10408000;
      10801: inst = 32'hc404b51;
      10802: inst = 32'h8220000;
      10803: inst = 32'h10408000;
      10804: inst = 32'hc404b52;
      10805: inst = 32'h8220000;
      10806: inst = 32'h10408000;
      10807: inst = 32'hc404b53;
      10808: inst = 32'h8220000;
      10809: inst = 32'h10408000;
      10810: inst = 32'hc404b54;
      10811: inst = 32'h8220000;
      10812: inst = 32'h10408000;
      10813: inst = 32'hc404b55;
      10814: inst = 32'h8220000;
      10815: inst = 32'h10408000;
      10816: inst = 32'hc404b56;
      10817: inst = 32'h8220000;
      10818: inst = 32'h10408000;
      10819: inst = 32'hc404b57;
      10820: inst = 32'h8220000;
      10821: inst = 32'h10408000;
      10822: inst = 32'hc404b58;
      10823: inst = 32'h8220000;
      10824: inst = 32'h10408000;
      10825: inst = 32'hc404b59;
      10826: inst = 32'h8220000;
      10827: inst = 32'h10408000;
      10828: inst = 32'hc404b5a;
      10829: inst = 32'h8220000;
      10830: inst = 32'h10408000;
      10831: inst = 32'hc404b5b;
      10832: inst = 32'h8220000;
      10833: inst = 32'h10408000;
      10834: inst = 32'hc404b5c;
      10835: inst = 32'h8220000;
      10836: inst = 32'h10408000;
      10837: inst = 32'hc404b5d;
      10838: inst = 32'h8220000;
      10839: inst = 32'h10408000;
      10840: inst = 32'hc404b5e;
      10841: inst = 32'h8220000;
      10842: inst = 32'h10408000;
      10843: inst = 32'hc404b5f;
      10844: inst = 32'h8220000;
      10845: inst = 32'h10408000;
      10846: inst = 32'hc404b60;
      10847: inst = 32'h8220000;
      10848: inst = 32'h10408000;
      10849: inst = 32'hc404b61;
      10850: inst = 32'h8220000;
      10851: inst = 32'h10408000;
      10852: inst = 32'hc404b62;
      10853: inst = 32'h8220000;
      10854: inst = 32'h10408000;
      10855: inst = 32'hc404b63;
      10856: inst = 32'h8220000;
      10857: inst = 32'h10408000;
      10858: inst = 32'hc404b9c;
      10859: inst = 32'h8220000;
      10860: inst = 32'h10408000;
      10861: inst = 32'hc404b9d;
      10862: inst = 32'h8220000;
      10863: inst = 32'h10408000;
      10864: inst = 32'hc404b9e;
      10865: inst = 32'h8220000;
      10866: inst = 32'h10408000;
      10867: inst = 32'hc404b9f;
      10868: inst = 32'h8220000;
      10869: inst = 32'h10408000;
      10870: inst = 32'hc404ba0;
      10871: inst = 32'h8220000;
      10872: inst = 32'h10408000;
      10873: inst = 32'hc404ba1;
      10874: inst = 32'h8220000;
      10875: inst = 32'h10408000;
      10876: inst = 32'hc404ba2;
      10877: inst = 32'h8220000;
      10878: inst = 32'h10408000;
      10879: inst = 32'hc404ba3;
      10880: inst = 32'h8220000;
      10881: inst = 32'h10408000;
      10882: inst = 32'hc404ba4;
      10883: inst = 32'h8220000;
      10884: inst = 32'h10408000;
      10885: inst = 32'hc404ba5;
      10886: inst = 32'h8220000;
      10887: inst = 32'h10408000;
      10888: inst = 32'hc404ba6;
      10889: inst = 32'h8220000;
      10890: inst = 32'h10408000;
      10891: inst = 32'hc404ba7;
      10892: inst = 32'h8220000;
      10893: inst = 32'h10408000;
      10894: inst = 32'hc404ba8;
      10895: inst = 32'h8220000;
      10896: inst = 32'h10408000;
      10897: inst = 32'hc404ba9;
      10898: inst = 32'h8220000;
      10899: inst = 32'h10408000;
      10900: inst = 32'hc404baa;
      10901: inst = 32'h8220000;
      10902: inst = 32'h10408000;
      10903: inst = 32'hc404bab;
      10904: inst = 32'h8220000;
      10905: inst = 32'h10408000;
      10906: inst = 32'hc404bac;
      10907: inst = 32'h8220000;
      10908: inst = 32'h10408000;
      10909: inst = 32'hc404bad;
      10910: inst = 32'h8220000;
      10911: inst = 32'h10408000;
      10912: inst = 32'hc404bae;
      10913: inst = 32'h8220000;
      10914: inst = 32'h10408000;
      10915: inst = 32'hc404baf;
      10916: inst = 32'h8220000;
      10917: inst = 32'h10408000;
      10918: inst = 32'hc404bb0;
      10919: inst = 32'h8220000;
      10920: inst = 32'h10408000;
      10921: inst = 32'hc404bb1;
      10922: inst = 32'h8220000;
      10923: inst = 32'h10408000;
      10924: inst = 32'hc404bb2;
      10925: inst = 32'h8220000;
      10926: inst = 32'h10408000;
      10927: inst = 32'hc404bb3;
      10928: inst = 32'h8220000;
      10929: inst = 32'h10408000;
      10930: inst = 32'hc404bb4;
      10931: inst = 32'h8220000;
      10932: inst = 32'h10408000;
      10933: inst = 32'hc404bb5;
      10934: inst = 32'h8220000;
      10935: inst = 32'h10408000;
      10936: inst = 32'hc404bb6;
      10937: inst = 32'h8220000;
      10938: inst = 32'h10408000;
      10939: inst = 32'hc404bb7;
      10940: inst = 32'h8220000;
      10941: inst = 32'h10408000;
      10942: inst = 32'hc404bb8;
      10943: inst = 32'h8220000;
      10944: inst = 32'h10408000;
      10945: inst = 32'hc404bb9;
      10946: inst = 32'h8220000;
      10947: inst = 32'h10408000;
      10948: inst = 32'hc404bba;
      10949: inst = 32'h8220000;
      10950: inst = 32'h10408000;
      10951: inst = 32'hc404bbb;
      10952: inst = 32'h8220000;
      10953: inst = 32'h10408000;
      10954: inst = 32'hc404bbc;
      10955: inst = 32'h8220000;
      10956: inst = 32'h10408000;
      10957: inst = 32'hc404bbd;
      10958: inst = 32'h8220000;
      10959: inst = 32'h10408000;
      10960: inst = 32'hc404bbe;
      10961: inst = 32'h8220000;
      10962: inst = 32'h10408000;
      10963: inst = 32'hc404bbf;
      10964: inst = 32'h8220000;
      10965: inst = 32'h10408000;
      10966: inst = 32'hc404bc0;
      10967: inst = 32'h8220000;
      10968: inst = 32'h10408000;
      10969: inst = 32'hc404bc1;
      10970: inst = 32'h8220000;
      10971: inst = 32'h10408000;
      10972: inst = 32'hc404bc2;
      10973: inst = 32'h8220000;
      10974: inst = 32'h10408000;
      10975: inst = 32'hc404bc3;
      10976: inst = 32'h8220000;
      10977: inst = 32'hc20ee75;
      10978: inst = 32'h10408000;
      10979: inst = 32'hc4042ea;
      10980: inst = 32'h8220000;
      10981: inst = 32'h10408000;
      10982: inst = 32'hc4043a7;
      10983: inst = 32'h8220000;
      10984: inst = 32'hc20d42c;
      10985: inst = 32'h10408000;
      10986: inst = 32'hc4042eb;
      10987: inst = 32'h8220000;
      10988: inst = 32'h10408000;
      10989: inst = 32'hc4042ec;
      10990: inst = 32'h8220000;
      10991: inst = 32'h10408000;
      10992: inst = 32'hc4043a8;
      10993: inst = 32'h8220000;
      10994: inst = 32'hc20ee55;
      10995: inst = 32'h10408000;
      10996: inst = 32'hc4042ed;
      10997: inst = 32'h8220000;
      10998: inst = 32'h10408000;
      10999: inst = 32'hc4043b0;
      11000: inst = 32'h8220000;
      11001: inst = 32'hc20e571;
      11002: inst = 32'h10408000;
      11003: inst = 32'hc404349;
      11004: inst = 32'h8220000;
      11005: inst = 32'h10408000;
      11006: inst = 32'hc40434e;
      11007: inst = 32'h8220000;
      11008: inst = 32'h10408000;
      11009: inst = 32'hc404406;
      11010: inst = 32'h8220000;
      11011: inst = 32'h10408000;
      11012: inst = 32'hc404411;
      11013: inst = 32'h8220000;
      11014: inst = 32'hc20cb28;
      11015: inst = 32'h10408000;
      11016: inst = 32'hc40434a;
      11017: inst = 32'h8220000;
      11018: inst = 32'h10408000;
      11019: inst = 32'hc40434d;
      11020: inst = 32'h8220000;
      11021: inst = 32'h10408000;
      11022: inst = 32'hc404407;
      11023: inst = 32'h8220000;
      11024: inst = 32'h10408000;
      11025: inst = 32'hc404410;
      11026: inst = 32'h8220000;
      11027: inst = 32'hc20cac7;
      11028: inst = 32'h10408000;
      11029: inst = 32'hc40434b;
      11030: inst = 32'h8220000;
      11031: inst = 32'h10408000;
      11032: inst = 32'hc40434c;
      11033: inst = 32'h8220000;
      11034: inst = 32'h10408000;
      11035: inst = 32'hc4043a9;
      11036: inst = 32'h8220000;
      11037: inst = 32'h10408000;
      11038: inst = 32'hc4043aa;
      11039: inst = 32'h8220000;
      11040: inst = 32'h10408000;
      11041: inst = 32'hc4043ab;
      11042: inst = 32'h8220000;
      11043: inst = 32'h10408000;
      11044: inst = 32'hc4043ac;
      11045: inst = 32'h8220000;
      11046: inst = 32'h10408000;
      11047: inst = 32'hc4043ad;
      11048: inst = 32'h8220000;
      11049: inst = 32'h10408000;
      11050: inst = 32'hc4043ae;
      11051: inst = 32'h8220000;
      11052: inst = 32'h10408000;
      11053: inst = 32'hc404408;
      11054: inst = 32'h8220000;
      11055: inst = 32'h10408000;
      11056: inst = 32'hc404409;
      11057: inst = 32'h8220000;
      11058: inst = 32'h10408000;
      11059: inst = 32'hc40440a;
      11060: inst = 32'h8220000;
      11061: inst = 32'h10408000;
      11062: inst = 32'hc40440b;
      11063: inst = 32'h8220000;
      11064: inst = 32'h10408000;
      11065: inst = 32'hc40440c;
      11066: inst = 32'h8220000;
      11067: inst = 32'h10408000;
      11068: inst = 32'hc40440d;
      11069: inst = 32'h8220000;
      11070: inst = 32'h10408000;
      11071: inst = 32'hc40440e;
      11072: inst = 32'h8220000;
      11073: inst = 32'h10408000;
      11074: inst = 32'hc40440f;
      11075: inst = 32'h8220000;
      11076: inst = 32'hc20d40c;
      11077: inst = 32'h10408000;
      11078: inst = 32'hc4043af;
      11079: inst = 32'h8220000;
      11080: inst = 32'hc20ee8e;
      11081: inst = 32'h10408000;
      11082: inst = 32'hc40446a;
      11083: inst = 32'h8220000;
      11084: inst = 32'h10408000;
      11085: inst = 32'hc4044b5;
      11086: inst = 32'h8220000;
      11087: inst = 32'hc20ee48;
      11088: inst = 32'h10408000;
      11089: inst = 32'hc40446b;
      11090: inst = 32'h8220000;
      11091: inst = 32'h10408000;
      11092: inst = 32'hc40446c;
      11093: inst = 32'h8220000;
      11094: inst = 32'h10408000;
      11095: inst = 32'hc4044b3;
      11096: inst = 32'h8220000;
      11097: inst = 32'h10408000;
      11098: inst = 32'hc4044b4;
      11099: inst = 32'h8220000;
      11100: inst = 32'hc20ee90;
      11101: inst = 32'h10408000;
      11102: inst = 32'hc40446d;
      11103: inst = 32'h8220000;
      11104: inst = 32'h10408000;
      11105: inst = 32'hc4044b2;
      11106: inst = 32'h8220000;
      11107: inst = 32'hc20eeb5;
      11108: inst = 32'h10408000;
      11109: inst = 32'hc4044cb;
      11110: inst = 32'h8220000;
      11111: inst = 32'h10408000;
      11112: inst = 32'hc4044cc;
      11113: inst = 32'h8220000;
      11114: inst = 32'h10408000;
      11115: inst = 32'hc404513;
      11116: inst = 32'h8220000;
      11117: inst = 32'h10408000;
      11118: inst = 32'hc404514;
      11119: inst = 32'h8220000;
      11120: inst = 32'hc20c2e2;
      11121: inst = 32'h10408000;
      11122: inst = 32'hc4046ef;
      11123: inst = 32'h8220000;
      11124: inst = 32'h10408000;
      11125: inst = 32'hc4046f0;
      11126: inst = 32'h8220000;
      11127: inst = 32'h10408000;
      11128: inst = 32'hc4046f1;
      11129: inst = 32'h8220000;
      11130: inst = 32'h10408000;
      11131: inst = 32'hc4046f2;
      11132: inst = 32'h8220000;
      11133: inst = 32'h10408000;
      11134: inst = 32'hc4046f3;
      11135: inst = 32'h8220000;
      11136: inst = 32'h10408000;
      11137: inst = 32'hc4046f4;
      11138: inst = 32'h8220000;
      11139: inst = 32'h10408000;
      11140: inst = 32'hc4046f5;
      11141: inst = 32'h8220000;
      11142: inst = 32'h10408000;
      11143: inst = 32'hc4046f6;
      11144: inst = 32'h8220000;
      11145: inst = 32'h10408000;
      11146: inst = 32'hc4046f7;
      11147: inst = 32'h8220000;
      11148: inst = 32'h10408000;
      11149: inst = 32'hc4046f8;
      11150: inst = 32'h8220000;
      11151: inst = 32'h10408000;
      11152: inst = 32'hc4046f9;
      11153: inst = 32'h8220000;
      11154: inst = 32'h10408000;
      11155: inst = 32'hc4046fa;
      11156: inst = 32'h8220000;
      11157: inst = 32'h10408000;
      11158: inst = 32'hc4046fb;
      11159: inst = 32'h8220000;
      11160: inst = 32'h10408000;
      11161: inst = 32'hc4046fc;
      11162: inst = 32'h8220000;
      11163: inst = 32'h10408000;
      11164: inst = 32'hc4046fd;
      11165: inst = 32'h8220000;
      11166: inst = 32'h10408000;
      11167: inst = 32'hc4046fe;
      11168: inst = 32'h8220000;
      11169: inst = 32'h10408000;
      11170: inst = 32'hc4046ff;
      11171: inst = 32'h8220000;
      11172: inst = 32'h10408000;
      11173: inst = 32'hc40474f;
      11174: inst = 32'h8220000;
      11175: inst = 32'h10408000;
      11176: inst = 32'hc40475f;
      11177: inst = 32'h8220000;
      11178: inst = 32'h10408000;
      11179: inst = 32'hc4047af;
      11180: inst = 32'h8220000;
      11181: inst = 32'h10408000;
      11182: inst = 32'hc4047bf;
      11183: inst = 32'h8220000;
      11184: inst = 32'h10408000;
      11185: inst = 32'hc40480f;
      11186: inst = 32'h8220000;
      11187: inst = 32'h10408000;
      11188: inst = 32'hc40481f;
      11189: inst = 32'h8220000;
      11190: inst = 32'h10408000;
      11191: inst = 32'hc40486f;
      11192: inst = 32'h8220000;
      11193: inst = 32'h10408000;
      11194: inst = 32'hc40487f;
      11195: inst = 32'h8220000;
      11196: inst = 32'h10408000;
      11197: inst = 32'hc4048cf;
      11198: inst = 32'h8220000;
      11199: inst = 32'h10408000;
      11200: inst = 32'hc4048df;
      11201: inst = 32'h8220000;
      11202: inst = 32'h10408000;
      11203: inst = 32'hc40492f;
      11204: inst = 32'h8220000;
      11205: inst = 32'h10408000;
      11206: inst = 32'hc40493f;
      11207: inst = 32'h8220000;
      11208: inst = 32'h10408000;
      11209: inst = 32'hc40498f;
      11210: inst = 32'h8220000;
      11211: inst = 32'h10408000;
      11212: inst = 32'hc40499f;
      11213: inst = 32'h8220000;
      11214: inst = 32'h10408000;
      11215: inst = 32'hc4049ef;
      11216: inst = 32'h8220000;
      11217: inst = 32'h10408000;
      11218: inst = 32'hc4049ff;
      11219: inst = 32'h8220000;
      11220: inst = 32'h10408000;
      11221: inst = 32'hc404a4f;
      11222: inst = 32'h8220000;
      11223: inst = 32'h10408000;
      11224: inst = 32'hc404a5f;
      11225: inst = 32'h8220000;
      11226: inst = 32'h10408000;
      11227: inst = 32'hc404aaf;
      11228: inst = 32'h8220000;
      11229: inst = 32'h10408000;
      11230: inst = 32'hc404abf;
      11231: inst = 32'h8220000;
      11232: inst = 32'h10408000;
      11233: inst = 32'hc404b0f;
      11234: inst = 32'h8220000;
      11235: inst = 32'h10408000;
      11236: inst = 32'hc404b1f;
      11237: inst = 32'h8220000;
      11238: inst = 32'h10408000;
      11239: inst = 32'hc404b6f;
      11240: inst = 32'h8220000;
      11241: inst = 32'h10408000;
      11242: inst = 32'hc404b7f;
      11243: inst = 32'h8220000;
      11244: inst = 32'h10408000;
      11245: inst = 32'hc404bcf;
      11246: inst = 32'h8220000;
      11247: inst = 32'h10408000;
      11248: inst = 32'hc404bdf;
      11249: inst = 32'h8220000;
      11250: inst = 32'h10408000;
      11251: inst = 32'hc404c2f;
      11252: inst = 32'h8220000;
      11253: inst = 32'h10408000;
      11254: inst = 32'hc404c3f;
      11255: inst = 32'h8220000;
      11256: inst = 32'h10408000;
      11257: inst = 32'hc404c8f;
      11258: inst = 32'h8220000;
      11259: inst = 32'h10408000;
      11260: inst = 32'hc404c9f;
      11261: inst = 32'h8220000;
      11262: inst = 32'h10408000;
      11263: inst = 32'hc404cef;
      11264: inst = 32'h8220000;
      11265: inst = 32'h10408000;
      11266: inst = 32'hc404cff;
      11267: inst = 32'h8220000;
      11268: inst = 32'h10408000;
      11269: inst = 32'hc404d4f;
      11270: inst = 32'h8220000;
      11271: inst = 32'h10408000;
      11272: inst = 32'hc404d5f;
      11273: inst = 32'h8220000;
      11274: inst = 32'h10408000;
      11275: inst = 32'hc404daf;
      11276: inst = 32'h8220000;
      11277: inst = 32'h10408000;
      11278: inst = 32'hc404dbf;
      11279: inst = 32'h8220000;
      11280: inst = 32'h10408000;
      11281: inst = 32'hc404e0f;
      11282: inst = 32'h8220000;
      11283: inst = 32'h10408000;
      11284: inst = 32'hc404e1f;
      11285: inst = 32'h8220000;
      11286: inst = 32'h10408000;
      11287: inst = 32'hc404e6f;
      11288: inst = 32'h8220000;
      11289: inst = 32'h10408000;
      11290: inst = 32'hc404e7f;
      11291: inst = 32'h8220000;
      11292: inst = 32'h10408000;
      11293: inst = 32'hc404ecf;
      11294: inst = 32'h8220000;
      11295: inst = 32'h10408000;
      11296: inst = 32'hc404edf;
      11297: inst = 32'h8220000;
      11298: inst = 32'h10408000;
      11299: inst = 32'hc404f2f;
      11300: inst = 32'h8220000;
      11301: inst = 32'h10408000;
      11302: inst = 32'hc404f3f;
      11303: inst = 32'h8220000;
      11304: inst = 32'h10408000;
      11305: inst = 32'hc404f8f;
      11306: inst = 32'h8220000;
      11307: inst = 32'h10408000;
      11308: inst = 32'hc404f9f;
      11309: inst = 32'h8220000;
      11310: inst = 32'h10408000;
      11311: inst = 32'hc404fef;
      11312: inst = 32'h8220000;
      11313: inst = 32'h10408000;
      11314: inst = 32'hc404fff;
      11315: inst = 32'h8220000;
      11316: inst = 32'h10408000;
      11317: inst = 32'hc40504f;
      11318: inst = 32'h8220000;
      11319: inst = 32'h10408000;
      11320: inst = 32'hc40505f;
      11321: inst = 32'h8220000;
      11322: inst = 32'h10408000;
      11323: inst = 32'hc4050af;
      11324: inst = 32'h8220000;
      11325: inst = 32'h10408000;
      11326: inst = 32'hc4050bf;
      11327: inst = 32'h8220000;
      11328: inst = 32'h10408000;
      11329: inst = 32'hc40510f;
      11330: inst = 32'h8220000;
      11331: inst = 32'h10408000;
      11332: inst = 32'hc40511f;
      11333: inst = 32'h8220000;
      11334: inst = 32'h10408000;
      11335: inst = 32'hc40516f;
      11336: inst = 32'h8220000;
      11337: inst = 32'h10408000;
      11338: inst = 32'hc40517f;
      11339: inst = 32'h8220000;
      11340: inst = 32'h10408000;
      11341: inst = 32'hc4051cf;
      11342: inst = 32'h8220000;
      11343: inst = 32'h10408000;
      11344: inst = 32'hc4051df;
      11345: inst = 32'h8220000;
      11346: inst = 32'h10408000;
      11347: inst = 32'hc40522f;
      11348: inst = 32'h8220000;
      11349: inst = 32'h10408000;
      11350: inst = 32'hc40523f;
      11351: inst = 32'h8220000;
      11352: inst = 32'h10408000;
      11353: inst = 32'hc40528f;
      11354: inst = 32'h8220000;
      11355: inst = 32'h10408000;
      11356: inst = 32'hc40529f;
      11357: inst = 32'h8220000;
      11358: inst = 32'h10408000;
      11359: inst = 32'hc4052ef;
      11360: inst = 32'h8220000;
      11361: inst = 32'h10408000;
      11362: inst = 32'hc4052f0;
      11363: inst = 32'h8220000;
      11364: inst = 32'h10408000;
      11365: inst = 32'hc4052f1;
      11366: inst = 32'h8220000;
      11367: inst = 32'h10408000;
      11368: inst = 32'hc4052f2;
      11369: inst = 32'h8220000;
      11370: inst = 32'h10408000;
      11371: inst = 32'hc4052f3;
      11372: inst = 32'h8220000;
      11373: inst = 32'h10408000;
      11374: inst = 32'hc4052f4;
      11375: inst = 32'h8220000;
      11376: inst = 32'h10408000;
      11377: inst = 32'hc4052f5;
      11378: inst = 32'h8220000;
      11379: inst = 32'h10408000;
      11380: inst = 32'hc4052f6;
      11381: inst = 32'h8220000;
      11382: inst = 32'h10408000;
      11383: inst = 32'hc4052f7;
      11384: inst = 32'h8220000;
      11385: inst = 32'h10408000;
      11386: inst = 32'hc4052f8;
      11387: inst = 32'h8220000;
      11388: inst = 32'h10408000;
      11389: inst = 32'hc4052f9;
      11390: inst = 32'h8220000;
      11391: inst = 32'h10408000;
      11392: inst = 32'hc4052fa;
      11393: inst = 32'h8220000;
      11394: inst = 32'h10408000;
      11395: inst = 32'hc4052fb;
      11396: inst = 32'h8220000;
      11397: inst = 32'h10408000;
      11398: inst = 32'hc4052fc;
      11399: inst = 32'h8220000;
      11400: inst = 32'h10408000;
      11401: inst = 32'hc4052fd;
      11402: inst = 32'h8220000;
      11403: inst = 32'h10408000;
      11404: inst = 32'hc4052fe;
      11405: inst = 32'h8220000;
      11406: inst = 32'h10408000;
      11407: inst = 32'hc4052ff;
      11408: inst = 32'h8220000;
      11409: inst = 32'hc20dbc5;
      11410: inst = 32'h10408000;
      11411: inst = 32'hc404750;
      11412: inst = 32'h8220000;
      11413: inst = 32'h10408000;
      11414: inst = 32'hc404751;
      11415: inst = 32'h8220000;
      11416: inst = 32'h10408000;
      11417: inst = 32'hc404752;
      11418: inst = 32'h8220000;
      11419: inst = 32'h10408000;
      11420: inst = 32'hc404753;
      11421: inst = 32'h8220000;
      11422: inst = 32'h10408000;
      11423: inst = 32'hc404754;
      11424: inst = 32'h8220000;
      11425: inst = 32'h10408000;
      11426: inst = 32'hc404755;
      11427: inst = 32'h8220000;
      11428: inst = 32'h10408000;
      11429: inst = 32'hc404756;
      11430: inst = 32'h8220000;
      11431: inst = 32'h10408000;
      11432: inst = 32'hc404757;
      11433: inst = 32'h8220000;
      11434: inst = 32'h10408000;
      11435: inst = 32'hc404758;
      11436: inst = 32'h8220000;
      11437: inst = 32'h10408000;
      11438: inst = 32'hc404759;
      11439: inst = 32'h8220000;
      11440: inst = 32'h10408000;
      11441: inst = 32'hc40475a;
      11442: inst = 32'h8220000;
      11443: inst = 32'h10408000;
      11444: inst = 32'hc40475b;
      11445: inst = 32'h8220000;
      11446: inst = 32'h10408000;
      11447: inst = 32'hc40475c;
      11448: inst = 32'h8220000;
      11449: inst = 32'h10408000;
      11450: inst = 32'hc40475d;
      11451: inst = 32'h8220000;
      11452: inst = 32'h10408000;
      11453: inst = 32'hc40475e;
      11454: inst = 32'h8220000;
      11455: inst = 32'h10408000;
      11456: inst = 32'hc4047b0;
      11457: inst = 32'h8220000;
      11458: inst = 32'h10408000;
      11459: inst = 32'hc4047b1;
      11460: inst = 32'h8220000;
      11461: inst = 32'h10408000;
      11462: inst = 32'hc4047b2;
      11463: inst = 32'h8220000;
      11464: inst = 32'h10408000;
      11465: inst = 32'hc4047b3;
      11466: inst = 32'h8220000;
      11467: inst = 32'h10408000;
      11468: inst = 32'hc4047b4;
      11469: inst = 32'h8220000;
      11470: inst = 32'h10408000;
      11471: inst = 32'hc4047b5;
      11472: inst = 32'h8220000;
      11473: inst = 32'h10408000;
      11474: inst = 32'hc4047b6;
      11475: inst = 32'h8220000;
      11476: inst = 32'h10408000;
      11477: inst = 32'hc4047b7;
      11478: inst = 32'h8220000;
      11479: inst = 32'h10408000;
      11480: inst = 32'hc4047b8;
      11481: inst = 32'h8220000;
      11482: inst = 32'h10408000;
      11483: inst = 32'hc4047b9;
      11484: inst = 32'h8220000;
      11485: inst = 32'h10408000;
      11486: inst = 32'hc4047ba;
      11487: inst = 32'h8220000;
      11488: inst = 32'h10408000;
      11489: inst = 32'hc4047bb;
      11490: inst = 32'h8220000;
      11491: inst = 32'h10408000;
      11492: inst = 32'hc4047bc;
      11493: inst = 32'h8220000;
      11494: inst = 32'h10408000;
      11495: inst = 32'hc4047bd;
      11496: inst = 32'h8220000;
      11497: inst = 32'h10408000;
      11498: inst = 32'hc4047be;
      11499: inst = 32'h8220000;
      11500: inst = 32'h10408000;
      11501: inst = 32'hc404810;
      11502: inst = 32'h8220000;
      11503: inst = 32'h10408000;
      11504: inst = 32'hc404811;
      11505: inst = 32'h8220000;
      11506: inst = 32'h10408000;
      11507: inst = 32'hc404812;
      11508: inst = 32'h8220000;
      11509: inst = 32'h10408000;
      11510: inst = 32'hc404813;
      11511: inst = 32'h8220000;
      11512: inst = 32'h10408000;
      11513: inst = 32'hc404814;
      11514: inst = 32'h8220000;
      11515: inst = 32'h10408000;
      11516: inst = 32'hc404815;
      11517: inst = 32'h8220000;
      11518: inst = 32'h10408000;
      11519: inst = 32'hc404816;
      11520: inst = 32'h8220000;
      11521: inst = 32'h10408000;
      11522: inst = 32'hc404817;
      11523: inst = 32'h8220000;
      11524: inst = 32'h10408000;
      11525: inst = 32'hc404818;
      11526: inst = 32'h8220000;
      11527: inst = 32'h10408000;
      11528: inst = 32'hc404819;
      11529: inst = 32'h8220000;
      11530: inst = 32'h10408000;
      11531: inst = 32'hc40481a;
      11532: inst = 32'h8220000;
      11533: inst = 32'h10408000;
      11534: inst = 32'hc40481b;
      11535: inst = 32'h8220000;
      11536: inst = 32'h10408000;
      11537: inst = 32'hc40481c;
      11538: inst = 32'h8220000;
      11539: inst = 32'h10408000;
      11540: inst = 32'hc40481d;
      11541: inst = 32'h8220000;
      11542: inst = 32'h10408000;
      11543: inst = 32'hc40481e;
      11544: inst = 32'h8220000;
      11545: inst = 32'h10408000;
      11546: inst = 32'hc404870;
      11547: inst = 32'h8220000;
      11548: inst = 32'h10408000;
      11549: inst = 32'hc404871;
      11550: inst = 32'h8220000;
      11551: inst = 32'h10408000;
      11552: inst = 32'hc404872;
      11553: inst = 32'h8220000;
      11554: inst = 32'h10408000;
      11555: inst = 32'hc404873;
      11556: inst = 32'h8220000;
      11557: inst = 32'h10408000;
      11558: inst = 32'hc404874;
      11559: inst = 32'h8220000;
      11560: inst = 32'h10408000;
      11561: inst = 32'hc404875;
      11562: inst = 32'h8220000;
      11563: inst = 32'h10408000;
      11564: inst = 32'hc404876;
      11565: inst = 32'h8220000;
      11566: inst = 32'h10408000;
      11567: inst = 32'hc404877;
      11568: inst = 32'h8220000;
      11569: inst = 32'h10408000;
      11570: inst = 32'hc404878;
      11571: inst = 32'h8220000;
      11572: inst = 32'h10408000;
      11573: inst = 32'hc404879;
      11574: inst = 32'h8220000;
      11575: inst = 32'h10408000;
      11576: inst = 32'hc40487a;
      11577: inst = 32'h8220000;
      11578: inst = 32'h10408000;
      11579: inst = 32'hc40487b;
      11580: inst = 32'h8220000;
      11581: inst = 32'h10408000;
      11582: inst = 32'hc40487c;
      11583: inst = 32'h8220000;
      11584: inst = 32'h10408000;
      11585: inst = 32'hc40487d;
      11586: inst = 32'h8220000;
      11587: inst = 32'h10408000;
      11588: inst = 32'hc40487e;
      11589: inst = 32'h8220000;
      11590: inst = 32'h10408000;
      11591: inst = 32'hc4048d0;
      11592: inst = 32'h8220000;
      11593: inst = 32'h10408000;
      11594: inst = 32'hc4048d1;
      11595: inst = 32'h8220000;
      11596: inst = 32'h10408000;
      11597: inst = 32'hc4048d2;
      11598: inst = 32'h8220000;
      11599: inst = 32'h10408000;
      11600: inst = 32'hc4048d3;
      11601: inst = 32'h8220000;
      11602: inst = 32'h10408000;
      11603: inst = 32'hc4048d4;
      11604: inst = 32'h8220000;
      11605: inst = 32'h10408000;
      11606: inst = 32'hc4048d5;
      11607: inst = 32'h8220000;
      11608: inst = 32'h10408000;
      11609: inst = 32'hc4048d6;
      11610: inst = 32'h8220000;
      11611: inst = 32'h10408000;
      11612: inst = 32'hc4048d7;
      11613: inst = 32'h8220000;
      11614: inst = 32'h10408000;
      11615: inst = 32'hc4048d8;
      11616: inst = 32'h8220000;
      11617: inst = 32'h10408000;
      11618: inst = 32'hc4048d9;
      11619: inst = 32'h8220000;
      11620: inst = 32'h10408000;
      11621: inst = 32'hc4048da;
      11622: inst = 32'h8220000;
      11623: inst = 32'h10408000;
      11624: inst = 32'hc4048db;
      11625: inst = 32'h8220000;
      11626: inst = 32'h10408000;
      11627: inst = 32'hc4048dc;
      11628: inst = 32'h8220000;
      11629: inst = 32'h10408000;
      11630: inst = 32'hc4048dd;
      11631: inst = 32'h8220000;
      11632: inst = 32'h10408000;
      11633: inst = 32'hc4048de;
      11634: inst = 32'h8220000;
      11635: inst = 32'h10408000;
      11636: inst = 32'hc404930;
      11637: inst = 32'h8220000;
      11638: inst = 32'h10408000;
      11639: inst = 32'hc404931;
      11640: inst = 32'h8220000;
      11641: inst = 32'h10408000;
      11642: inst = 32'hc404936;
      11643: inst = 32'h8220000;
      11644: inst = 32'h10408000;
      11645: inst = 32'hc404937;
      11646: inst = 32'h8220000;
      11647: inst = 32'h10408000;
      11648: inst = 32'hc404938;
      11649: inst = 32'h8220000;
      11650: inst = 32'h10408000;
      11651: inst = 32'hc404939;
      11652: inst = 32'h8220000;
      11653: inst = 32'h10408000;
      11654: inst = 32'hc40493a;
      11655: inst = 32'h8220000;
      11656: inst = 32'h10408000;
      11657: inst = 32'hc40493b;
      11658: inst = 32'h8220000;
      11659: inst = 32'h10408000;
      11660: inst = 32'hc40493c;
      11661: inst = 32'h8220000;
      11662: inst = 32'h10408000;
      11663: inst = 32'hc40493d;
      11664: inst = 32'h8220000;
      11665: inst = 32'h10408000;
      11666: inst = 32'hc40493e;
      11667: inst = 32'h8220000;
      11668: inst = 32'h10408000;
      11669: inst = 32'hc404990;
      11670: inst = 32'h8220000;
      11671: inst = 32'h10408000;
      11672: inst = 32'hc404991;
      11673: inst = 32'h8220000;
      11674: inst = 32'h10408000;
      11675: inst = 32'hc404996;
      11676: inst = 32'h8220000;
      11677: inst = 32'h10408000;
      11678: inst = 32'hc404997;
      11679: inst = 32'h8220000;
      11680: inst = 32'h10408000;
      11681: inst = 32'hc404998;
      11682: inst = 32'h8220000;
      11683: inst = 32'h10408000;
      11684: inst = 32'hc404999;
      11685: inst = 32'h8220000;
      11686: inst = 32'h10408000;
      11687: inst = 32'hc40499a;
      11688: inst = 32'h8220000;
      11689: inst = 32'h10408000;
      11690: inst = 32'hc40499b;
      11691: inst = 32'h8220000;
      11692: inst = 32'h10408000;
      11693: inst = 32'hc40499c;
      11694: inst = 32'h8220000;
      11695: inst = 32'h10408000;
      11696: inst = 32'hc40499d;
      11697: inst = 32'h8220000;
      11698: inst = 32'h10408000;
      11699: inst = 32'hc40499e;
      11700: inst = 32'h8220000;
      11701: inst = 32'h10408000;
      11702: inst = 32'hc4049f0;
      11703: inst = 32'h8220000;
      11704: inst = 32'h10408000;
      11705: inst = 32'hc4049f1;
      11706: inst = 32'h8220000;
      11707: inst = 32'h10408000;
      11708: inst = 32'hc4049f6;
      11709: inst = 32'h8220000;
      11710: inst = 32'h10408000;
      11711: inst = 32'hc4049f7;
      11712: inst = 32'h8220000;
      11713: inst = 32'h10408000;
      11714: inst = 32'hc4049f8;
      11715: inst = 32'h8220000;
      11716: inst = 32'h10408000;
      11717: inst = 32'hc4049f9;
      11718: inst = 32'h8220000;
      11719: inst = 32'h10408000;
      11720: inst = 32'hc4049fa;
      11721: inst = 32'h8220000;
      11722: inst = 32'h10408000;
      11723: inst = 32'hc4049fb;
      11724: inst = 32'h8220000;
      11725: inst = 32'h10408000;
      11726: inst = 32'hc4049fc;
      11727: inst = 32'h8220000;
      11728: inst = 32'h10408000;
      11729: inst = 32'hc4049fd;
      11730: inst = 32'h8220000;
      11731: inst = 32'h10408000;
      11732: inst = 32'hc4049fe;
      11733: inst = 32'h8220000;
      11734: inst = 32'h10408000;
      11735: inst = 32'hc404a50;
      11736: inst = 32'h8220000;
      11737: inst = 32'h10408000;
      11738: inst = 32'hc404a51;
      11739: inst = 32'h8220000;
      11740: inst = 32'h10408000;
      11741: inst = 32'hc404a56;
      11742: inst = 32'h8220000;
      11743: inst = 32'h10408000;
      11744: inst = 32'hc404a57;
      11745: inst = 32'h8220000;
      11746: inst = 32'h10408000;
      11747: inst = 32'hc404a58;
      11748: inst = 32'h8220000;
      11749: inst = 32'h10408000;
      11750: inst = 32'hc404a59;
      11751: inst = 32'h8220000;
      11752: inst = 32'h10408000;
      11753: inst = 32'hc404a5a;
      11754: inst = 32'h8220000;
      11755: inst = 32'h10408000;
      11756: inst = 32'hc404a5b;
      11757: inst = 32'h8220000;
      11758: inst = 32'h10408000;
      11759: inst = 32'hc404a5c;
      11760: inst = 32'h8220000;
      11761: inst = 32'h10408000;
      11762: inst = 32'hc404a5d;
      11763: inst = 32'h8220000;
      11764: inst = 32'h10408000;
      11765: inst = 32'hc404a5e;
      11766: inst = 32'h8220000;
      11767: inst = 32'h10408000;
      11768: inst = 32'hc404ab0;
      11769: inst = 32'h8220000;
      11770: inst = 32'h10408000;
      11771: inst = 32'hc404ab1;
      11772: inst = 32'h8220000;
      11773: inst = 32'h10408000;
      11774: inst = 32'hc404ab6;
      11775: inst = 32'h8220000;
      11776: inst = 32'h10408000;
      11777: inst = 32'hc404ab7;
      11778: inst = 32'h8220000;
      11779: inst = 32'h10408000;
      11780: inst = 32'hc404ab8;
      11781: inst = 32'h8220000;
      11782: inst = 32'h10408000;
      11783: inst = 32'hc404ab9;
      11784: inst = 32'h8220000;
      11785: inst = 32'h10408000;
      11786: inst = 32'hc404aba;
      11787: inst = 32'h8220000;
      11788: inst = 32'h10408000;
      11789: inst = 32'hc404abb;
      11790: inst = 32'h8220000;
      11791: inst = 32'h10408000;
      11792: inst = 32'hc404abc;
      11793: inst = 32'h8220000;
      11794: inst = 32'h10408000;
      11795: inst = 32'hc404abd;
      11796: inst = 32'h8220000;
      11797: inst = 32'h10408000;
      11798: inst = 32'hc404abe;
      11799: inst = 32'h8220000;
      11800: inst = 32'h10408000;
      11801: inst = 32'hc404b10;
      11802: inst = 32'h8220000;
      11803: inst = 32'h10408000;
      11804: inst = 32'hc404b11;
      11805: inst = 32'h8220000;
      11806: inst = 32'h10408000;
      11807: inst = 32'hc404b16;
      11808: inst = 32'h8220000;
      11809: inst = 32'h10408000;
      11810: inst = 32'hc404b17;
      11811: inst = 32'h8220000;
      11812: inst = 32'h10408000;
      11813: inst = 32'hc404b18;
      11814: inst = 32'h8220000;
      11815: inst = 32'h10408000;
      11816: inst = 32'hc404b19;
      11817: inst = 32'h8220000;
      11818: inst = 32'h10408000;
      11819: inst = 32'hc404b1a;
      11820: inst = 32'h8220000;
      11821: inst = 32'h10408000;
      11822: inst = 32'hc404b1b;
      11823: inst = 32'h8220000;
      11824: inst = 32'h10408000;
      11825: inst = 32'hc404b1c;
      11826: inst = 32'h8220000;
      11827: inst = 32'h10408000;
      11828: inst = 32'hc404b1d;
      11829: inst = 32'h8220000;
      11830: inst = 32'h10408000;
      11831: inst = 32'hc404b1e;
      11832: inst = 32'h8220000;
      11833: inst = 32'h10408000;
      11834: inst = 32'hc404b70;
      11835: inst = 32'h8220000;
      11836: inst = 32'h10408000;
      11837: inst = 32'hc404b71;
      11838: inst = 32'h8220000;
      11839: inst = 32'h10408000;
      11840: inst = 32'hc404b76;
      11841: inst = 32'h8220000;
      11842: inst = 32'h10408000;
      11843: inst = 32'hc404b77;
      11844: inst = 32'h8220000;
      11845: inst = 32'h10408000;
      11846: inst = 32'hc404b78;
      11847: inst = 32'h8220000;
      11848: inst = 32'h10408000;
      11849: inst = 32'hc404b79;
      11850: inst = 32'h8220000;
      11851: inst = 32'h10408000;
      11852: inst = 32'hc404b7a;
      11853: inst = 32'h8220000;
      11854: inst = 32'h10408000;
      11855: inst = 32'hc404b7b;
      11856: inst = 32'h8220000;
      11857: inst = 32'h10408000;
      11858: inst = 32'hc404b7c;
      11859: inst = 32'h8220000;
      11860: inst = 32'h10408000;
      11861: inst = 32'hc404b7d;
      11862: inst = 32'h8220000;
      11863: inst = 32'h10408000;
      11864: inst = 32'hc404b7e;
      11865: inst = 32'h8220000;
      11866: inst = 32'h10408000;
      11867: inst = 32'hc404bd0;
      11868: inst = 32'h8220000;
      11869: inst = 32'h10408000;
      11870: inst = 32'hc404bd1;
      11871: inst = 32'h8220000;
      11872: inst = 32'h10408000;
      11873: inst = 32'hc404bd2;
      11874: inst = 32'h8220000;
      11875: inst = 32'h10408000;
      11876: inst = 32'hc404bd3;
      11877: inst = 32'h8220000;
      11878: inst = 32'h10408000;
      11879: inst = 32'hc404bd4;
      11880: inst = 32'h8220000;
      11881: inst = 32'h10408000;
      11882: inst = 32'hc404bd5;
      11883: inst = 32'h8220000;
      11884: inst = 32'h10408000;
      11885: inst = 32'hc404bd6;
      11886: inst = 32'h8220000;
      11887: inst = 32'h10408000;
      11888: inst = 32'hc404bd7;
      11889: inst = 32'h8220000;
      11890: inst = 32'h10408000;
      11891: inst = 32'hc404bd8;
      11892: inst = 32'h8220000;
      11893: inst = 32'h10408000;
      11894: inst = 32'hc404bd9;
      11895: inst = 32'h8220000;
      11896: inst = 32'h10408000;
      11897: inst = 32'hc404bda;
      11898: inst = 32'h8220000;
      11899: inst = 32'h10408000;
      11900: inst = 32'hc404bdb;
      11901: inst = 32'h8220000;
      11902: inst = 32'h10408000;
      11903: inst = 32'hc404bdc;
      11904: inst = 32'h8220000;
      11905: inst = 32'h10408000;
      11906: inst = 32'hc404bdd;
      11907: inst = 32'h8220000;
      11908: inst = 32'h10408000;
      11909: inst = 32'hc404bde;
      11910: inst = 32'h8220000;
      11911: inst = 32'h10408000;
      11912: inst = 32'hc404c30;
      11913: inst = 32'h8220000;
      11914: inst = 32'h10408000;
      11915: inst = 32'hc404c31;
      11916: inst = 32'h8220000;
      11917: inst = 32'h10408000;
      11918: inst = 32'hc404c32;
      11919: inst = 32'h8220000;
      11920: inst = 32'h10408000;
      11921: inst = 32'hc404c33;
      11922: inst = 32'h8220000;
      11923: inst = 32'h10408000;
      11924: inst = 32'hc404c34;
      11925: inst = 32'h8220000;
      11926: inst = 32'h10408000;
      11927: inst = 32'hc404c35;
      11928: inst = 32'h8220000;
      11929: inst = 32'h10408000;
      11930: inst = 32'hc404c36;
      11931: inst = 32'h8220000;
      11932: inst = 32'h10408000;
      11933: inst = 32'hc404c37;
      11934: inst = 32'h8220000;
      11935: inst = 32'h10408000;
      11936: inst = 32'hc404c38;
      11937: inst = 32'h8220000;
      11938: inst = 32'h10408000;
      11939: inst = 32'hc404c39;
      11940: inst = 32'h8220000;
      11941: inst = 32'h10408000;
      11942: inst = 32'hc404c3a;
      11943: inst = 32'h8220000;
      11944: inst = 32'h10408000;
      11945: inst = 32'hc404c3b;
      11946: inst = 32'h8220000;
      11947: inst = 32'h10408000;
      11948: inst = 32'hc404c3c;
      11949: inst = 32'h8220000;
      11950: inst = 32'h10408000;
      11951: inst = 32'hc404c3d;
      11952: inst = 32'h8220000;
      11953: inst = 32'h10408000;
      11954: inst = 32'hc404c3e;
      11955: inst = 32'h8220000;
      11956: inst = 32'h10408000;
      11957: inst = 32'hc404c90;
      11958: inst = 32'h8220000;
      11959: inst = 32'h10408000;
      11960: inst = 32'hc404c91;
      11961: inst = 32'h8220000;
      11962: inst = 32'h10408000;
      11963: inst = 32'hc404c92;
      11964: inst = 32'h8220000;
      11965: inst = 32'h10408000;
      11966: inst = 32'hc404c93;
      11967: inst = 32'h8220000;
      11968: inst = 32'h10408000;
      11969: inst = 32'hc404c94;
      11970: inst = 32'h8220000;
      11971: inst = 32'h10408000;
      11972: inst = 32'hc404c95;
      11973: inst = 32'h8220000;
      11974: inst = 32'h10408000;
      11975: inst = 32'hc404c96;
      11976: inst = 32'h8220000;
      11977: inst = 32'h10408000;
      11978: inst = 32'hc404c97;
      11979: inst = 32'h8220000;
      11980: inst = 32'h10408000;
      11981: inst = 32'hc404c98;
      11982: inst = 32'h8220000;
      11983: inst = 32'h10408000;
      11984: inst = 32'hc404c99;
      11985: inst = 32'h8220000;
      11986: inst = 32'h10408000;
      11987: inst = 32'hc404c9a;
      11988: inst = 32'h8220000;
      11989: inst = 32'h10408000;
      11990: inst = 32'hc404c9b;
      11991: inst = 32'h8220000;
      11992: inst = 32'h10408000;
      11993: inst = 32'hc404c9c;
      11994: inst = 32'h8220000;
      11995: inst = 32'h10408000;
      11996: inst = 32'hc404c9d;
      11997: inst = 32'h8220000;
      11998: inst = 32'h10408000;
      11999: inst = 32'hc404c9e;
      12000: inst = 32'h8220000;
      12001: inst = 32'h10408000;
      12002: inst = 32'hc404cf0;
      12003: inst = 32'h8220000;
      12004: inst = 32'h10408000;
      12005: inst = 32'hc404cf1;
      12006: inst = 32'h8220000;
      12007: inst = 32'h10408000;
      12008: inst = 32'hc404cf2;
      12009: inst = 32'h8220000;
      12010: inst = 32'h10408000;
      12011: inst = 32'hc404cf3;
      12012: inst = 32'h8220000;
      12013: inst = 32'h10408000;
      12014: inst = 32'hc404cf4;
      12015: inst = 32'h8220000;
      12016: inst = 32'h10408000;
      12017: inst = 32'hc404cf5;
      12018: inst = 32'h8220000;
      12019: inst = 32'h10408000;
      12020: inst = 32'hc404cf6;
      12021: inst = 32'h8220000;
      12022: inst = 32'h10408000;
      12023: inst = 32'hc404cf7;
      12024: inst = 32'h8220000;
      12025: inst = 32'h10408000;
      12026: inst = 32'hc404cf8;
      12027: inst = 32'h8220000;
      12028: inst = 32'h10408000;
      12029: inst = 32'hc404cf9;
      12030: inst = 32'h8220000;
      12031: inst = 32'h10408000;
      12032: inst = 32'hc404cfa;
      12033: inst = 32'h8220000;
      12034: inst = 32'h10408000;
      12035: inst = 32'hc404cfe;
      12036: inst = 32'h8220000;
      12037: inst = 32'h10408000;
      12038: inst = 32'hc404d50;
      12039: inst = 32'h8220000;
      12040: inst = 32'h10408000;
      12041: inst = 32'hc404d51;
      12042: inst = 32'h8220000;
      12043: inst = 32'h10408000;
      12044: inst = 32'hc404d52;
      12045: inst = 32'h8220000;
      12046: inst = 32'h10408000;
      12047: inst = 32'hc404d53;
      12048: inst = 32'h8220000;
      12049: inst = 32'h10408000;
      12050: inst = 32'hc404d54;
      12051: inst = 32'h8220000;
      12052: inst = 32'h10408000;
      12053: inst = 32'hc404d55;
      12054: inst = 32'h8220000;
      12055: inst = 32'h10408000;
      12056: inst = 32'hc404d56;
      12057: inst = 32'h8220000;
      12058: inst = 32'h10408000;
      12059: inst = 32'hc404d57;
      12060: inst = 32'h8220000;
      12061: inst = 32'h10408000;
      12062: inst = 32'hc404d58;
      12063: inst = 32'h8220000;
      12064: inst = 32'h10408000;
      12065: inst = 32'hc404d59;
      12066: inst = 32'h8220000;
      12067: inst = 32'h10408000;
      12068: inst = 32'hc404d5a;
      12069: inst = 32'h8220000;
      12070: inst = 32'h10408000;
      12071: inst = 32'hc404d5c;
      12072: inst = 32'h8220000;
      12073: inst = 32'h10408000;
      12074: inst = 32'hc404d5d;
      12075: inst = 32'h8220000;
      12076: inst = 32'h10408000;
      12077: inst = 32'hc404d5e;
      12078: inst = 32'h8220000;
      12079: inst = 32'h10408000;
      12080: inst = 32'hc404db0;
      12081: inst = 32'h8220000;
      12082: inst = 32'h10408000;
      12083: inst = 32'hc404db1;
      12084: inst = 32'h8220000;
      12085: inst = 32'h10408000;
      12086: inst = 32'hc404db2;
      12087: inst = 32'h8220000;
      12088: inst = 32'h10408000;
      12089: inst = 32'hc404db3;
      12090: inst = 32'h8220000;
      12091: inst = 32'h10408000;
      12092: inst = 32'hc404db4;
      12093: inst = 32'h8220000;
      12094: inst = 32'h10408000;
      12095: inst = 32'hc404db5;
      12096: inst = 32'h8220000;
      12097: inst = 32'h10408000;
      12098: inst = 32'hc404db6;
      12099: inst = 32'h8220000;
      12100: inst = 32'h10408000;
      12101: inst = 32'hc404db7;
      12102: inst = 32'h8220000;
      12103: inst = 32'h10408000;
      12104: inst = 32'hc404db8;
      12105: inst = 32'h8220000;
      12106: inst = 32'h10408000;
      12107: inst = 32'hc404db9;
      12108: inst = 32'h8220000;
      12109: inst = 32'h10408000;
      12110: inst = 32'hc404dba;
      12111: inst = 32'h8220000;
      12112: inst = 32'h10408000;
      12113: inst = 32'hc404dbb;
      12114: inst = 32'h8220000;
      12115: inst = 32'h10408000;
      12116: inst = 32'hc404dbc;
      12117: inst = 32'h8220000;
      12118: inst = 32'h10408000;
      12119: inst = 32'hc404dbd;
      12120: inst = 32'h8220000;
      12121: inst = 32'h10408000;
      12122: inst = 32'hc404dbe;
      12123: inst = 32'h8220000;
      12124: inst = 32'h10408000;
      12125: inst = 32'hc404e10;
      12126: inst = 32'h8220000;
      12127: inst = 32'h10408000;
      12128: inst = 32'hc404e11;
      12129: inst = 32'h8220000;
      12130: inst = 32'h10408000;
      12131: inst = 32'hc404e12;
      12132: inst = 32'h8220000;
      12133: inst = 32'h10408000;
      12134: inst = 32'hc404e13;
      12135: inst = 32'h8220000;
      12136: inst = 32'h10408000;
      12137: inst = 32'hc404e14;
      12138: inst = 32'h8220000;
      12139: inst = 32'h10408000;
      12140: inst = 32'hc404e15;
      12141: inst = 32'h8220000;
      12142: inst = 32'h10408000;
      12143: inst = 32'hc404e16;
      12144: inst = 32'h8220000;
      12145: inst = 32'h10408000;
      12146: inst = 32'hc404e17;
      12147: inst = 32'h8220000;
      12148: inst = 32'h10408000;
      12149: inst = 32'hc404e18;
      12150: inst = 32'h8220000;
      12151: inst = 32'h10408000;
      12152: inst = 32'hc404e19;
      12153: inst = 32'h8220000;
      12154: inst = 32'h10408000;
      12155: inst = 32'hc404e1a;
      12156: inst = 32'h8220000;
      12157: inst = 32'h10408000;
      12158: inst = 32'hc404e1b;
      12159: inst = 32'h8220000;
      12160: inst = 32'h10408000;
      12161: inst = 32'hc404e1c;
      12162: inst = 32'h8220000;
      12163: inst = 32'h10408000;
      12164: inst = 32'hc404e1d;
      12165: inst = 32'h8220000;
      12166: inst = 32'h10408000;
      12167: inst = 32'hc404e1e;
      12168: inst = 32'h8220000;
      12169: inst = 32'h10408000;
      12170: inst = 32'hc404e70;
      12171: inst = 32'h8220000;
      12172: inst = 32'h10408000;
      12173: inst = 32'hc404e71;
      12174: inst = 32'h8220000;
      12175: inst = 32'h10408000;
      12176: inst = 32'hc404e72;
      12177: inst = 32'h8220000;
      12178: inst = 32'h10408000;
      12179: inst = 32'hc404e73;
      12180: inst = 32'h8220000;
      12181: inst = 32'h10408000;
      12182: inst = 32'hc404e74;
      12183: inst = 32'h8220000;
      12184: inst = 32'h10408000;
      12185: inst = 32'hc404e75;
      12186: inst = 32'h8220000;
      12187: inst = 32'h10408000;
      12188: inst = 32'hc404e76;
      12189: inst = 32'h8220000;
      12190: inst = 32'h10408000;
      12191: inst = 32'hc404e77;
      12192: inst = 32'h8220000;
      12193: inst = 32'h10408000;
      12194: inst = 32'hc404e78;
      12195: inst = 32'h8220000;
      12196: inst = 32'h10408000;
      12197: inst = 32'hc404e79;
      12198: inst = 32'h8220000;
      12199: inst = 32'h10408000;
      12200: inst = 32'hc404e7a;
      12201: inst = 32'h8220000;
      12202: inst = 32'h10408000;
      12203: inst = 32'hc404e7b;
      12204: inst = 32'h8220000;
      12205: inst = 32'h10408000;
      12206: inst = 32'hc404e7c;
      12207: inst = 32'h8220000;
      12208: inst = 32'h10408000;
      12209: inst = 32'hc404e7d;
      12210: inst = 32'h8220000;
      12211: inst = 32'h10408000;
      12212: inst = 32'hc404e7e;
      12213: inst = 32'h8220000;
      12214: inst = 32'h10408000;
      12215: inst = 32'hc404ed0;
      12216: inst = 32'h8220000;
      12217: inst = 32'h10408000;
      12218: inst = 32'hc404ed1;
      12219: inst = 32'h8220000;
      12220: inst = 32'h10408000;
      12221: inst = 32'hc404ed2;
      12222: inst = 32'h8220000;
      12223: inst = 32'h10408000;
      12224: inst = 32'hc404ed3;
      12225: inst = 32'h8220000;
      12226: inst = 32'h10408000;
      12227: inst = 32'hc404ed4;
      12228: inst = 32'h8220000;
      12229: inst = 32'h10408000;
      12230: inst = 32'hc404ed5;
      12231: inst = 32'h8220000;
      12232: inst = 32'h10408000;
      12233: inst = 32'hc404ed6;
      12234: inst = 32'h8220000;
      12235: inst = 32'h10408000;
      12236: inst = 32'hc404ed7;
      12237: inst = 32'h8220000;
      12238: inst = 32'h10408000;
      12239: inst = 32'hc404ed8;
      12240: inst = 32'h8220000;
      12241: inst = 32'h10408000;
      12242: inst = 32'hc404ed9;
      12243: inst = 32'h8220000;
      12244: inst = 32'h10408000;
      12245: inst = 32'hc404eda;
      12246: inst = 32'h8220000;
      12247: inst = 32'h10408000;
      12248: inst = 32'hc404edb;
      12249: inst = 32'h8220000;
      12250: inst = 32'h10408000;
      12251: inst = 32'hc404edc;
      12252: inst = 32'h8220000;
      12253: inst = 32'h10408000;
      12254: inst = 32'hc404edd;
      12255: inst = 32'h8220000;
      12256: inst = 32'h10408000;
      12257: inst = 32'hc404ede;
      12258: inst = 32'h8220000;
      12259: inst = 32'h10408000;
      12260: inst = 32'hc404f30;
      12261: inst = 32'h8220000;
      12262: inst = 32'h10408000;
      12263: inst = 32'hc404f31;
      12264: inst = 32'h8220000;
      12265: inst = 32'h10408000;
      12266: inst = 32'hc404f32;
      12267: inst = 32'h8220000;
      12268: inst = 32'h10408000;
      12269: inst = 32'hc404f33;
      12270: inst = 32'h8220000;
      12271: inst = 32'h10408000;
      12272: inst = 32'hc404f34;
      12273: inst = 32'h8220000;
      12274: inst = 32'h10408000;
      12275: inst = 32'hc404f35;
      12276: inst = 32'h8220000;
      12277: inst = 32'h10408000;
      12278: inst = 32'hc404f36;
      12279: inst = 32'h8220000;
      12280: inst = 32'h10408000;
      12281: inst = 32'hc404f37;
      12282: inst = 32'h8220000;
      12283: inst = 32'h10408000;
      12284: inst = 32'hc404f38;
      12285: inst = 32'h8220000;
      12286: inst = 32'h10408000;
      12287: inst = 32'hc404f39;
      12288: inst = 32'h8220000;
      12289: inst = 32'h10408000;
      12290: inst = 32'hc404f3a;
      12291: inst = 32'h8220000;
      12292: inst = 32'h10408000;
      12293: inst = 32'hc404f3b;
      12294: inst = 32'h8220000;
      12295: inst = 32'h10408000;
      12296: inst = 32'hc404f3c;
      12297: inst = 32'h8220000;
      12298: inst = 32'h10408000;
      12299: inst = 32'hc404f3d;
      12300: inst = 32'h8220000;
      12301: inst = 32'h10408000;
      12302: inst = 32'hc404f3e;
      12303: inst = 32'h8220000;
      12304: inst = 32'h10408000;
      12305: inst = 32'hc404f90;
      12306: inst = 32'h8220000;
      12307: inst = 32'h10408000;
      12308: inst = 32'hc404f91;
      12309: inst = 32'h8220000;
      12310: inst = 32'h10408000;
      12311: inst = 32'hc404f92;
      12312: inst = 32'h8220000;
      12313: inst = 32'h10408000;
      12314: inst = 32'hc404f93;
      12315: inst = 32'h8220000;
      12316: inst = 32'h10408000;
      12317: inst = 32'hc404f94;
      12318: inst = 32'h8220000;
      12319: inst = 32'h10408000;
      12320: inst = 32'hc404f95;
      12321: inst = 32'h8220000;
      12322: inst = 32'h10408000;
      12323: inst = 32'hc404f96;
      12324: inst = 32'h8220000;
      12325: inst = 32'h10408000;
      12326: inst = 32'hc404f97;
      12327: inst = 32'h8220000;
      12328: inst = 32'h10408000;
      12329: inst = 32'hc404f98;
      12330: inst = 32'h8220000;
      12331: inst = 32'h10408000;
      12332: inst = 32'hc404f99;
      12333: inst = 32'h8220000;
      12334: inst = 32'h10408000;
      12335: inst = 32'hc404f9a;
      12336: inst = 32'h8220000;
      12337: inst = 32'h10408000;
      12338: inst = 32'hc404f9b;
      12339: inst = 32'h8220000;
      12340: inst = 32'h10408000;
      12341: inst = 32'hc404f9c;
      12342: inst = 32'h8220000;
      12343: inst = 32'h10408000;
      12344: inst = 32'hc404f9d;
      12345: inst = 32'h8220000;
      12346: inst = 32'h10408000;
      12347: inst = 32'hc404f9e;
      12348: inst = 32'h8220000;
      12349: inst = 32'h10408000;
      12350: inst = 32'hc404ff0;
      12351: inst = 32'h8220000;
      12352: inst = 32'h10408000;
      12353: inst = 32'hc404ff1;
      12354: inst = 32'h8220000;
      12355: inst = 32'h10408000;
      12356: inst = 32'hc404ff2;
      12357: inst = 32'h8220000;
      12358: inst = 32'h10408000;
      12359: inst = 32'hc404ff3;
      12360: inst = 32'h8220000;
      12361: inst = 32'h10408000;
      12362: inst = 32'hc404ff4;
      12363: inst = 32'h8220000;
      12364: inst = 32'h10408000;
      12365: inst = 32'hc404ff5;
      12366: inst = 32'h8220000;
      12367: inst = 32'h10408000;
      12368: inst = 32'hc404ff6;
      12369: inst = 32'h8220000;
      12370: inst = 32'h10408000;
      12371: inst = 32'hc404ff7;
      12372: inst = 32'h8220000;
      12373: inst = 32'h10408000;
      12374: inst = 32'hc404ff8;
      12375: inst = 32'h8220000;
      12376: inst = 32'h10408000;
      12377: inst = 32'hc404ff9;
      12378: inst = 32'h8220000;
      12379: inst = 32'h10408000;
      12380: inst = 32'hc404ffa;
      12381: inst = 32'h8220000;
      12382: inst = 32'h10408000;
      12383: inst = 32'hc404ffb;
      12384: inst = 32'h8220000;
      12385: inst = 32'h10408000;
      12386: inst = 32'hc404ffc;
      12387: inst = 32'h8220000;
      12388: inst = 32'h10408000;
      12389: inst = 32'hc404ffd;
      12390: inst = 32'h8220000;
      12391: inst = 32'h10408000;
      12392: inst = 32'hc404ffe;
      12393: inst = 32'h8220000;
      12394: inst = 32'h10408000;
      12395: inst = 32'hc405050;
      12396: inst = 32'h8220000;
      12397: inst = 32'h10408000;
      12398: inst = 32'hc405051;
      12399: inst = 32'h8220000;
      12400: inst = 32'h10408000;
      12401: inst = 32'hc405052;
      12402: inst = 32'h8220000;
      12403: inst = 32'h10408000;
      12404: inst = 32'hc405053;
      12405: inst = 32'h8220000;
      12406: inst = 32'h10408000;
      12407: inst = 32'hc405054;
      12408: inst = 32'h8220000;
      12409: inst = 32'h10408000;
      12410: inst = 32'hc405055;
      12411: inst = 32'h8220000;
      12412: inst = 32'h10408000;
      12413: inst = 32'hc405056;
      12414: inst = 32'h8220000;
      12415: inst = 32'h10408000;
      12416: inst = 32'hc405057;
      12417: inst = 32'h8220000;
      12418: inst = 32'h10408000;
      12419: inst = 32'hc405058;
      12420: inst = 32'h8220000;
      12421: inst = 32'h10408000;
      12422: inst = 32'hc405059;
      12423: inst = 32'h8220000;
      12424: inst = 32'h10408000;
      12425: inst = 32'hc40505a;
      12426: inst = 32'h8220000;
      12427: inst = 32'h10408000;
      12428: inst = 32'hc40505b;
      12429: inst = 32'h8220000;
      12430: inst = 32'h10408000;
      12431: inst = 32'hc40505c;
      12432: inst = 32'h8220000;
      12433: inst = 32'h10408000;
      12434: inst = 32'hc40505d;
      12435: inst = 32'h8220000;
      12436: inst = 32'h10408000;
      12437: inst = 32'hc40505e;
      12438: inst = 32'h8220000;
      12439: inst = 32'h10408000;
      12440: inst = 32'hc4050b0;
      12441: inst = 32'h8220000;
      12442: inst = 32'h10408000;
      12443: inst = 32'hc4050b1;
      12444: inst = 32'h8220000;
      12445: inst = 32'h10408000;
      12446: inst = 32'hc4050b2;
      12447: inst = 32'h8220000;
      12448: inst = 32'h10408000;
      12449: inst = 32'hc4050b3;
      12450: inst = 32'h8220000;
      12451: inst = 32'h10408000;
      12452: inst = 32'hc4050b4;
      12453: inst = 32'h8220000;
      12454: inst = 32'h10408000;
      12455: inst = 32'hc4050b5;
      12456: inst = 32'h8220000;
      12457: inst = 32'h10408000;
      12458: inst = 32'hc4050b6;
      12459: inst = 32'h8220000;
      12460: inst = 32'h10408000;
      12461: inst = 32'hc4050b7;
      12462: inst = 32'h8220000;
      12463: inst = 32'h10408000;
      12464: inst = 32'hc4050b8;
      12465: inst = 32'h8220000;
      12466: inst = 32'h10408000;
      12467: inst = 32'hc4050b9;
      12468: inst = 32'h8220000;
      12469: inst = 32'h10408000;
      12470: inst = 32'hc4050ba;
      12471: inst = 32'h8220000;
      12472: inst = 32'h10408000;
      12473: inst = 32'hc4050bb;
      12474: inst = 32'h8220000;
      12475: inst = 32'h10408000;
      12476: inst = 32'hc4050bc;
      12477: inst = 32'h8220000;
      12478: inst = 32'h10408000;
      12479: inst = 32'hc4050bd;
      12480: inst = 32'h8220000;
      12481: inst = 32'h10408000;
      12482: inst = 32'hc4050be;
      12483: inst = 32'h8220000;
      12484: inst = 32'h10408000;
      12485: inst = 32'hc405110;
      12486: inst = 32'h8220000;
      12487: inst = 32'h10408000;
      12488: inst = 32'hc405111;
      12489: inst = 32'h8220000;
      12490: inst = 32'h10408000;
      12491: inst = 32'hc405112;
      12492: inst = 32'h8220000;
      12493: inst = 32'h10408000;
      12494: inst = 32'hc405113;
      12495: inst = 32'h8220000;
      12496: inst = 32'h10408000;
      12497: inst = 32'hc405114;
      12498: inst = 32'h8220000;
      12499: inst = 32'h10408000;
      12500: inst = 32'hc405115;
      12501: inst = 32'h8220000;
      12502: inst = 32'h10408000;
      12503: inst = 32'hc405116;
      12504: inst = 32'h8220000;
      12505: inst = 32'h10408000;
      12506: inst = 32'hc405117;
      12507: inst = 32'h8220000;
      12508: inst = 32'h10408000;
      12509: inst = 32'hc405118;
      12510: inst = 32'h8220000;
      12511: inst = 32'h10408000;
      12512: inst = 32'hc405119;
      12513: inst = 32'h8220000;
      12514: inst = 32'h10408000;
      12515: inst = 32'hc40511a;
      12516: inst = 32'h8220000;
      12517: inst = 32'h10408000;
      12518: inst = 32'hc40511b;
      12519: inst = 32'h8220000;
      12520: inst = 32'h10408000;
      12521: inst = 32'hc40511c;
      12522: inst = 32'h8220000;
      12523: inst = 32'h10408000;
      12524: inst = 32'hc40511d;
      12525: inst = 32'h8220000;
      12526: inst = 32'h10408000;
      12527: inst = 32'hc40511e;
      12528: inst = 32'h8220000;
      12529: inst = 32'h10408000;
      12530: inst = 32'hc405170;
      12531: inst = 32'h8220000;
      12532: inst = 32'h10408000;
      12533: inst = 32'hc405171;
      12534: inst = 32'h8220000;
      12535: inst = 32'h10408000;
      12536: inst = 32'hc405172;
      12537: inst = 32'h8220000;
      12538: inst = 32'h10408000;
      12539: inst = 32'hc405173;
      12540: inst = 32'h8220000;
      12541: inst = 32'h10408000;
      12542: inst = 32'hc405174;
      12543: inst = 32'h8220000;
      12544: inst = 32'h10408000;
      12545: inst = 32'hc405175;
      12546: inst = 32'h8220000;
      12547: inst = 32'h10408000;
      12548: inst = 32'hc405176;
      12549: inst = 32'h8220000;
      12550: inst = 32'h10408000;
      12551: inst = 32'hc405177;
      12552: inst = 32'h8220000;
      12553: inst = 32'h10408000;
      12554: inst = 32'hc405178;
      12555: inst = 32'h8220000;
      12556: inst = 32'h10408000;
      12557: inst = 32'hc405179;
      12558: inst = 32'h8220000;
      12559: inst = 32'h10408000;
      12560: inst = 32'hc40517a;
      12561: inst = 32'h8220000;
      12562: inst = 32'h10408000;
      12563: inst = 32'hc40517b;
      12564: inst = 32'h8220000;
      12565: inst = 32'h10408000;
      12566: inst = 32'hc40517c;
      12567: inst = 32'h8220000;
      12568: inst = 32'h10408000;
      12569: inst = 32'hc40517d;
      12570: inst = 32'h8220000;
      12571: inst = 32'h10408000;
      12572: inst = 32'hc40517e;
      12573: inst = 32'h8220000;
      12574: inst = 32'h10408000;
      12575: inst = 32'hc4051d0;
      12576: inst = 32'h8220000;
      12577: inst = 32'h10408000;
      12578: inst = 32'hc4051d1;
      12579: inst = 32'h8220000;
      12580: inst = 32'h10408000;
      12581: inst = 32'hc4051d2;
      12582: inst = 32'h8220000;
      12583: inst = 32'h10408000;
      12584: inst = 32'hc4051d3;
      12585: inst = 32'h8220000;
      12586: inst = 32'h10408000;
      12587: inst = 32'hc4051d4;
      12588: inst = 32'h8220000;
      12589: inst = 32'h10408000;
      12590: inst = 32'hc4051d5;
      12591: inst = 32'h8220000;
      12592: inst = 32'h10408000;
      12593: inst = 32'hc4051d6;
      12594: inst = 32'h8220000;
      12595: inst = 32'h10408000;
      12596: inst = 32'hc4051d7;
      12597: inst = 32'h8220000;
      12598: inst = 32'h10408000;
      12599: inst = 32'hc4051d8;
      12600: inst = 32'h8220000;
      12601: inst = 32'h10408000;
      12602: inst = 32'hc4051d9;
      12603: inst = 32'h8220000;
      12604: inst = 32'h10408000;
      12605: inst = 32'hc4051da;
      12606: inst = 32'h8220000;
      12607: inst = 32'h10408000;
      12608: inst = 32'hc4051db;
      12609: inst = 32'h8220000;
      12610: inst = 32'h10408000;
      12611: inst = 32'hc4051dc;
      12612: inst = 32'h8220000;
      12613: inst = 32'h10408000;
      12614: inst = 32'hc4051dd;
      12615: inst = 32'h8220000;
      12616: inst = 32'h10408000;
      12617: inst = 32'hc4051de;
      12618: inst = 32'h8220000;
      12619: inst = 32'h10408000;
      12620: inst = 32'hc405230;
      12621: inst = 32'h8220000;
      12622: inst = 32'h10408000;
      12623: inst = 32'hc405231;
      12624: inst = 32'h8220000;
      12625: inst = 32'h10408000;
      12626: inst = 32'hc405232;
      12627: inst = 32'h8220000;
      12628: inst = 32'h10408000;
      12629: inst = 32'hc405233;
      12630: inst = 32'h8220000;
      12631: inst = 32'h10408000;
      12632: inst = 32'hc405234;
      12633: inst = 32'h8220000;
      12634: inst = 32'h10408000;
      12635: inst = 32'hc405235;
      12636: inst = 32'h8220000;
      12637: inst = 32'h10408000;
      12638: inst = 32'hc405236;
      12639: inst = 32'h8220000;
      12640: inst = 32'h10408000;
      12641: inst = 32'hc405237;
      12642: inst = 32'h8220000;
      12643: inst = 32'h10408000;
      12644: inst = 32'hc405238;
      12645: inst = 32'h8220000;
      12646: inst = 32'h10408000;
      12647: inst = 32'hc405239;
      12648: inst = 32'h8220000;
      12649: inst = 32'h10408000;
      12650: inst = 32'hc40523a;
      12651: inst = 32'h8220000;
      12652: inst = 32'h10408000;
      12653: inst = 32'hc40523b;
      12654: inst = 32'h8220000;
      12655: inst = 32'h10408000;
      12656: inst = 32'hc40523c;
      12657: inst = 32'h8220000;
      12658: inst = 32'h10408000;
      12659: inst = 32'hc40523d;
      12660: inst = 32'h8220000;
      12661: inst = 32'h10408000;
      12662: inst = 32'hc40523e;
      12663: inst = 32'h8220000;
      12664: inst = 32'h10408000;
      12665: inst = 32'hc405290;
      12666: inst = 32'h8220000;
      12667: inst = 32'h10408000;
      12668: inst = 32'hc405291;
      12669: inst = 32'h8220000;
      12670: inst = 32'h10408000;
      12671: inst = 32'hc405292;
      12672: inst = 32'h8220000;
      12673: inst = 32'h10408000;
      12674: inst = 32'hc405293;
      12675: inst = 32'h8220000;
      12676: inst = 32'h10408000;
      12677: inst = 32'hc405294;
      12678: inst = 32'h8220000;
      12679: inst = 32'h10408000;
      12680: inst = 32'hc405295;
      12681: inst = 32'h8220000;
      12682: inst = 32'h10408000;
      12683: inst = 32'hc405296;
      12684: inst = 32'h8220000;
      12685: inst = 32'h10408000;
      12686: inst = 32'hc405297;
      12687: inst = 32'h8220000;
      12688: inst = 32'h10408000;
      12689: inst = 32'hc405298;
      12690: inst = 32'h8220000;
      12691: inst = 32'h10408000;
      12692: inst = 32'hc405299;
      12693: inst = 32'h8220000;
      12694: inst = 32'h10408000;
      12695: inst = 32'hc40529a;
      12696: inst = 32'h8220000;
      12697: inst = 32'h10408000;
      12698: inst = 32'hc40529b;
      12699: inst = 32'h8220000;
      12700: inst = 32'h10408000;
      12701: inst = 32'hc40529c;
      12702: inst = 32'h8220000;
      12703: inst = 32'h10408000;
      12704: inst = 32'hc40529d;
      12705: inst = 32'h8220000;
      12706: inst = 32'h10408000;
      12707: inst = 32'hc40529e;
      12708: inst = 32'h8220000;
      12709: inst = 32'hc20ef7c;
      12710: inst = 32'h10408000;
      12711: inst = 32'hc404932;
      12712: inst = 32'h8220000;
      12713: inst = 32'h10408000;
      12714: inst = 32'hc404933;
      12715: inst = 32'h8220000;
      12716: inst = 32'h10408000;
      12717: inst = 32'hc404934;
      12718: inst = 32'h8220000;
      12719: inst = 32'h10408000;
      12720: inst = 32'hc404935;
      12721: inst = 32'h8220000;
      12722: inst = 32'h10408000;
      12723: inst = 32'hc404993;
      12724: inst = 32'h8220000;
      12725: inst = 32'h10408000;
      12726: inst = 32'hc404994;
      12727: inst = 32'h8220000;
      12728: inst = 32'h10408000;
      12729: inst = 32'hc404995;
      12730: inst = 32'h8220000;
      12731: inst = 32'h10408000;
      12732: inst = 32'hc4049f3;
      12733: inst = 32'h8220000;
      12734: inst = 32'h10408000;
      12735: inst = 32'hc4049f4;
      12736: inst = 32'h8220000;
      12737: inst = 32'h10408000;
      12738: inst = 32'hc4049f5;
      12739: inst = 32'h8220000;
      12740: inst = 32'h10408000;
      12741: inst = 32'hc404a53;
      12742: inst = 32'h8220000;
      12743: inst = 32'h10408000;
      12744: inst = 32'hc404a54;
      12745: inst = 32'h8220000;
      12746: inst = 32'h10408000;
      12747: inst = 32'hc404a55;
      12748: inst = 32'h8220000;
      12749: inst = 32'h10408000;
      12750: inst = 32'hc404ab2;
      12751: inst = 32'h8220000;
      12752: inst = 32'h10408000;
      12753: inst = 32'hc404ab3;
      12754: inst = 32'h8220000;
      12755: inst = 32'h10408000;
      12756: inst = 32'hc404ab5;
      12757: inst = 32'h8220000;
      12758: inst = 32'h10408000;
      12759: inst = 32'hc404b12;
      12760: inst = 32'h8220000;
      12761: inst = 32'h10408000;
      12762: inst = 32'hc404b13;
      12763: inst = 32'h8220000;
      12764: inst = 32'h10408000;
      12765: inst = 32'hc404b15;
      12766: inst = 32'h8220000;
      12767: inst = 32'h10408000;
      12768: inst = 32'hc404b72;
      12769: inst = 32'h8220000;
      12770: inst = 32'h10408000;
      12771: inst = 32'hc404b73;
      12772: inst = 32'h8220000;
      12773: inst = 32'h10408000;
      12774: inst = 32'hc404b74;
      12775: inst = 32'h8220000;
      12776: inst = 32'h10408000;
      12777: inst = 32'hc404b75;
      12778: inst = 32'h8220000;
      12779: inst = 32'hc20eed7;
      12780: inst = 32'h10408000;
      12781: inst = 32'hc404a08;
      12782: inst = 32'h8220000;
      12783: inst = 32'h10408000;
      12784: inst = 32'hc404a0e;
      12785: inst = 32'h8220000;
      12786: inst = 32'hc20e6fa;
      12787: inst = 32'h10408000;
      12788: inst = 32'hc404a09;
      12789: inst = 32'h8220000;
      12790: inst = 32'h10408000;
      12791: inst = 32'hc404a0d;
      12792: inst = 32'h8220000;
      12793: inst = 32'h10408000;
      12794: inst = 32'hc404be7;
      12795: inst = 32'h8220000;
      12796: inst = 32'hc20e6fb;
      12797: inst = 32'h10408000;
      12798: inst = 32'hc404a0a;
      12799: inst = 32'h8220000;
      12800: inst = 32'h10408000;
      12801: inst = 32'hc404a0c;
      12802: inst = 32'h8220000;
      12803: inst = 32'h10408000;
      12804: inst = 32'hc404ac7;
      12805: inst = 32'h8220000;
      12806: inst = 32'h10408000;
      12807: inst = 32'hc404acf;
      12808: inst = 32'h8220000;
      12809: inst = 32'h10408000;
      12810: inst = 32'hc404b87;
      12811: inst = 32'h8220000;
      12812: inst = 32'h10408000;
      12813: inst = 32'hc404b8f;
      12814: inst = 32'h8220000;
      12815: inst = 32'h10408000;
      12816: inst = 32'hc404c4d;
      12817: inst = 32'h8220000;
      12818: inst = 32'hc20defb;
      12819: inst = 32'h10408000;
      12820: inst = 32'hc404a0b;
      12821: inst = 32'h8220000;
      12822: inst = 32'h10408000;
      12823: inst = 32'hc404a68;
      12824: inst = 32'h8220000;
      12825: inst = 32'h10408000;
      12826: inst = 32'hc404a69;
      12827: inst = 32'h8220000;
      12828: inst = 32'h10408000;
      12829: inst = 32'hc404a6a;
      12830: inst = 32'h8220000;
      12831: inst = 32'h10408000;
      12832: inst = 32'hc404a6b;
      12833: inst = 32'h8220000;
      12834: inst = 32'h10408000;
      12835: inst = 32'hc404a6c;
      12836: inst = 32'h8220000;
      12837: inst = 32'h10408000;
      12838: inst = 32'hc404a6d;
      12839: inst = 32'h8220000;
      12840: inst = 32'h10408000;
      12841: inst = 32'hc404a6e;
      12842: inst = 32'h8220000;
      12843: inst = 32'h10408000;
      12844: inst = 32'hc404ac8;
      12845: inst = 32'h8220000;
      12846: inst = 32'h10408000;
      12847: inst = 32'hc404ac9;
      12848: inst = 32'h8220000;
      12849: inst = 32'h10408000;
      12850: inst = 32'hc404aca;
      12851: inst = 32'h8220000;
      12852: inst = 32'h10408000;
      12853: inst = 32'hc404acb;
      12854: inst = 32'h8220000;
      12855: inst = 32'h10408000;
      12856: inst = 32'hc404acc;
      12857: inst = 32'h8220000;
      12858: inst = 32'h10408000;
      12859: inst = 32'hc404acd;
      12860: inst = 32'h8220000;
      12861: inst = 32'h10408000;
      12862: inst = 32'hc404ace;
      12863: inst = 32'h8220000;
      12864: inst = 32'h10408000;
      12865: inst = 32'hc404b27;
      12866: inst = 32'h8220000;
      12867: inst = 32'h10408000;
      12868: inst = 32'hc404b2a;
      12869: inst = 32'h8220000;
      12870: inst = 32'h10408000;
      12871: inst = 32'hc404b2d;
      12872: inst = 32'h8220000;
      12873: inst = 32'h10408000;
      12874: inst = 32'hc404b2e;
      12875: inst = 32'h8220000;
      12876: inst = 32'h10408000;
      12877: inst = 32'hc404b2f;
      12878: inst = 32'h8220000;
      12879: inst = 32'h10408000;
      12880: inst = 32'hc404b8a;
      12881: inst = 32'h8220000;
      12882: inst = 32'h10408000;
      12883: inst = 32'hc404b8d;
      12884: inst = 32'h8220000;
      12885: inst = 32'h10408000;
      12886: inst = 32'hc404b8e;
      12887: inst = 32'h8220000;
      12888: inst = 32'h10408000;
      12889: inst = 32'hc404be8;
      12890: inst = 32'h8220000;
      12891: inst = 32'h10408000;
      12892: inst = 32'hc404be9;
      12893: inst = 32'h8220000;
      12894: inst = 32'h10408000;
      12895: inst = 32'hc404bea;
      12896: inst = 32'h8220000;
      12897: inst = 32'h10408000;
      12898: inst = 32'hc404beb;
      12899: inst = 32'h8220000;
      12900: inst = 32'h10408000;
      12901: inst = 32'hc404bec;
      12902: inst = 32'h8220000;
      12903: inst = 32'h10408000;
      12904: inst = 32'hc404bed;
      12905: inst = 32'h8220000;
      12906: inst = 32'h10408000;
      12907: inst = 32'hc404bee;
      12908: inst = 32'h8220000;
      12909: inst = 32'h10408000;
      12910: inst = 32'hc404c49;
      12911: inst = 32'h8220000;
      12912: inst = 32'h10408000;
      12913: inst = 32'hc404c4b;
      12914: inst = 32'h8220000;
      12915: inst = 32'h10408000;
      12916: inst = 32'hc404ca9;
      12917: inst = 32'h8220000;
      12918: inst = 32'h10408000;
      12919: inst = 32'hc404cab;
      12920: inst = 32'h8220000;
      12921: inst = 32'hc20eed8;
      12922: inst = 32'h10408000;
      12923: inst = 32'hc404a67;
      12924: inst = 32'h8220000;
      12925: inst = 32'h10408000;
      12926: inst = 32'hc404a6f;
      12927: inst = 32'h8220000;
      12928: inst = 32'hc204a69;
      12929: inst = 32'h10408000;
      12930: inst = 32'hc404b28;
      12931: inst = 32'h8220000;
      12932: inst = 32'h10408000;
      12933: inst = 32'hc404b29;
      12934: inst = 32'h8220000;
      12935: inst = 32'h10408000;
      12936: inst = 32'hc404b2b;
      12937: inst = 32'h8220000;
      12938: inst = 32'h10408000;
      12939: inst = 32'hc404b2c;
      12940: inst = 32'h8220000;
      12941: inst = 32'h10408000;
      12942: inst = 32'hc404b88;
      12943: inst = 32'h8220000;
      12944: inst = 32'h10408000;
      12945: inst = 32'hc404b89;
      12946: inst = 32'h8220000;
      12947: inst = 32'h10408000;
      12948: inst = 32'hc404b8b;
      12949: inst = 32'h8220000;
      12950: inst = 32'h10408000;
      12951: inst = 32'hc404b8c;
      12952: inst = 32'h8220000;
      12953: inst = 32'h10408000;
      12954: inst = 32'hc404c48;
      12955: inst = 32'h8220000;
      12956: inst = 32'h10408000;
      12957: inst = 32'hc404c4a;
      12958: inst = 32'h8220000;
      12959: inst = 32'h10408000;
      12960: inst = 32'hc404c4c;
      12961: inst = 32'h8220000;
      12962: inst = 32'h10408000;
      12963: inst = 32'hc404ca8;
      12964: inst = 32'h8220000;
      12965: inst = 32'h10408000;
      12966: inst = 32'hc404caa;
      12967: inst = 32'h8220000;
      12968: inst = 32'h10408000;
      12969: inst = 32'hc404cac;
      12970: inst = 32'h8220000;
      12971: inst = 32'h10408000;
      12972: inst = 32'hc405085;
      12973: inst = 32'h8220000;
      12974: inst = 32'h10408000;
      12975: inst = 32'hc40509a;
      12976: inst = 32'h8220000;
      12977: inst = 32'h10408000;
      12978: inst = 32'hc4050e4;
      12979: inst = 32'h8220000;
      12980: inst = 32'h10408000;
      12981: inst = 32'hc4050e5;
      12982: inst = 32'h8220000;
      12983: inst = 32'h10408000;
      12984: inst = 32'hc4050fa;
      12985: inst = 32'h8220000;
      12986: inst = 32'h10408000;
      12987: inst = 32'hc4050fb;
      12988: inst = 32'h8220000;
      12989: inst = 32'h10408000;
      12990: inst = 32'hc405143;
      12991: inst = 32'h8220000;
      12992: inst = 32'h10408000;
      12993: inst = 32'hc405144;
      12994: inst = 32'h8220000;
      12995: inst = 32'h10408000;
      12996: inst = 32'hc405145;
      12997: inst = 32'h8220000;
      12998: inst = 32'h10408000;
      12999: inst = 32'hc40515a;
      13000: inst = 32'h8220000;
      13001: inst = 32'h10408000;
      13002: inst = 32'hc40515b;
      13003: inst = 32'h8220000;
      13004: inst = 32'h10408000;
      13005: inst = 32'hc40515c;
      13006: inst = 32'h8220000;
      13007: inst = 32'h10408000;
      13008: inst = 32'hc4051a2;
      13009: inst = 32'h8220000;
      13010: inst = 32'h10408000;
      13011: inst = 32'hc4051a3;
      13012: inst = 32'h8220000;
      13013: inst = 32'h10408000;
      13014: inst = 32'hc4051a4;
      13015: inst = 32'h8220000;
      13016: inst = 32'h10408000;
      13017: inst = 32'hc4051a5;
      13018: inst = 32'h8220000;
      13019: inst = 32'h10408000;
      13020: inst = 32'hc4051ba;
      13021: inst = 32'h8220000;
      13022: inst = 32'h10408000;
      13023: inst = 32'hc4051bb;
      13024: inst = 32'h8220000;
      13025: inst = 32'h10408000;
      13026: inst = 32'hc4051bc;
      13027: inst = 32'h8220000;
      13028: inst = 32'h10408000;
      13029: inst = 32'hc4051bd;
      13030: inst = 32'h8220000;
      13031: inst = 32'h10408000;
      13032: inst = 32'hc405202;
      13033: inst = 32'h8220000;
      13034: inst = 32'h10408000;
      13035: inst = 32'hc405203;
      13036: inst = 32'h8220000;
      13037: inst = 32'h10408000;
      13038: inst = 32'hc405204;
      13039: inst = 32'h8220000;
      13040: inst = 32'h10408000;
      13041: inst = 32'hc405205;
      13042: inst = 32'h8220000;
      13043: inst = 32'h10408000;
      13044: inst = 32'hc40521a;
      13045: inst = 32'h8220000;
      13046: inst = 32'h10408000;
      13047: inst = 32'hc40521b;
      13048: inst = 32'h8220000;
      13049: inst = 32'h10408000;
      13050: inst = 32'hc40521c;
      13051: inst = 32'h8220000;
      13052: inst = 32'h10408000;
      13053: inst = 32'hc40521d;
      13054: inst = 32'h8220000;
      13055: inst = 32'h10408000;
      13056: inst = 32'hc405262;
      13057: inst = 32'h8220000;
      13058: inst = 32'h10408000;
      13059: inst = 32'hc405263;
      13060: inst = 32'h8220000;
      13061: inst = 32'h10408000;
      13062: inst = 32'hc405264;
      13063: inst = 32'h8220000;
      13064: inst = 32'h10408000;
      13065: inst = 32'hc405265;
      13066: inst = 32'h8220000;
      13067: inst = 32'h10408000;
      13068: inst = 32'hc40527a;
      13069: inst = 32'h8220000;
      13070: inst = 32'h10408000;
      13071: inst = 32'hc40527b;
      13072: inst = 32'h8220000;
      13073: inst = 32'h10408000;
      13074: inst = 32'hc40527c;
      13075: inst = 32'h8220000;
      13076: inst = 32'h10408000;
      13077: inst = 32'hc40527d;
      13078: inst = 32'h8220000;
      13079: inst = 32'h10408000;
      13080: inst = 32'hc4052c2;
      13081: inst = 32'h8220000;
      13082: inst = 32'h10408000;
      13083: inst = 32'hc4052c3;
      13084: inst = 32'h8220000;
      13085: inst = 32'h10408000;
      13086: inst = 32'hc4052c4;
      13087: inst = 32'h8220000;
      13088: inst = 32'h10408000;
      13089: inst = 32'hc4052db;
      13090: inst = 32'h8220000;
      13091: inst = 32'h10408000;
      13092: inst = 32'hc4052dc;
      13093: inst = 32'h8220000;
      13094: inst = 32'h10408000;
      13095: inst = 32'hc4052dd;
      13096: inst = 32'h8220000;
      13097: inst = 32'h10408000;
      13098: inst = 32'hc405322;
      13099: inst = 32'h8220000;
      13100: inst = 32'h10408000;
      13101: inst = 32'hc405323;
      13102: inst = 32'h8220000;
      13103: inst = 32'h10408000;
      13104: inst = 32'hc405324;
      13105: inst = 32'h8220000;
      13106: inst = 32'h10408000;
      13107: inst = 32'hc40533b;
      13108: inst = 32'h8220000;
      13109: inst = 32'h10408000;
      13110: inst = 32'hc40533c;
      13111: inst = 32'h8220000;
      13112: inst = 32'h10408000;
      13113: inst = 32'hc40533d;
      13114: inst = 32'h8220000;
      13115: inst = 32'h10408000;
      13116: inst = 32'hc40537f;
      13117: inst = 32'h8220000;
      13118: inst = 32'h10408000;
      13119: inst = 32'hc405382;
      13120: inst = 32'h8220000;
      13121: inst = 32'h10408000;
      13122: inst = 32'hc405383;
      13123: inst = 32'h8220000;
      13124: inst = 32'h10408000;
      13125: inst = 32'hc405384;
      13126: inst = 32'h8220000;
      13127: inst = 32'h10408000;
      13128: inst = 32'hc40539b;
      13129: inst = 32'h8220000;
      13130: inst = 32'h10408000;
      13131: inst = 32'hc40539c;
      13132: inst = 32'h8220000;
      13133: inst = 32'h10408000;
      13134: inst = 32'hc40539d;
      13135: inst = 32'h8220000;
      13136: inst = 32'h10408000;
      13137: inst = 32'hc4053a0;
      13138: inst = 32'h8220000;
      13139: inst = 32'h10408000;
      13140: inst = 32'hc4053de;
      13141: inst = 32'h8220000;
      13142: inst = 32'h10408000;
      13143: inst = 32'hc4053df;
      13144: inst = 32'h8220000;
      13145: inst = 32'h10408000;
      13146: inst = 32'hc4053e2;
      13147: inst = 32'h8220000;
      13148: inst = 32'h10408000;
      13149: inst = 32'hc4053e3;
      13150: inst = 32'h8220000;
      13151: inst = 32'h10408000;
      13152: inst = 32'hc4053fc;
      13153: inst = 32'h8220000;
      13154: inst = 32'h10408000;
      13155: inst = 32'hc4053fd;
      13156: inst = 32'h8220000;
      13157: inst = 32'h10408000;
      13158: inst = 32'hc405400;
      13159: inst = 32'h8220000;
      13160: inst = 32'h10408000;
      13161: inst = 32'hc405401;
      13162: inst = 32'h8220000;
      13163: inst = 32'h10408000;
      13164: inst = 32'hc40543d;
      13165: inst = 32'h8220000;
      13166: inst = 32'h10408000;
      13167: inst = 32'hc40543e;
      13168: inst = 32'h8220000;
      13169: inst = 32'h10408000;
      13170: inst = 32'hc40543f;
      13171: inst = 32'h8220000;
      13172: inst = 32'h10408000;
      13173: inst = 32'hc405442;
      13174: inst = 32'h8220000;
      13175: inst = 32'h10408000;
      13176: inst = 32'hc405443;
      13177: inst = 32'h8220000;
      13178: inst = 32'h10408000;
      13179: inst = 32'hc40545c;
      13180: inst = 32'h8220000;
      13181: inst = 32'h10408000;
      13182: inst = 32'hc40545d;
      13183: inst = 32'h8220000;
      13184: inst = 32'h10408000;
      13185: inst = 32'hc405460;
      13186: inst = 32'h8220000;
      13187: inst = 32'h10408000;
      13188: inst = 32'hc405461;
      13189: inst = 32'h8220000;
      13190: inst = 32'h10408000;
      13191: inst = 32'hc405462;
      13192: inst = 32'h8220000;
      13193: inst = 32'h10408000;
      13194: inst = 32'hc40549d;
      13195: inst = 32'h8220000;
      13196: inst = 32'h10408000;
      13197: inst = 32'hc40549e;
      13198: inst = 32'h8220000;
      13199: inst = 32'h10408000;
      13200: inst = 32'hc4054a0;
      13201: inst = 32'h8220000;
      13202: inst = 32'h10408000;
      13203: inst = 32'hc4054a1;
      13204: inst = 32'h8220000;
      13205: inst = 32'h10408000;
      13206: inst = 32'hc4054a2;
      13207: inst = 32'h8220000;
      13208: inst = 32'h10408000;
      13209: inst = 32'hc4054a3;
      13210: inst = 32'h8220000;
      13211: inst = 32'h10408000;
      13212: inst = 32'hc4054bc;
      13213: inst = 32'h8220000;
      13214: inst = 32'h10408000;
      13215: inst = 32'hc4054bd;
      13216: inst = 32'h8220000;
      13217: inst = 32'h10408000;
      13218: inst = 32'hc4054be;
      13219: inst = 32'h8220000;
      13220: inst = 32'h10408000;
      13221: inst = 32'hc4054bf;
      13222: inst = 32'h8220000;
      13223: inst = 32'h10408000;
      13224: inst = 32'hc4054c1;
      13225: inst = 32'h8220000;
      13226: inst = 32'h10408000;
      13227: inst = 32'hc4054c2;
      13228: inst = 32'h8220000;
      13229: inst = 32'h10408000;
      13230: inst = 32'hc4054fc;
      13231: inst = 32'h8220000;
      13232: inst = 32'h10408000;
      13233: inst = 32'hc4054fd;
      13234: inst = 32'h8220000;
      13235: inst = 32'h10408000;
      13236: inst = 32'hc4054fe;
      13237: inst = 32'h8220000;
      13238: inst = 32'h10408000;
      13239: inst = 32'hc405502;
      13240: inst = 32'h8220000;
      13241: inst = 32'h10408000;
      13242: inst = 32'hc40551d;
      13243: inst = 32'h8220000;
      13244: inst = 32'h10408000;
      13245: inst = 32'hc405521;
      13246: inst = 32'h8220000;
      13247: inst = 32'h10408000;
      13248: inst = 32'hc405522;
      13249: inst = 32'h8220000;
      13250: inst = 32'h10408000;
      13251: inst = 32'hc405523;
      13252: inst = 32'h8220000;
      13253: inst = 32'h10408000;
      13254: inst = 32'hc40555b;
      13255: inst = 32'h8220000;
      13256: inst = 32'h10408000;
      13257: inst = 32'hc40555c;
      13258: inst = 32'h8220000;
      13259: inst = 32'h10408000;
      13260: inst = 32'hc40555d;
      13261: inst = 32'h8220000;
      13262: inst = 32'h10408000;
      13263: inst = 32'hc405562;
      13264: inst = 32'h8220000;
      13265: inst = 32'h10408000;
      13266: inst = 32'hc40557d;
      13267: inst = 32'h8220000;
      13268: inst = 32'h10408000;
      13269: inst = 32'hc405582;
      13270: inst = 32'h8220000;
      13271: inst = 32'h10408000;
      13272: inst = 32'hc405583;
      13273: inst = 32'h8220000;
      13274: inst = 32'h10408000;
      13275: inst = 32'hc405584;
      13276: inst = 32'h8220000;
      13277: inst = 32'h10408000;
      13278: inst = 32'hc4055ba;
      13279: inst = 32'h8220000;
      13280: inst = 32'h10408000;
      13281: inst = 32'hc4055bb;
      13282: inst = 32'h8220000;
      13283: inst = 32'h10408000;
      13284: inst = 32'hc4055bc;
      13285: inst = 32'h8220000;
      13286: inst = 32'h10408000;
      13287: inst = 32'hc4055bd;
      13288: inst = 32'h8220000;
      13289: inst = 32'h10408000;
      13290: inst = 32'hc4055c2;
      13291: inst = 32'h8220000;
      13292: inst = 32'h10408000;
      13293: inst = 32'hc4055dd;
      13294: inst = 32'h8220000;
      13295: inst = 32'h10408000;
      13296: inst = 32'hc4055e2;
      13297: inst = 32'h8220000;
      13298: inst = 32'h10408000;
      13299: inst = 32'hc4055e3;
      13300: inst = 32'h8220000;
      13301: inst = 32'h10408000;
      13302: inst = 32'hc4055e4;
      13303: inst = 32'h8220000;
      13304: inst = 32'h10408000;
      13305: inst = 32'hc4055e5;
      13306: inst = 32'h8220000;
      13307: inst = 32'h10408000;
      13308: inst = 32'hc40561a;
      13309: inst = 32'h8220000;
      13310: inst = 32'h10408000;
      13311: inst = 32'hc40561b;
      13312: inst = 32'h8220000;
      13313: inst = 32'h10408000;
      13314: inst = 32'hc40561c;
      13315: inst = 32'h8220000;
      13316: inst = 32'h10408000;
      13317: inst = 32'hc40561d;
      13318: inst = 32'h8220000;
      13319: inst = 32'h10408000;
      13320: inst = 32'hc405642;
      13321: inst = 32'h8220000;
      13322: inst = 32'h10408000;
      13323: inst = 32'hc405643;
      13324: inst = 32'h8220000;
      13325: inst = 32'h10408000;
      13326: inst = 32'hc405644;
      13327: inst = 32'h8220000;
      13328: inst = 32'h10408000;
      13329: inst = 32'hc405645;
      13330: inst = 32'h8220000;
      13331: inst = 32'h10408000;
      13332: inst = 32'hc405679;
      13333: inst = 32'h8220000;
      13334: inst = 32'h10408000;
      13335: inst = 32'hc40567a;
      13336: inst = 32'h8220000;
      13337: inst = 32'h10408000;
      13338: inst = 32'hc40567b;
      13339: inst = 32'h8220000;
      13340: inst = 32'h10408000;
      13341: inst = 32'hc40567c;
      13342: inst = 32'h8220000;
      13343: inst = 32'h10408000;
      13344: inst = 32'hc4056a3;
      13345: inst = 32'h8220000;
      13346: inst = 32'h10408000;
      13347: inst = 32'hc4056a4;
      13348: inst = 32'h8220000;
      13349: inst = 32'h10408000;
      13350: inst = 32'hc4056a5;
      13351: inst = 32'h8220000;
      13352: inst = 32'h10408000;
      13353: inst = 32'hc4056a6;
      13354: inst = 32'h8220000;
      13355: inst = 32'hc20e6d9;
      13356: inst = 32'h10408000;
      13357: inst = 32'hc404bef;
      13358: inst = 32'h8220000;
      13359: inst = 32'h10408000;
      13360: inst = 32'hc404c4e;
      13361: inst = 32'h8220000;
      13362: inst = 32'hc20eeb7;
      13363: inst = 32'h10408000;
      13364: inst = 32'hc404c47;
      13365: inst = 32'h8220000;
      13366: inst = 32'hc20d615;
      13367: inst = 32'h10408000;
      13368: inst = 32'hc404ca2;
      13369: inst = 32'h8220000;
      13370: inst = 32'h10408000;
      13371: inst = 32'hc404d00;
      13372: inst = 32'h8220000;
      13373: inst = 32'hc209c91;
      13374: inst = 32'h10408000;
      13375: inst = 32'hc404ca3;
      13376: inst = 32'h8220000;
      13377: inst = 32'h10408000;
      13378: inst = 32'hc404d01;
      13379: inst = 32'h8220000;
      13380: inst = 32'hc207bf0;
      13381: inst = 32'h10408000;
      13382: inst = 32'hc404ca4;
      13383: inst = 32'h8220000;
      13384: inst = 32'h10408000;
      13385: inst = 32'hc404ca5;
      13386: inst = 32'h8220000;
      13387: inst = 32'h10408000;
      13388: inst = 32'hc404ca6;
      13389: inst = 32'h8220000;
      13390: inst = 32'h10408000;
      13391: inst = 32'hc404ca7;
      13392: inst = 32'h8220000;
      13393: inst = 32'h10408000;
      13394: inst = 32'hc404d02;
      13395: inst = 32'h8220000;
      13396: inst = 32'h10408000;
      13397: inst = 32'hc404d03;
      13398: inst = 32'h8220000;
      13399: inst = 32'h10408000;
      13400: inst = 32'hc404d04;
      13401: inst = 32'h8220000;
      13402: inst = 32'h10408000;
      13403: inst = 32'hc404d05;
      13404: inst = 32'h8220000;
      13405: inst = 32'h10408000;
      13406: inst = 32'hc404d06;
      13407: inst = 32'h8220000;
      13408: inst = 32'h10408000;
      13409: inst = 32'hc404d07;
      13410: inst = 32'h8220000;
      13411: inst = 32'h10408000;
      13412: inst = 32'hc404d08;
      13413: inst = 32'h8220000;
      13414: inst = 32'h10408000;
      13415: inst = 32'hc404d09;
      13416: inst = 32'h8220000;
      13417: inst = 32'h10408000;
      13418: inst = 32'hc404d0a;
      13419: inst = 32'h8220000;
      13420: inst = 32'h10408000;
      13421: inst = 32'hc404d0b;
      13422: inst = 32'h8220000;
      13423: inst = 32'h10408000;
      13424: inst = 32'hc404d0c;
      13425: inst = 32'h8220000;
      13426: inst = 32'h10408000;
      13427: inst = 32'hc404d0d;
      13428: inst = 32'h8220000;
      13429: inst = 32'h10408000;
      13430: inst = 32'hc404d0e;
      13431: inst = 32'h8220000;
      13432: inst = 32'h10408000;
      13433: inst = 32'hc404d0f;
      13434: inst = 32'h8220000;
      13435: inst = 32'h10408000;
      13436: inst = 32'hc404d10;
      13437: inst = 32'h8220000;
      13438: inst = 32'h10408000;
      13439: inst = 32'hc404d11;
      13440: inst = 32'h8220000;
      13441: inst = 32'h10408000;
      13442: inst = 32'hc404d12;
      13443: inst = 32'h8220000;
      13444: inst = 32'h10408000;
      13445: inst = 32'hc404d13;
      13446: inst = 32'h8220000;
      13447: inst = 32'h10408000;
      13448: inst = 32'hc404d14;
      13449: inst = 32'h8220000;
      13450: inst = 32'h10408000;
      13451: inst = 32'hc4055c3;
      13452: inst = 32'h8220000;
      13453: inst = 32'h10408000;
      13454: inst = 32'hc4055dc;
      13455: inst = 32'h8220000;
      13456: inst = 32'hc20ad55;
      13457: inst = 32'h10408000;
      13458: inst = 32'hc404cad;
      13459: inst = 32'h8220000;
      13460: inst = 32'hc208410;
      13461: inst = 32'h10408000;
      13462: inst = 32'hc404cae;
      13463: inst = 32'h8220000;
      13464: inst = 32'h10408000;
      13465: inst = 32'hc404caf;
      13466: inst = 32'h8220000;
      13467: inst = 32'h10408000;
      13468: inst = 32'hc404cb0;
      13469: inst = 32'h8220000;
      13470: inst = 32'h10408000;
      13471: inst = 32'hc404cb1;
      13472: inst = 32'h8220000;
      13473: inst = 32'h10408000;
      13474: inst = 32'hc404cb2;
      13475: inst = 32'h8220000;
      13476: inst = 32'h10408000;
      13477: inst = 32'hc404cb3;
      13478: inst = 32'h8220000;
      13479: inst = 32'h10408000;
      13480: inst = 32'hc404cb4;
      13481: inst = 32'h8220000;
      13482: inst = 32'h10408000;
      13483: inst = 32'hc404cb5;
      13484: inst = 32'h8220000;
      13485: inst = 32'h10408000;
      13486: inst = 32'hc40537d;
      13487: inst = 32'h8220000;
      13488: inst = 32'h10408000;
      13489: inst = 32'hc405385;
      13490: inst = 32'h8220000;
      13491: inst = 32'h10408000;
      13492: inst = 32'hc40539a;
      13493: inst = 32'h8220000;
      13494: inst = 32'h10408000;
      13495: inst = 32'hc4053a2;
      13496: inst = 32'h8220000;
      13497: inst = 32'h10408000;
      13498: inst = 32'hc4054a4;
      13499: inst = 32'h8220000;
      13500: inst = 32'h10408000;
      13501: inst = 32'hc4054bb;
      13502: inst = 32'h8220000;
      13503: inst = 32'h10408000;
      13504: inst = 32'hc405741;
      13505: inst = 32'h8220000;
      13506: inst = 32'h10408000;
      13507: inst = 32'hc40575e;
      13508: inst = 32'h8220000;
      13509: inst = 32'hc209470;
      13510: inst = 32'h10408000;
      13511: inst = 32'hc404cb6;
      13512: inst = 32'h8220000;
      13513: inst = 32'h10408000;
      13514: inst = 32'hc404d15;
      13515: inst = 32'h8220000;
      13516: inst = 32'hc20a534;
      13517: inst = 32'h10408000;
      13518: inst = 32'hc404cfb;
      13519: inst = 32'h8220000;
      13520: inst = 32'hc208c51;
      13521: inst = 32'h10408000;
      13522: inst = 32'hc404cfc;
      13523: inst = 32'h8220000;
      13524: inst = 32'h10408000;
      13525: inst = 32'hc404cfd;
      13526: inst = 32'h8220000;
      13527: inst = 32'h10408000;
      13528: inst = 32'hc4053da;
      13529: inst = 32'h8220000;
      13530: inst = 32'h10408000;
      13531: inst = 32'hc4053dc;
      13532: inst = 32'h8220000;
      13533: inst = 32'h10408000;
      13534: inst = 32'hc405403;
      13535: inst = 32'h8220000;
      13536: inst = 32'h10408000;
      13537: inst = 32'hc405405;
      13538: inst = 32'h8220000;
      13539: inst = 32'h10408000;
      13540: inst = 32'hc4054fa;
      13541: inst = 32'h8220000;
      13542: inst = 32'h10408000;
      13543: inst = 32'hc405525;
      13544: inst = 32'h8220000;
      13545: inst = 32'h10408000;
      13546: inst = 32'hc405557;
      13547: inst = 32'h8220000;
      13548: inst = 32'h10408000;
      13549: inst = 32'hc40555f;
      13550: inst = 32'h8220000;
      13551: inst = 32'h10408000;
      13552: inst = 32'hc405580;
      13553: inst = 32'h8220000;
      13554: inst = 32'h10408000;
      13555: inst = 32'hc405588;
      13556: inst = 32'h8220000;
      13557: inst = 32'h10408000;
      13558: inst = 32'hc405618;
      13559: inst = 32'h8220000;
      13560: inst = 32'h10408000;
      13561: inst = 32'hc405627;
      13562: inst = 32'h8220000;
      13563: inst = 32'h10408000;
      13564: inst = 32'hc405638;
      13565: inst = 32'h8220000;
      13566: inst = 32'h10408000;
      13567: inst = 32'hc405647;
      13568: inst = 32'h8220000;
      13569: inst = 32'h10408000;
      13570: inst = 32'hc40570b;
      13571: inst = 32'h8220000;
      13572: inst = 32'hc206b6d;
      13573: inst = 32'h10408000;
      13574: inst = 32'hc404d16;
      13575: inst = 32'h8220000;
      13576: inst = 32'h10408000;
      13577: inst = 32'hc404d75;
      13578: inst = 32'h8220000;
      13579: inst = 32'h10408000;
      13580: inst = 32'hc404d76;
      13581: inst = 32'h8220000;
      13582: inst = 32'h10408000;
      13583: inst = 32'hc404dd5;
      13584: inst = 32'h8220000;
      13585: inst = 32'h10408000;
      13586: inst = 32'hc404dd6;
      13587: inst = 32'h8220000;
      13588: inst = 32'h10408000;
      13589: inst = 32'hc404e35;
      13590: inst = 32'h8220000;
      13591: inst = 32'h10408000;
      13592: inst = 32'hc404e36;
      13593: inst = 32'h8220000;
      13594: inst = 32'h10408000;
      13595: inst = 32'hc404e95;
      13596: inst = 32'h8220000;
      13597: inst = 32'h10408000;
      13598: inst = 32'hc404e96;
      13599: inst = 32'h8220000;
      13600: inst = 32'h10408000;
      13601: inst = 32'hc404ef5;
      13602: inst = 32'h8220000;
      13603: inst = 32'h10408000;
      13604: inst = 32'hc404ef6;
      13605: inst = 32'h8220000;
      13606: inst = 32'h10408000;
      13607: inst = 32'hc404f55;
      13608: inst = 32'h8220000;
      13609: inst = 32'h10408000;
      13610: inst = 32'hc404f56;
      13611: inst = 32'h8220000;
      13612: inst = 32'h10408000;
      13613: inst = 32'hc404fb5;
      13614: inst = 32'h8220000;
      13615: inst = 32'h10408000;
      13616: inst = 32'hc404fb6;
      13617: inst = 32'h8220000;
      13618: inst = 32'h10408000;
      13619: inst = 32'hc405015;
      13620: inst = 32'h8220000;
      13621: inst = 32'h10408000;
      13622: inst = 32'hc405016;
      13623: inst = 32'h8220000;
      13624: inst = 32'h10408000;
      13625: inst = 32'hc405075;
      13626: inst = 32'h8220000;
      13627: inst = 32'h10408000;
      13628: inst = 32'hc405076;
      13629: inst = 32'h8220000;
      13630: inst = 32'h10408000;
      13631: inst = 32'hc4050d5;
      13632: inst = 32'h8220000;
      13633: inst = 32'h10408000;
      13634: inst = 32'hc4050d6;
      13635: inst = 32'h8220000;
      13636: inst = 32'h10408000;
      13637: inst = 32'hc405135;
      13638: inst = 32'h8220000;
      13639: inst = 32'h10408000;
      13640: inst = 32'hc405136;
      13641: inst = 32'h8220000;
      13642: inst = 32'h10408000;
      13643: inst = 32'hc405195;
      13644: inst = 32'h8220000;
      13645: inst = 32'h10408000;
      13646: inst = 32'hc405196;
      13647: inst = 32'h8220000;
      13648: inst = 32'h10408000;
      13649: inst = 32'hc4051f5;
      13650: inst = 32'h8220000;
      13651: inst = 32'h10408000;
      13652: inst = 32'hc4051f6;
      13653: inst = 32'h8220000;
      13654: inst = 32'h10408000;
      13655: inst = 32'hc405255;
      13656: inst = 32'h8220000;
      13657: inst = 32'h10408000;
      13658: inst = 32'hc405256;
      13659: inst = 32'h8220000;
      13660: inst = 32'h10408000;
      13661: inst = 32'hc4052b5;
      13662: inst = 32'h8220000;
      13663: inst = 32'h10408000;
      13664: inst = 32'hc4052b6;
      13665: inst = 32'h8220000;
      13666: inst = 32'h10408000;
      13667: inst = 32'hc405325;
      13668: inst = 32'h8220000;
      13669: inst = 32'h10408000;
      13670: inst = 32'hc40533a;
      13671: inst = 32'h8220000;
      13672: inst = 32'hc20c638;
      13673: inst = 32'h10408000;
      13674: inst = 32'hc404d5b;
      13675: inst = 32'h8220000;
      13676: inst = 32'hc208c71;
      13677: inst = 32'h10408000;
      13678: inst = 32'hc404d60;
      13679: inst = 32'h8220000;
      13680: inst = 32'h10408000;
      13681: inst = 32'hc404d61;
      13682: inst = 32'h8220000;
      13683: inst = 32'h10408000;
      13684: inst = 32'hc404d62;
      13685: inst = 32'h8220000;
      13686: inst = 32'h10408000;
      13687: inst = 32'hc404d63;
      13688: inst = 32'h8220000;
      13689: inst = 32'h10408000;
      13690: inst = 32'hc404d64;
      13691: inst = 32'h8220000;
      13692: inst = 32'h10408000;
      13693: inst = 32'hc404d65;
      13694: inst = 32'h8220000;
      13695: inst = 32'h10408000;
      13696: inst = 32'hc404d66;
      13697: inst = 32'h8220000;
      13698: inst = 32'h10408000;
      13699: inst = 32'hc404d67;
      13700: inst = 32'h8220000;
      13701: inst = 32'h10408000;
      13702: inst = 32'hc404d68;
      13703: inst = 32'h8220000;
      13704: inst = 32'h10408000;
      13705: inst = 32'hc404d69;
      13706: inst = 32'h8220000;
      13707: inst = 32'h10408000;
      13708: inst = 32'hc404d6a;
      13709: inst = 32'h8220000;
      13710: inst = 32'h10408000;
      13711: inst = 32'hc404d6b;
      13712: inst = 32'h8220000;
      13713: inst = 32'h10408000;
      13714: inst = 32'hc404d6c;
      13715: inst = 32'h8220000;
      13716: inst = 32'h10408000;
      13717: inst = 32'hc404d6d;
      13718: inst = 32'h8220000;
      13719: inst = 32'h10408000;
      13720: inst = 32'hc404d6e;
      13721: inst = 32'h8220000;
      13722: inst = 32'h10408000;
      13723: inst = 32'hc404d6f;
      13724: inst = 32'h8220000;
      13725: inst = 32'h10408000;
      13726: inst = 32'hc404d70;
      13727: inst = 32'h8220000;
      13728: inst = 32'h10408000;
      13729: inst = 32'hc404d71;
      13730: inst = 32'h8220000;
      13731: inst = 32'h10408000;
      13732: inst = 32'hc404d72;
      13733: inst = 32'h8220000;
      13734: inst = 32'h10408000;
      13735: inst = 32'hc404d73;
      13736: inst = 32'h8220000;
      13737: inst = 32'h10408000;
      13738: inst = 32'hc404d74;
      13739: inst = 32'h8220000;
      13740: inst = 32'h10408000;
      13741: inst = 32'hc404dc0;
      13742: inst = 32'h8220000;
      13743: inst = 32'h10408000;
      13744: inst = 32'hc404dca;
      13745: inst = 32'h8220000;
      13746: inst = 32'h10408000;
      13747: inst = 32'hc404dd4;
      13748: inst = 32'h8220000;
      13749: inst = 32'h10408000;
      13750: inst = 32'hc404e20;
      13751: inst = 32'h8220000;
      13752: inst = 32'h10408000;
      13753: inst = 32'hc404e2a;
      13754: inst = 32'h8220000;
      13755: inst = 32'h10408000;
      13756: inst = 32'hc404e34;
      13757: inst = 32'h8220000;
      13758: inst = 32'h10408000;
      13759: inst = 32'hc404e80;
      13760: inst = 32'h8220000;
      13761: inst = 32'h10408000;
      13762: inst = 32'hc404e8a;
      13763: inst = 32'h8220000;
      13764: inst = 32'h10408000;
      13765: inst = 32'hc404e94;
      13766: inst = 32'h8220000;
      13767: inst = 32'h10408000;
      13768: inst = 32'hc404ee0;
      13769: inst = 32'h8220000;
      13770: inst = 32'h10408000;
      13771: inst = 32'hc404eea;
      13772: inst = 32'h8220000;
      13773: inst = 32'h10408000;
      13774: inst = 32'hc404ef4;
      13775: inst = 32'h8220000;
      13776: inst = 32'h10408000;
      13777: inst = 32'hc404f40;
      13778: inst = 32'h8220000;
      13779: inst = 32'h10408000;
      13780: inst = 32'hc404f4a;
      13781: inst = 32'h8220000;
      13782: inst = 32'h10408000;
      13783: inst = 32'hc404f54;
      13784: inst = 32'h8220000;
      13785: inst = 32'h10408000;
      13786: inst = 32'hc404fa0;
      13787: inst = 32'h8220000;
      13788: inst = 32'h10408000;
      13789: inst = 32'hc404faa;
      13790: inst = 32'h8220000;
      13791: inst = 32'h10408000;
      13792: inst = 32'hc404fb4;
      13793: inst = 32'h8220000;
      13794: inst = 32'h10408000;
      13795: inst = 32'hc405000;
      13796: inst = 32'h8220000;
      13797: inst = 32'h10408000;
      13798: inst = 32'hc40500a;
      13799: inst = 32'h8220000;
      13800: inst = 32'h10408000;
      13801: inst = 32'hc405014;
      13802: inst = 32'h8220000;
      13803: inst = 32'h10408000;
      13804: inst = 32'hc405060;
      13805: inst = 32'h8220000;
      13806: inst = 32'h10408000;
      13807: inst = 32'hc40506a;
      13808: inst = 32'h8220000;
      13809: inst = 32'h10408000;
      13810: inst = 32'hc405074;
      13811: inst = 32'h8220000;
      13812: inst = 32'h10408000;
      13813: inst = 32'hc4050c0;
      13814: inst = 32'h8220000;
      13815: inst = 32'h10408000;
      13816: inst = 32'hc4050ca;
      13817: inst = 32'h8220000;
      13818: inst = 32'h10408000;
      13819: inst = 32'hc4050d4;
      13820: inst = 32'h8220000;
      13821: inst = 32'h10408000;
      13822: inst = 32'hc405120;
      13823: inst = 32'h8220000;
      13824: inst = 32'h10408000;
      13825: inst = 32'hc40512a;
      13826: inst = 32'h8220000;
      13827: inst = 32'h10408000;
      13828: inst = 32'hc405134;
      13829: inst = 32'h8220000;
      13830: inst = 32'h10408000;
      13831: inst = 32'hc405180;
      13832: inst = 32'h8220000;
      13833: inst = 32'h10408000;
      13834: inst = 32'hc40518a;
      13835: inst = 32'h8220000;
      13836: inst = 32'h10408000;
      13837: inst = 32'hc405194;
      13838: inst = 32'h8220000;
      13839: inst = 32'h10408000;
      13840: inst = 32'hc4051a8;
      13841: inst = 32'h8220000;
      13842: inst = 32'h10408000;
      13843: inst = 32'hc4051a9;
      13844: inst = 32'h8220000;
      13845: inst = 32'h10408000;
      13846: inst = 32'hc4051b7;
      13847: inst = 32'h8220000;
      13848: inst = 32'h10408000;
      13849: inst = 32'hc4051e0;
      13850: inst = 32'h8220000;
      13851: inst = 32'h10408000;
      13852: inst = 32'hc4051ea;
      13853: inst = 32'h8220000;
      13854: inst = 32'h10408000;
      13855: inst = 32'hc4051f4;
      13856: inst = 32'h8220000;
      13857: inst = 32'h10408000;
      13858: inst = 32'hc405208;
      13859: inst = 32'h8220000;
      13860: inst = 32'h10408000;
      13861: inst = 32'hc405217;
      13862: inst = 32'h8220000;
      13863: inst = 32'h10408000;
      13864: inst = 32'hc405240;
      13865: inst = 32'h8220000;
      13866: inst = 32'h10408000;
      13867: inst = 32'hc40524a;
      13868: inst = 32'h8220000;
      13869: inst = 32'h10408000;
      13870: inst = 32'hc405254;
      13871: inst = 32'h8220000;
      13872: inst = 32'h10408000;
      13873: inst = 32'hc40525e;
      13874: inst = 32'h8220000;
      13875: inst = 32'h10408000;
      13876: inst = 32'hc405268;
      13877: inst = 32'h8220000;
      13878: inst = 32'h10408000;
      13879: inst = 32'hc405277;
      13880: inst = 32'h8220000;
      13881: inst = 32'h10408000;
      13882: inst = 32'hc405281;
      13883: inst = 32'h8220000;
      13884: inst = 32'h10408000;
      13885: inst = 32'hc4052a0;
      13886: inst = 32'h8220000;
      13887: inst = 32'h10408000;
      13888: inst = 32'hc4052a1;
      13889: inst = 32'h8220000;
      13890: inst = 32'h10408000;
      13891: inst = 32'hc4052a2;
      13892: inst = 32'h8220000;
      13893: inst = 32'h10408000;
      13894: inst = 32'hc4052a3;
      13895: inst = 32'h8220000;
      13896: inst = 32'h10408000;
      13897: inst = 32'hc4052a4;
      13898: inst = 32'h8220000;
      13899: inst = 32'h10408000;
      13900: inst = 32'hc4052a5;
      13901: inst = 32'h8220000;
      13902: inst = 32'h10408000;
      13903: inst = 32'hc4052a6;
      13904: inst = 32'h8220000;
      13905: inst = 32'h10408000;
      13906: inst = 32'hc4052a7;
      13907: inst = 32'h8220000;
      13908: inst = 32'h10408000;
      13909: inst = 32'hc4052a8;
      13910: inst = 32'h8220000;
      13911: inst = 32'h10408000;
      13912: inst = 32'hc4052a9;
      13913: inst = 32'h8220000;
      13914: inst = 32'h10408000;
      13915: inst = 32'hc4052aa;
      13916: inst = 32'h8220000;
      13917: inst = 32'h10408000;
      13918: inst = 32'hc4052ab;
      13919: inst = 32'h8220000;
      13920: inst = 32'h10408000;
      13921: inst = 32'hc4052ac;
      13922: inst = 32'h8220000;
      13923: inst = 32'h10408000;
      13924: inst = 32'hc4052ad;
      13925: inst = 32'h8220000;
      13926: inst = 32'h10408000;
      13927: inst = 32'hc4052ae;
      13928: inst = 32'h8220000;
      13929: inst = 32'h10408000;
      13930: inst = 32'hc4052af;
      13931: inst = 32'h8220000;
      13932: inst = 32'h10408000;
      13933: inst = 32'hc4052b0;
      13934: inst = 32'h8220000;
      13935: inst = 32'h10408000;
      13936: inst = 32'hc4052b1;
      13937: inst = 32'h8220000;
      13938: inst = 32'h10408000;
      13939: inst = 32'hc4052b2;
      13940: inst = 32'h8220000;
      13941: inst = 32'h10408000;
      13942: inst = 32'hc4052b3;
      13943: inst = 32'h8220000;
      13944: inst = 32'h10408000;
      13945: inst = 32'hc4052b4;
      13946: inst = 32'h8220000;
      13947: inst = 32'h10408000;
      13948: inst = 32'hc4052bd;
      13949: inst = 32'h8220000;
      13950: inst = 32'h10408000;
      13951: inst = 32'hc4052be;
      13952: inst = 32'h8220000;
      13953: inst = 32'h10408000;
      13954: inst = 32'hc4052c8;
      13955: inst = 32'h8220000;
      13956: inst = 32'h10408000;
      13957: inst = 32'hc4052d7;
      13958: inst = 32'h8220000;
      13959: inst = 32'h10408000;
      13960: inst = 32'hc4052e1;
      13961: inst = 32'h8220000;
      13962: inst = 32'h10408000;
      13963: inst = 32'hc4052e2;
      13964: inst = 32'h8220000;
      13965: inst = 32'h10408000;
      13966: inst = 32'hc40531c;
      13967: inst = 32'h8220000;
      13968: inst = 32'h10408000;
      13969: inst = 32'hc40531d;
      13970: inst = 32'h8220000;
      13971: inst = 32'h10408000;
      13972: inst = 32'hc40531e;
      13973: inst = 32'h8220000;
      13974: inst = 32'h10408000;
      13975: inst = 32'hc40531f;
      13976: inst = 32'h8220000;
      13977: inst = 32'h10408000;
      13978: inst = 32'hc405320;
      13979: inst = 32'h8220000;
      13980: inst = 32'h10408000;
      13981: inst = 32'hc405326;
      13982: inst = 32'h8220000;
      13983: inst = 32'h10408000;
      13984: inst = 32'hc405327;
      13985: inst = 32'h8220000;
      13986: inst = 32'h10408000;
      13987: inst = 32'hc405328;
      13988: inst = 32'h8220000;
      13989: inst = 32'h10408000;
      13990: inst = 32'hc405337;
      13991: inst = 32'h8220000;
      13992: inst = 32'h10408000;
      13993: inst = 32'hc405338;
      13994: inst = 32'h8220000;
      13995: inst = 32'h10408000;
      13996: inst = 32'hc405339;
      13997: inst = 32'h8220000;
      13998: inst = 32'h10408000;
      13999: inst = 32'hc40533f;
      14000: inst = 32'h8220000;
      14001: inst = 32'h10408000;
      14002: inst = 32'hc405340;
      14003: inst = 32'h8220000;
      14004: inst = 32'h10408000;
      14005: inst = 32'hc405341;
      14006: inst = 32'h8220000;
      14007: inst = 32'h10408000;
      14008: inst = 32'hc405342;
      14009: inst = 32'h8220000;
      14010: inst = 32'h10408000;
      14011: inst = 32'hc405343;
      14012: inst = 32'h8220000;
      14013: inst = 32'h10408000;
      14014: inst = 32'hc40537b;
      14015: inst = 32'h8220000;
      14016: inst = 32'h10408000;
      14017: inst = 32'hc40537c;
      14018: inst = 32'h8220000;
      14019: inst = 32'h10408000;
      14020: inst = 32'hc405386;
      14021: inst = 32'h8220000;
      14022: inst = 32'h10408000;
      14023: inst = 32'hc405387;
      14024: inst = 32'h8220000;
      14025: inst = 32'h10408000;
      14026: inst = 32'hc405388;
      14027: inst = 32'h8220000;
      14028: inst = 32'h10408000;
      14029: inst = 32'hc405397;
      14030: inst = 32'h8220000;
      14031: inst = 32'h10408000;
      14032: inst = 32'hc405398;
      14033: inst = 32'h8220000;
      14034: inst = 32'h10408000;
      14035: inst = 32'hc405399;
      14036: inst = 32'h8220000;
      14037: inst = 32'h10408000;
      14038: inst = 32'hc4053a3;
      14039: inst = 32'h8220000;
      14040: inst = 32'h10408000;
      14041: inst = 32'hc4053a4;
      14042: inst = 32'h8220000;
      14043: inst = 32'h10408000;
      14044: inst = 32'hc4053db;
      14045: inst = 32'h8220000;
      14046: inst = 32'h10408000;
      14047: inst = 32'hc4053e5;
      14048: inst = 32'h8220000;
      14049: inst = 32'h10408000;
      14050: inst = 32'hc4053e6;
      14051: inst = 32'h8220000;
      14052: inst = 32'h10408000;
      14053: inst = 32'hc4053e7;
      14054: inst = 32'h8220000;
      14055: inst = 32'h10408000;
      14056: inst = 32'hc4053f8;
      14057: inst = 32'h8220000;
      14058: inst = 32'h10408000;
      14059: inst = 32'hc4053f9;
      14060: inst = 32'h8220000;
      14061: inst = 32'h10408000;
      14062: inst = 32'hc4053fa;
      14063: inst = 32'h8220000;
      14064: inst = 32'h10408000;
      14065: inst = 32'hc405404;
      14066: inst = 32'h8220000;
      14067: inst = 32'h10408000;
      14068: inst = 32'hc40543a;
      14069: inst = 32'h8220000;
      14070: inst = 32'h10408000;
      14071: inst = 32'hc40543b;
      14072: inst = 32'h8220000;
      14073: inst = 32'h10408000;
      14074: inst = 32'hc405445;
      14075: inst = 32'h8220000;
      14076: inst = 32'h10408000;
      14077: inst = 32'hc405446;
      14078: inst = 32'h8220000;
      14079: inst = 32'h10408000;
      14080: inst = 32'hc405447;
      14081: inst = 32'h8220000;
      14082: inst = 32'h10408000;
      14083: inst = 32'hc405458;
      14084: inst = 32'h8220000;
      14085: inst = 32'h10408000;
      14086: inst = 32'hc405459;
      14087: inst = 32'h8220000;
      14088: inst = 32'h10408000;
      14089: inst = 32'hc40545a;
      14090: inst = 32'h8220000;
      14091: inst = 32'h10408000;
      14092: inst = 32'hc405464;
      14093: inst = 32'h8220000;
      14094: inst = 32'h10408000;
      14095: inst = 32'hc405465;
      14096: inst = 32'h8220000;
      14097: inst = 32'h10408000;
      14098: inst = 32'hc405499;
      14099: inst = 32'h8220000;
      14100: inst = 32'h10408000;
      14101: inst = 32'hc40549a;
      14102: inst = 32'h8220000;
      14103: inst = 32'h10408000;
      14104: inst = 32'hc4054a5;
      14105: inst = 32'h8220000;
      14106: inst = 32'h10408000;
      14107: inst = 32'hc4054a6;
      14108: inst = 32'h8220000;
      14109: inst = 32'h10408000;
      14110: inst = 32'hc4054a7;
      14111: inst = 32'h8220000;
      14112: inst = 32'h10408000;
      14113: inst = 32'hc4054b8;
      14114: inst = 32'h8220000;
      14115: inst = 32'h10408000;
      14116: inst = 32'hc4054b9;
      14117: inst = 32'h8220000;
      14118: inst = 32'h10408000;
      14119: inst = 32'hc4054ba;
      14120: inst = 32'h8220000;
      14121: inst = 32'h10408000;
      14122: inst = 32'hc4054c5;
      14123: inst = 32'h8220000;
      14124: inst = 32'h10408000;
      14125: inst = 32'hc4054c6;
      14126: inst = 32'h8220000;
      14127: inst = 32'h10408000;
      14128: inst = 32'hc4054f8;
      14129: inst = 32'h8220000;
      14130: inst = 32'h10408000;
      14131: inst = 32'hc4054f9;
      14132: inst = 32'h8220000;
      14133: inst = 32'h10408000;
      14134: inst = 32'hc405500;
      14135: inst = 32'h8220000;
      14136: inst = 32'h10408000;
      14137: inst = 32'hc405504;
      14138: inst = 32'h8220000;
      14139: inst = 32'h10408000;
      14140: inst = 32'hc405505;
      14141: inst = 32'h8220000;
      14142: inst = 32'h10408000;
      14143: inst = 32'hc405506;
      14144: inst = 32'h8220000;
      14145: inst = 32'h10408000;
      14146: inst = 32'hc405507;
      14147: inst = 32'h8220000;
      14148: inst = 32'h10408000;
      14149: inst = 32'hc405518;
      14150: inst = 32'h8220000;
      14151: inst = 32'h10408000;
      14152: inst = 32'hc405519;
      14153: inst = 32'h8220000;
      14154: inst = 32'h10408000;
      14155: inst = 32'hc40551a;
      14156: inst = 32'h8220000;
      14157: inst = 32'h10408000;
      14158: inst = 32'hc40551b;
      14159: inst = 32'h8220000;
      14160: inst = 32'h10408000;
      14161: inst = 32'hc40551f;
      14162: inst = 32'h8220000;
      14163: inst = 32'h10408000;
      14164: inst = 32'hc405526;
      14165: inst = 32'h8220000;
      14166: inst = 32'h10408000;
      14167: inst = 32'hc405527;
      14168: inst = 32'h8220000;
      14169: inst = 32'h10408000;
      14170: inst = 32'hc405558;
      14171: inst = 32'h8220000;
      14172: inst = 32'h10408000;
      14173: inst = 32'hc405559;
      14174: inst = 32'h8220000;
      14175: inst = 32'h10408000;
      14176: inst = 32'hc405560;
      14177: inst = 32'h8220000;
      14178: inst = 32'h10408000;
      14179: inst = 32'hc405564;
      14180: inst = 32'h8220000;
      14181: inst = 32'h10408000;
      14182: inst = 32'hc405565;
      14183: inst = 32'h8220000;
      14184: inst = 32'h10408000;
      14185: inst = 32'hc405566;
      14186: inst = 32'h8220000;
      14187: inst = 32'h10408000;
      14188: inst = 32'hc405567;
      14189: inst = 32'h8220000;
      14190: inst = 32'h10408000;
      14191: inst = 32'hc405578;
      14192: inst = 32'h8220000;
      14193: inst = 32'h10408000;
      14194: inst = 32'hc405579;
      14195: inst = 32'h8220000;
      14196: inst = 32'h10408000;
      14197: inst = 32'hc40557a;
      14198: inst = 32'h8220000;
      14199: inst = 32'h10408000;
      14200: inst = 32'hc40557b;
      14201: inst = 32'h8220000;
      14202: inst = 32'h10408000;
      14203: inst = 32'hc40557f;
      14204: inst = 32'h8220000;
      14205: inst = 32'h10408000;
      14206: inst = 32'hc405586;
      14207: inst = 32'h8220000;
      14208: inst = 32'h10408000;
      14209: inst = 32'hc405587;
      14210: inst = 32'h8220000;
      14211: inst = 32'h10408000;
      14212: inst = 32'hc4055b7;
      14213: inst = 32'h8220000;
      14214: inst = 32'h10408000;
      14215: inst = 32'hc4055b8;
      14216: inst = 32'h8220000;
      14217: inst = 32'h10408000;
      14218: inst = 32'hc4055bf;
      14219: inst = 32'h8220000;
      14220: inst = 32'h10408000;
      14221: inst = 32'hc4055c0;
      14222: inst = 32'h8220000;
      14223: inst = 32'h10408000;
      14224: inst = 32'hc4055c4;
      14225: inst = 32'h8220000;
      14226: inst = 32'h10408000;
      14227: inst = 32'hc4055c5;
      14228: inst = 32'h8220000;
      14229: inst = 32'h10408000;
      14230: inst = 32'hc4055c6;
      14231: inst = 32'h8220000;
      14232: inst = 32'h10408000;
      14233: inst = 32'hc4055c7;
      14234: inst = 32'h8220000;
      14235: inst = 32'h10408000;
      14236: inst = 32'hc4055d8;
      14237: inst = 32'h8220000;
      14238: inst = 32'h10408000;
      14239: inst = 32'hc4055d9;
      14240: inst = 32'h8220000;
      14241: inst = 32'h10408000;
      14242: inst = 32'hc4055da;
      14243: inst = 32'h8220000;
      14244: inst = 32'h10408000;
      14245: inst = 32'hc4055db;
      14246: inst = 32'h8220000;
      14247: inst = 32'h10408000;
      14248: inst = 32'hc4055df;
      14249: inst = 32'h8220000;
      14250: inst = 32'h10408000;
      14251: inst = 32'hc4055e0;
      14252: inst = 32'h8220000;
      14253: inst = 32'h10408000;
      14254: inst = 32'hc4055e7;
      14255: inst = 32'h8220000;
      14256: inst = 32'h10408000;
      14257: inst = 32'hc4055e8;
      14258: inst = 32'h8220000;
      14259: inst = 32'h10408000;
      14260: inst = 32'hc405616;
      14261: inst = 32'h8220000;
      14262: inst = 32'h10408000;
      14263: inst = 32'hc405617;
      14264: inst = 32'h8220000;
      14265: inst = 32'h10408000;
      14266: inst = 32'hc40561f;
      14267: inst = 32'h8220000;
      14268: inst = 32'h10408000;
      14269: inst = 32'hc405620;
      14270: inst = 32'h8220000;
      14271: inst = 32'h10408000;
      14272: inst = 32'hc405623;
      14273: inst = 32'h8220000;
      14274: inst = 32'h10408000;
      14275: inst = 32'hc405624;
      14276: inst = 32'h8220000;
      14277: inst = 32'h10408000;
      14278: inst = 32'hc405625;
      14279: inst = 32'h8220000;
      14280: inst = 32'h10408000;
      14281: inst = 32'hc405626;
      14282: inst = 32'h8220000;
      14283: inst = 32'h10408000;
      14284: inst = 32'hc405639;
      14285: inst = 32'h8220000;
      14286: inst = 32'h10408000;
      14287: inst = 32'hc40563a;
      14288: inst = 32'h8220000;
      14289: inst = 32'h10408000;
      14290: inst = 32'hc40563b;
      14291: inst = 32'h8220000;
      14292: inst = 32'h10408000;
      14293: inst = 32'hc40563c;
      14294: inst = 32'h8220000;
      14295: inst = 32'h10408000;
      14296: inst = 32'hc40563f;
      14297: inst = 32'h8220000;
      14298: inst = 32'h10408000;
      14299: inst = 32'hc405640;
      14300: inst = 32'h8220000;
      14301: inst = 32'h10408000;
      14302: inst = 32'hc405648;
      14303: inst = 32'h8220000;
      14304: inst = 32'h10408000;
      14305: inst = 32'hc405649;
      14306: inst = 32'h8220000;
      14307: inst = 32'h10408000;
      14308: inst = 32'hc405675;
      14309: inst = 32'h8220000;
      14310: inst = 32'h10408000;
      14311: inst = 32'hc405676;
      14312: inst = 32'h8220000;
      14313: inst = 32'h10408000;
      14314: inst = 32'hc405677;
      14315: inst = 32'h8220000;
      14316: inst = 32'h10408000;
      14317: inst = 32'hc40567e;
      14318: inst = 32'h8220000;
      14319: inst = 32'h10408000;
      14320: inst = 32'hc40567f;
      14321: inst = 32'h8220000;
      14322: inst = 32'h10408000;
      14323: inst = 32'hc405680;
      14324: inst = 32'h8220000;
      14325: inst = 32'h10408000;
      14326: inst = 32'hc405683;
      14327: inst = 32'h8220000;
      14328: inst = 32'h10408000;
      14329: inst = 32'hc405684;
      14330: inst = 32'h8220000;
      14331: inst = 32'h10408000;
      14332: inst = 32'hc405685;
      14333: inst = 32'h8220000;
      14334: inst = 32'h10408000;
      14335: inst = 32'hc405686;
      14336: inst = 32'h8220000;
      14337: inst = 32'h10408000;
      14338: inst = 32'hc405699;
      14339: inst = 32'h8220000;
      14340: inst = 32'h10408000;
      14341: inst = 32'hc40569a;
      14342: inst = 32'h8220000;
      14343: inst = 32'h10408000;
      14344: inst = 32'hc40569b;
      14345: inst = 32'h8220000;
      14346: inst = 32'h10408000;
      14347: inst = 32'hc40569c;
      14348: inst = 32'h8220000;
      14349: inst = 32'h10408000;
      14350: inst = 32'hc40569f;
      14351: inst = 32'h8220000;
      14352: inst = 32'h10408000;
      14353: inst = 32'hc4056a0;
      14354: inst = 32'h8220000;
      14355: inst = 32'h10408000;
      14356: inst = 32'hc4056a1;
      14357: inst = 32'h8220000;
      14358: inst = 32'h10408000;
      14359: inst = 32'hc4056a8;
      14360: inst = 32'h8220000;
      14361: inst = 32'h10408000;
      14362: inst = 32'hc4056a9;
      14363: inst = 32'h8220000;
      14364: inst = 32'h10408000;
      14365: inst = 32'hc4056aa;
      14366: inst = 32'h8220000;
      14367: inst = 32'h10408000;
      14368: inst = 32'hc4056d4;
      14369: inst = 32'h8220000;
      14370: inst = 32'h10408000;
      14371: inst = 32'hc4056d5;
      14372: inst = 32'h8220000;
      14373: inst = 32'h10408000;
      14374: inst = 32'hc4056d6;
      14375: inst = 32'h8220000;
      14376: inst = 32'h10408000;
      14377: inst = 32'hc4056d7;
      14378: inst = 32'h8220000;
      14379: inst = 32'h10408000;
      14380: inst = 32'hc4056d8;
      14381: inst = 32'h8220000;
      14382: inst = 32'h10408000;
      14383: inst = 32'hc4056d9;
      14384: inst = 32'h8220000;
      14385: inst = 32'h10408000;
      14386: inst = 32'hc4056da;
      14387: inst = 32'h8220000;
      14388: inst = 32'h10408000;
      14389: inst = 32'hc4056db;
      14390: inst = 32'h8220000;
      14391: inst = 32'h10408000;
      14392: inst = 32'hc4056dc;
      14393: inst = 32'h8220000;
      14394: inst = 32'h10408000;
      14395: inst = 32'hc4056dd;
      14396: inst = 32'h8220000;
      14397: inst = 32'h10408000;
      14398: inst = 32'hc4056de;
      14399: inst = 32'h8220000;
      14400: inst = 32'h10408000;
      14401: inst = 32'hc4056df;
      14402: inst = 32'h8220000;
      14403: inst = 32'h10408000;
      14404: inst = 32'hc4056e0;
      14405: inst = 32'h8220000;
      14406: inst = 32'h10408000;
      14407: inst = 32'hc4056e3;
      14408: inst = 32'h8220000;
      14409: inst = 32'h10408000;
      14410: inst = 32'hc4056e4;
      14411: inst = 32'h8220000;
      14412: inst = 32'h10408000;
      14413: inst = 32'hc4056e5;
      14414: inst = 32'h8220000;
      14415: inst = 32'h10408000;
      14416: inst = 32'hc4056e6;
      14417: inst = 32'h8220000;
      14418: inst = 32'h10408000;
      14419: inst = 32'hc4056f9;
      14420: inst = 32'h8220000;
      14421: inst = 32'h10408000;
      14422: inst = 32'hc4056fa;
      14423: inst = 32'h8220000;
      14424: inst = 32'h10408000;
      14425: inst = 32'hc4056fb;
      14426: inst = 32'h8220000;
      14427: inst = 32'h10408000;
      14428: inst = 32'hc4056fc;
      14429: inst = 32'h8220000;
      14430: inst = 32'h10408000;
      14431: inst = 32'hc4056ff;
      14432: inst = 32'h8220000;
      14433: inst = 32'h10408000;
      14434: inst = 32'hc405700;
      14435: inst = 32'h8220000;
      14436: inst = 32'h10408000;
      14437: inst = 32'hc405701;
      14438: inst = 32'h8220000;
      14439: inst = 32'h10408000;
      14440: inst = 32'hc405702;
      14441: inst = 32'h8220000;
      14442: inst = 32'h10408000;
      14443: inst = 32'hc405703;
      14444: inst = 32'h8220000;
      14445: inst = 32'h10408000;
      14446: inst = 32'hc405704;
      14447: inst = 32'h8220000;
      14448: inst = 32'h10408000;
      14449: inst = 32'hc405705;
      14450: inst = 32'h8220000;
      14451: inst = 32'h10408000;
      14452: inst = 32'hc405706;
      14453: inst = 32'h8220000;
      14454: inst = 32'h10408000;
      14455: inst = 32'hc405707;
      14456: inst = 32'h8220000;
      14457: inst = 32'h10408000;
      14458: inst = 32'hc405708;
      14459: inst = 32'h8220000;
      14460: inst = 32'h10408000;
      14461: inst = 32'hc405709;
      14462: inst = 32'h8220000;
      14463: inst = 32'h10408000;
      14464: inst = 32'hc40570a;
      14465: inst = 32'h8220000;
      14466: inst = 32'h10408000;
      14467: inst = 32'hc405734;
      14468: inst = 32'h8220000;
      14469: inst = 32'h10408000;
      14470: inst = 32'hc405735;
      14471: inst = 32'h8220000;
      14472: inst = 32'h10408000;
      14473: inst = 32'hc405736;
      14474: inst = 32'h8220000;
      14475: inst = 32'h10408000;
      14476: inst = 32'hc405737;
      14477: inst = 32'h8220000;
      14478: inst = 32'h10408000;
      14479: inst = 32'hc405738;
      14480: inst = 32'h8220000;
      14481: inst = 32'h10408000;
      14482: inst = 32'hc405739;
      14483: inst = 32'h8220000;
      14484: inst = 32'h10408000;
      14485: inst = 32'hc40573a;
      14486: inst = 32'h8220000;
      14487: inst = 32'h10408000;
      14488: inst = 32'hc40573b;
      14489: inst = 32'h8220000;
      14490: inst = 32'h10408000;
      14491: inst = 32'hc40573c;
      14492: inst = 32'h8220000;
      14493: inst = 32'h10408000;
      14494: inst = 32'hc40573d;
      14495: inst = 32'h8220000;
      14496: inst = 32'h10408000;
      14497: inst = 32'hc40573e;
      14498: inst = 32'h8220000;
      14499: inst = 32'h10408000;
      14500: inst = 32'hc40573f;
      14501: inst = 32'h8220000;
      14502: inst = 32'h10408000;
      14503: inst = 32'hc405740;
      14504: inst = 32'h8220000;
      14505: inst = 32'h10408000;
      14506: inst = 32'hc405742;
      14507: inst = 32'h8220000;
      14508: inst = 32'h10408000;
      14509: inst = 32'hc405743;
      14510: inst = 32'h8220000;
      14511: inst = 32'h10408000;
      14512: inst = 32'hc405744;
      14513: inst = 32'h8220000;
      14514: inst = 32'h10408000;
      14515: inst = 32'hc405745;
      14516: inst = 32'h8220000;
      14517: inst = 32'h10408000;
      14518: inst = 32'hc405746;
      14519: inst = 32'h8220000;
      14520: inst = 32'h10408000;
      14521: inst = 32'hc405759;
      14522: inst = 32'h8220000;
      14523: inst = 32'h10408000;
      14524: inst = 32'hc40575a;
      14525: inst = 32'h8220000;
      14526: inst = 32'h10408000;
      14527: inst = 32'hc40575b;
      14528: inst = 32'h8220000;
      14529: inst = 32'h10408000;
      14530: inst = 32'hc40575c;
      14531: inst = 32'h8220000;
      14532: inst = 32'h10408000;
      14533: inst = 32'hc40575d;
      14534: inst = 32'h8220000;
      14535: inst = 32'h10408000;
      14536: inst = 32'hc40575f;
      14537: inst = 32'h8220000;
      14538: inst = 32'h10408000;
      14539: inst = 32'hc405760;
      14540: inst = 32'h8220000;
      14541: inst = 32'h10408000;
      14542: inst = 32'hc405761;
      14543: inst = 32'h8220000;
      14544: inst = 32'h10408000;
      14545: inst = 32'hc405762;
      14546: inst = 32'h8220000;
      14547: inst = 32'h10408000;
      14548: inst = 32'hc405763;
      14549: inst = 32'h8220000;
      14550: inst = 32'h10408000;
      14551: inst = 32'hc405764;
      14552: inst = 32'h8220000;
      14553: inst = 32'h10408000;
      14554: inst = 32'hc405765;
      14555: inst = 32'h8220000;
      14556: inst = 32'h10408000;
      14557: inst = 32'hc405766;
      14558: inst = 32'h8220000;
      14559: inst = 32'h10408000;
      14560: inst = 32'hc405767;
      14561: inst = 32'h8220000;
      14562: inst = 32'h10408000;
      14563: inst = 32'hc405768;
      14564: inst = 32'h8220000;
      14565: inst = 32'h10408000;
      14566: inst = 32'hc405769;
      14567: inst = 32'h8220000;
      14568: inst = 32'h10408000;
      14569: inst = 32'hc40576a;
      14570: inst = 32'h8220000;
      14571: inst = 32'h10408000;
      14572: inst = 32'hc40576b;
      14573: inst = 32'h8220000;
      14574: inst = 32'h10408000;
      14575: inst = 32'hc405793;
      14576: inst = 32'h8220000;
      14577: inst = 32'h10408000;
      14578: inst = 32'hc405794;
      14579: inst = 32'h8220000;
      14580: inst = 32'h10408000;
      14581: inst = 32'hc405795;
      14582: inst = 32'h8220000;
      14583: inst = 32'h10408000;
      14584: inst = 32'hc405796;
      14585: inst = 32'h8220000;
      14586: inst = 32'h10408000;
      14587: inst = 32'hc405797;
      14588: inst = 32'h8220000;
      14589: inst = 32'h10408000;
      14590: inst = 32'hc405798;
      14591: inst = 32'h8220000;
      14592: inst = 32'h10408000;
      14593: inst = 32'hc405799;
      14594: inst = 32'h8220000;
      14595: inst = 32'h10408000;
      14596: inst = 32'hc40579a;
      14597: inst = 32'h8220000;
      14598: inst = 32'h10408000;
      14599: inst = 32'hc40579b;
      14600: inst = 32'h8220000;
      14601: inst = 32'h10408000;
      14602: inst = 32'hc40579c;
      14603: inst = 32'h8220000;
      14604: inst = 32'h10408000;
      14605: inst = 32'hc40579d;
      14606: inst = 32'h8220000;
      14607: inst = 32'h10408000;
      14608: inst = 32'hc40579e;
      14609: inst = 32'h8220000;
      14610: inst = 32'h10408000;
      14611: inst = 32'hc40579f;
      14612: inst = 32'h8220000;
      14613: inst = 32'h10408000;
      14614: inst = 32'hc4057a0;
      14615: inst = 32'h8220000;
      14616: inst = 32'h10408000;
      14617: inst = 32'hc4057a1;
      14618: inst = 32'h8220000;
      14619: inst = 32'h10408000;
      14620: inst = 32'hc4057a2;
      14621: inst = 32'h8220000;
      14622: inst = 32'h10408000;
      14623: inst = 32'hc4057a3;
      14624: inst = 32'h8220000;
      14625: inst = 32'h10408000;
      14626: inst = 32'hc4057a4;
      14627: inst = 32'h8220000;
      14628: inst = 32'h10408000;
      14629: inst = 32'hc4057a5;
      14630: inst = 32'h8220000;
      14631: inst = 32'h10408000;
      14632: inst = 32'hc4057a6;
      14633: inst = 32'h8220000;
      14634: inst = 32'h10408000;
      14635: inst = 32'hc4057b9;
      14636: inst = 32'h8220000;
      14637: inst = 32'h10408000;
      14638: inst = 32'hc4057ba;
      14639: inst = 32'h8220000;
      14640: inst = 32'h10408000;
      14641: inst = 32'hc4057bb;
      14642: inst = 32'h8220000;
      14643: inst = 32'h10408000;
      14644: inst = 32'hc4057bc;
      14645: inst = 32'h8220000;
      14646: inst = 32'h10408000;
      14647: inst = 32'hc4057bd;
      14648: inst = 32'h8220000;
      14649: inst = 32'h10408000;
      14650: inst = 32'hc4057be;
      14651: inst = 32'h8220000;
      14652: inst = 32'h10408000;
      14653: inst = 32'hc4057bf;
      14654: inst = 32'h8220000;
      14655: inst = 32'h10408000;
      14656: inst = 32'hc4057c0;
      14657: inst = 32'h8220000;
      14658: inst = 32'h10408000;
      14659: inst = 32'hc4057c1;
      14660: inst = 32'h8220000;
      14661: inst = 32'h10408000;
      14662: inst = 32'hc4057c2;
      14663: inst = 32'h8220000;
      14664: inst = 32'h10408000;
      14665: inst = 32'hc4057c3;
      14666: inst = 32'h8220000;
      14667: inst = 32'h10408000;
      14668: inst = 32'hc4057c4;
      14669: inst = 32'h8220000;
      14670: inst = 32'h10408000;
      14671: inst = 32'hc4057c5;
      14672: inst = 32'h8220000;
      14673: inst = 32'h10408000;
      14674: inst = 32'hc4057c6;
      14675: inst = 32'h8220000;
      14676: inst = 32'h10408000;
      14677: inst = 32'hc4057c7;
      14678: inst = 32'h8220000;
      14679: inst = 32'h10408000;
      14680: inst = 32'hc4057c8;
      14681: inst = 32'h8220000;
      14682: inst = 32'h10408000;
      14683: inst = 32'hc4057c9;
      14684: inst = 32'h8220000;
      14685: inst = 32'h10408000;
      14686: inst = 32'hc4057ca;
      14687: inst = 32'h8220000;
      14688: inst = 32'h10408000;
      14689: inst = 32'hc4057cb;
      14690: inst = 32'h8220000;
      14691: inst = 32'h10408000;
      14692: inst = 32'hc4057cc;
      14693: inst = 32'h8220000;
      14694: inst = 32'hc20bdd7;
      14695: inst = 32'h10408000;
      14696: inst = 32'hc404dc1;
      14697: inst = 32'h8220000;
      14698: inst = 32'h10408000;
      14699: inst = 32'hc404dc2;
      14700: inst = 32'h8220000;
      14701: inst = 32'h10408000;
      14702: inst = 32'hc404dc3;
      14703: inst = 32'h8220000;
      14704: inst = 32'h10408000;
      14705: inst = 32'hc404dc4;
      14706: inst = 32'h8220000;
      14707: inst = 32'h10408000;
      14708: inst = 32'hc404dc5;
      14709: inst = 32'h8220000;
      14710: inst = 32'h10408000;
      14711: inst = 32'hc404dc6;
      14712: inst = 32'h8220000;
      14713: inst = 32'h10408000;
      14714: inst = 32'hc404dc7;
      14715: inst = 32'h8220000;
      14716: inst = 32'h10408000;
      14717: inst = 32'hc404dc8;
      14718: inst = 32'h8220000;
      14719: inst = 32'h10408000;
      14720: inst = 32'hc404dc9;
      14721: inst = 32'h8220000;
      14722: inst = 32'h10408000;
      14723: inst = 32'hc404dcb;
      14724: inst = 32'h8220000;
      14725: inst = 32'h10408000;
      14726: inst = 32'hc404dcc;
      14727: inst = 32'h8220000;
      14728: inst = 32'h10408000;
      14729: inst = 32'hc404dcd;
      14730: inst = 32'h8220000;
      14731: inst = 32'h10408000;
      14732: inst = 32'hc404dce;
      14733: inst = 32'h8220000;
      14734: inst = 32'h10408000;
      14735: inst = 32'hc404dcf;
      14736: inst = 32'h8220000;
      14737: inst = 32'h10408000;
      14738: inst = 32'hc404dd0;
      14739: inst = 32'h8220000;
      14740: inst = 32'h10408000;
      14741: inst = 32'hc404dd1;
      14742: inst = 32'h8220000;
      14743: inst = 32'h10408000;
      14744: inst = 32'hc404dd2;
      14745: inst = 32'h8220000;
      14746: inst = 32'h10408000;
      14747: inst = 32'hc404dd3;
      14748: inst = 32'h8220000;
      14749: inst = 32'h10408000;
      14750: inst = 32'hc404e21;
      14751: inst = 32'h8220000;
      14752: inst = 32'h10408000;
      14753: inst = 32'hc404e22;
      14754: inst = 32'h8220000;
      14755: inst = 32'h10408000;
      14756: inst = 32'hc404e23;
      14757: inst = 32'h8220000;
      14758: inst = 32'h10408000;
      14759: inst = 32'hc404e24;
      14760: inst = 32'h8220000;
      14761: inst = 32'h10408000;
      14762: inst = 32'hc404e25;
      14763: inst = 32'h8220000;
      14764: inst = 32'h10408000;
      14765: inst = 32'hc404e26;
      14766: inst = 32'h8220000;
      14767: inst = 32'h10408000;
      14768: inst = 32'hc404e27;
      14769: inst = 32'h8220000;
      14770: inst = 32'h10408000;
      14771: inst = 32'hc404e28;
      14772: inst = 32'h8220000;
      14773: inst = 32'h10408000;
      14774: inst = 32'hc404e29;
      14775: inst = 32'h8220000;
      14776: inst = 32'h10408000;
      14777: inst = 32'hc404e2b;
      14778: inst = 32'h8220000;
      14779: inst = 32'h10408000;
      14780: inst = 32'hc404e2c;
      14781: inst = 32'h8220000;
      14782: inst = 32'h10408000;
      14783: inst = 32'hc404e2d;
      14784: inst = 32'h8220000;
      14785: inst = 32'h10408000;
      14786: inst = 32'hc404e2e;
      14787: inst = 32'h8220000;
      14788: inst = 32'h10408000;
      14789: inst = 32'hc404e2f;
      14790: inst = 32'h8220000;
      14791: inst = 32'h10408000;
      14792: inst = 32'hc404e30;
      14793: inst = 32'h8220000;
      14794: inst = 32'h10408000;
      14795: inst = 32'hc404e31;
      14796: inst = 32'h8220000;
      14797: inst = 32'h10408000;
      14798: inst = 32'hc404e32;
      14799: inst = 32'h8220000;
      14800: inst = 32'h10408000;
      14801: inst = 32'hc404e33;
      14802: inst = 32'h8220000;
      14803: inst = 32'h10408000;
      14804: inst = 32'hc404e81;
      14805: inst = 32'h8220000;
      14806: inst = 32'h10408000;
      14807: inst = 32'hc404e82;
      14808: inst = 32'h8220000;
      14809: inst = 32'h10408000;
      14810: inst = 32'hc404e83;
      14811: inst = 32'h8220000;
      14812: inst = 32'h10408000;
      14813: inst = 32'hc404e84;
      14814: inst = 32'h8220000;
      14815: inst = 32'h10408000;
      14816: inst = 32'hc404e85;
      14817: inst = 32'h8220000;
      14818: inst = 32'h10408000;
      14819: inst = 32'hc404e86;
      14820: inst = 32'h8220000;
      14821: inst = 32'h10408000;
      14822: inst = 32'hc404e87;
      14823: inst = 32'h8220000;
      14824: inst = 32'h10408000;
      14825: inst = 32'hc404e88;
      14826: inst = 32'h8220000;
      14827: inst = 32'h10408000;
      14828: inst = 32'hc404e89;
      14829: inst = 32'h8220000;
      14830: inst = 32'h10408000;
      14831: inst = 32'hc404e8b;
      14832: inst = 32'h8220000;
      14833: inst = 32'h10408000;
      14834: inst = 32'hc404e8c;
      14835: inst = 32'h8220000;
      14836: inst = 32'h10408000;
      14837: inst = 32'hc404e8d;
      14838: inst = 32'h8220000;
      14839: inst = 32'h10408000;
      14840: inst = 32'hc404e8e;
      14841: inst = 32'h8220000;
      14842: inst = 32'h10408000;
      14843: inst = 32'hc404e8f;
      14844: inst = 32'h8220000;
      14845: inst = 32'h10408000;
      14846: inst = 32'hc404e90;
      14847: inst = 32'h8220000;
      14848: inst = 32'h10408000;
      14849: inst = 32'hc404e91;
      14850: inst = 32'h8220000;
      14851: inst = 32'h10408000;
      14852: inst = 32'hc404e92;
      14853: inst = 32'h8220000;
      14854: inst = 32'h10408000;
      14855: inst = 32'hc404e93;
      14856: inst = 32'h8220000;
      14857: inst = 32'h10408000;
      14858: inst = 32'hc404ee1;
      14859: inst = 32'h8220000;
      14860: inst = 32'h10408000;
      14861: inst = 32'hc404ee2;
      14862: inst = 32'h8220000;
      14863: inst = 32'h10408000;
      14864: inst = 32'hc404ee3;
      14865: inst = 32'h8220000;
      14866: inst = 32'h10408000;
      14867: inst = 32'hc404ee4;
      14868: inst = 32'h8220000;
      14869: inst = 32'h10408000;
      14870: inst = 32'hc404ee5;
      14871: inst = 32'h8220000;
      14872: inst = 32'h10408000;
      14873: inst = 32'hc404ee6;
      14874: inst = 32'h8220000;
      14875: inst = 32'h10408000;
      14876: inst = 32'hc404ee7;
      14877: inst = 32'h8220000;
      14878: inst = 32'h10408000;
      14879: inst = 32'hc404ee8;
      14880: inst = 32'h8220000;
      14881: inst = 32'h10408000;
      14882: inst = 32'hc404ee9;
      14883: inst = 32'h8220000;
      14884: inst = 32'h10408000;
      14885: inst = 32'hc404eeb;
      14886: inst = 32'h8220000;
      14887: inst = 32'h10408000;
      14888: inst = 32'hc404eec;
      14889: inst = 32'h8220000;
      14890: inst = 32'h10408000;
      14891: inst = 32'hc404eed;
      14892: inst = 32'h8220000;
      14893: inst = 32'h10408000;
      14894: inst = 32'hc404eee;
      14895: inst = 32'h8220000;
      14896: inst = 32'h10408000;
      14897: inst = 32'hc404eef;
      14898: inst = 32'h8220000;
      14899: inst = 32'h10408000;
      14900: inst = 32'hc404ef0;
      14901: inst = 32'h8220000;
      14902: inst = 32'h10408000;
      14903: inst = 32'hc404ef1;
      14904: inst = 32'h8220000;
      14905: inst = 32'h10408000;
      14906: inst = 32'hc404ef2;
      14907: inst = 32'h8220000;
      14908: inst = 32'h10408000;
      14909: inst = 32'hc404ef3;
      14910: inst = 32'h8220000;
      14911: inst = 32'h10408000;
      14912: inst = 32'hc404f41;
      14913: inst = 32'h8220000;
      14914: inst = 32'h10408000;
      14915: inst = 32'hc404f42;
      14916: inst = 32'h8220000;
      14917: inst = 32'h10408000;
      14918: inst = 32'hc404f43;
      14919: inst = 32'h8220000;
      14920: inst = 32'h10408000;
      14921: inst = 32'hc404f44;
      14922: inst = 32'h8220000;
      14923: inst = 32'h10408000;
      14924: inst = 32'hc404f45;
      14925: inst = 32'h8220000;
      14926: inst = 32'h10408000;
      14927: inst = 32'hc404f46;
      14928: inst = 32'h8220000;
      14929: inst = 32'h10408000;
      14930: inst = 32'hc404f47;
      14931: inst = 32'h8220000;
      14932: inst = 32'h10408000;
      14933: inst = 32'hc404f48;
      14934: inst = 32'h8220000;
      14935: inst = 32'h10408000;
      14936: inst = 32'hc404f49;
      14937: inst = 32'h8220000;
      14938: inst = 32'h10408000;
      14939: inst = 32'hc404f4b;
      14940: inst = 32'h8220000;
      14941: inst = 32'h10408000;
      14942: inst = 32'hc404f4c;
      14943: inst = 32'h8220000;
      14944: inst = 32'h10408000;
      14945: inst = 32'hc404f4d;
      14946: inst = 32'h8220000;
      14947: inst = 32'h10408000;
      14948: inst = 32'hc404f4e;
      14949: inst = 32'h8220000;
      14950: inst = 32'h10408000;
      14951: inst = 32'hc404f4f;
      14952: inst = 32'h8220000;
      14953: inst = 32'h10408000;
      14954: inst = 32'hc404f50;
      14955: inst = 32'h8220000;
      14956: inst = 32'h10408000;
      14957: inst = 32'hc404f51;
      14958: inst = 32'h8220000;
      14959: inst = 32'h10408000;
      14960: inst = 32'hc404f52;
      14961: inst = 32'h8220000;
      14962: inst = 32'h10408000;
      14963: inst = 32'hc404f53;
      14964: inst = 32'h8220000;
      14965: inst = 32'h10408000;
      14966: inst = 32'hc404fa1;
      14967: inst = 32'h8220000;
      14968: inst = 32'h10408000;
      14969: inst = 32'hc404fa2;
      14970: inst = 32'h8220000;
      14971: inst = 32'h10408000;
      14972: inst = 32'hc404fa3;
      14973: inst = 32'h8220000;
      14974: inst = 32'h10408000;
      14975: inst = 32'hc404fa4;
      14976: inst = 32'h8220000;
      14977: inst = 32'h10408000;
      14978: inst = 32'hc404fa5;
      14979: inst = 32'h8220000;
      14980: inst = 32'h10408000;
      14981: inst = 32'hc404fa6;
      14982: inst = 32'h8220000;
      14983: inst = 32'h10408000;
      14984: inst = 32'hc404fa7;
      14985: inst = 32'h8220000;
      14986: inst = 32'h10408000;
      14987: inst = 32'hc404fa9;
      14988: inst = 32'h8220000;
      14989: inst = 32'h10408000;
      14990: inst = 32'hc404fab;
      14991: inst = 32'h8220000;
      14992: inst = 32'h10408000;
      14993: inst = 32'hc404fad;
      14994: inst = 32'h8220000;
      14995: inst = 32'h10408000;
      14996: inst = 32'hc404fae;
      14997: inst = 32'h8220000;
      14998: inst = 32'h10408000;
      14999: inst = 32'hc404faf;
      15000: inst = 32'h8220000;
      15001: inst = 32'h10408000;
      15002: inst = 32'hc404fb0;
      15003: inst = 32'h8220000;
      15004: inst = 32'h10408000;
      15005: inst = 32'hc404fb1;
      15006: inst = 32'h8220000;
      15007: inst = 32'h10408000;
      15008: inst = 32'hc404fb2;
      15009: inst = 32'h8220000;
      15010: inst = 32'h10408000;
      15011: inst = 32'hc404fb3;
      15012: inst = 32'h8220000;
      15013: inst = 32'h10408000;
      15014: inst = 32'hc405001;
      15015: inst = 32'h8220000;
      15016: inst = 32'h10408000;
      15017: inst = 32'hc405002;
      15018: inst = 32'h8220000;
      15019: inst = 32'h10408000;
      15020: inst = 32'hc405003;
      15021: inst = 32'h8220000;
      15022: inst = 32'h10408000;
      15023: inst = 32'hc405004;
      15024: inst = 32'h8220000;
      15025: inst = 32'h10408000;
      15026: inst = 32'hc405005;
      15027: inst = 32'h8220000;
      15028: inst = 32'h10408000;
      15029: inst = 32'hc405006;
      15030: inst = 32'h8220000;
      15031: inst = 32'h10408000;
      15032: inst = 32'hc405007;
      15033: inst = 32'h8220000;
      15034: inst = 32'h10408000;
      15035: inst = 32'hc405009;
      15036: inst = 32'h8220000;
      15037: inst = 32'h10408000;
      15038: inst = 32'hc40500b;
      15039: inst = 32'h8220000;
      15040: inst = 32'h10408000;
      15041: inst = 32'hc40500d;
      15042: inst = 32'h8220000;
      15043: inst = 32'h10408000;
      15044: inst = 32'hc40500e;
      15045: inst = 32'h8220000;
      15046: inst = 32'h10408000;
      15047: inst = 32'hc40500f;
      15048: inst = 32'h8220000;
      15049: inst = 32'h10408000;
      15050: inst = 32'hc405010;
      15051: inst = 32'h8220000;
      15052: inst = 32'h10408000;
      15053: inst = 32'hc405011;
      15054: inst = 32'h8220000;
      15055: inst = 32'h10408000;
      15056: inst = 32'hc405012;
      15057: inst = 32'h8220000;
      15058: inst = 32'h10408000;
      15059: inst = 32'hc405013;
      15060: inst = 32'h8220000;
      15061: inst = 32'h10408000;
      15062: inst = 32'hc405061;
      15063: inst = 32'h8220000;
      15064: inst = 32'h10408000;
      15065: inst = 32'hc405062;
      15066: inst = 32'h8220000;
      15067: inst = 32'h10408000;
      15068: inst = 32'hc405063;
      15069: inst = 32'h8220000;
      15070: inst = 32'h10408000;
      15071: inst = 32'hc405064;
      15072: inst = 32'h8220000;
      15073: inst = 32'h10408000;
      15074: inst = 32'hc405065;
      15075: inst = 32'h8220000;
      15076: inst = 32'h10408000;
      15077: inst = 32'hc405066;
      15078: inst = 32'h8220000;
      15079: inst = 32'h10408000;
      15080: inst = 32'hc405067;
      15081: inst = 32'h8220000;
      15082: inst = 32'h10408000;
      15083: inst = 32'hc405068;
      15084: inst = 32'h8220000;
      15085: inst = 32'h10408000;
      15086: inst = 32'hc405069;
      15087: inst = 32'h8220000;
      15088: inst = 32'h10408000;
      15089: inst = 32'hc40506b;
      15090: inst = 32'h8220000;
      15091: inst = 32'h10408000;
      15092: inst = 32'hc40506c;
      15093: inst = 32'h8220000;
      15094: inst = 32'h10408000;
      15095: inst = 32'hc40506d;
      15096: inst = 32'h8220000;
      15097: inst = 32'h10408000;
      15098: inst = 32'hc40506e;
      15099: inst = 32'h8220000;
      15100: inst = 32'h10408000;
      15101: inst = 32'hc40506f;
      15102: inst = 32'h8220000;
      15103: inst = 32'h10408000;
      15104: inst = 32'hc405070;
      15105: inst = 32'h8220000;
      15106: inst = 32'h10408000;
      15107: inst = 32'hc405071;
      15108: inst = 32'h8220000;
      15109: inst = 32'h10408000;
      15110: inst = 32'hc405072;
      15111: inst = 32'h8220000;
      15112: inst = 32'h10408000;
      15113: inst = 32'hc405073;
      15114: inst = 32'h8220000;
      15115: inst = 32'h10408000;
      15116: inst = 32'hc4050c1;
      15117: inst = 32'h8220000;
      15118: inst = 32'h10408000;
      15119: inst = 32'hc4050c2;
      15120: inst = 32'h8220000;
      15121: inst = 32'h10408000;
      15122: inst = 32'hc4050c3;
      15123: inst = 32'h8220000;
      15124: inst = 32'h10408000;
      15125: inst = 32'hc4050c4;
      15126: inst = 32'h8220000;
      15127: inst = 32'h10408000;
      15128: inst = 32'hc4050c5;
      15129: inst = 32'h8220000;
      15130: inst = 32'h10408000;
      15131: inst = 32'hc4050c6;
      15132: inst = 32'h8220000;
      15133: inst = 32'h10408000;
      15134: inst = 32'hc4050c7;
      15135: inst = 32'h8220000;
      15136: inst = 32'h10408000;
      15137: inst = 32'hc4050c8;
      15138: inst = 32'h8220000;
      15139: inst = 32'h10408000;
      15140: inst = 32'hc4050c9;
      15141: inst = 32'h8220000;
      15142: inst = 32'h10408000;
      15143: inst = 32'hc4050cb;
      15144: inst = 32'h8220000;
      15145: inst = 32'h10408000;
      15146: inst = 32'hc4050cc;
      15147: inst = 32'h8220000;
      15148: inst = 32'h10408000;
      15149: inst = 32'hc4050cd;
      15150: inst = 32'h8220000;
      15151: inst = 32'h10408000;
      15152: inst = 32'hc4050ce;
      15153: inst = 32'h8220000;
      15154: inst = 32'h10408000;
      15155: inst = 32'hc4050cf;
      15156: inst = 32'h8220000;
      15157: inst = 32'h10408000;
      15158: inst = 32'hc4050d0;
      15159: inst = 32'h8220000;
      15160: inst = 32'h10408000;
      15161: inst = 32'hc4050d1;
      15162: inst = 32'h8220000;
      15163: inst = 32'h10408000;
      15164: inst = 32'hc4050d2;
      15165: inst = 32'h8220000;
      15166: inst = 32'h10408000;
      15167: inst = 32'hc4050d3;
      15168: inst = 32'h8220000;
      15169: inst = 32'h10408000;
      15170: inst = 32'hc405121;
      15171: inst = 32'h8220000;
      15172: inst = 32'h10408000;
      15173: inst = 32'hc405122;
      15174: inst = 32'h8220000;
      15175: inst = 32'h10408000;
      15176: inst = 32'hc405123;
      15177: inst = 32'h8220000;
      15178: inst = 32'h10408000;
      15179: inst = 32'hc405124;
      15180: inst = 32'h8220000;
      15181: inst = 32'h10408000;
      15182: inst = 32'hc405125;
      15183: inst = 32'h8220000;
      15184: inst = 32'h10408000;
      15185: inst = 32'hc405126;
      15186: inst = 32'h8220000;
      15187: inst = 32'h10408000;
      15188: inst = 32'hc405127;
      15189: inst = 32'h8220000;
      15190: inst = 32'h10408000;
      15191: inst = 32'hc405128;
      15192: inst = 32'h8220000;
      15193: inst = 32'h10408000;
      15194: inst = 32'hc405129;
      15195: inst = 32'h8220000;
      15196: inst = 32'h10408000;
      15197: inst = 32'hc40512b;
      15198: inst = 32'h8220000;
      15199: inst = 32'h10408000;
      15200: inst = 32'hc40512c;
      15201: inst = 32'h8220000;
      15202: inst = 32'h10408000;
      15203: inst = 32'hc40512d;
      15204: inst = 32'h8220000;
      15205: inst = 32'h10408000;
      15206: inst = 32'hc40512e;
      15207: inst = 32'h8220000;
      15208: inst = 32'h10408000;
      15209: inst = 32'hc40512f;
      15210: inst = 32'h8220000;
      15211: inst = 32'h10408000;
      15212: inst = 32'hc405130;
      15213: inst = 32'h8220000;
      15214: inst = 32'h10408000;
      15215: inst = 32'hc405131;
      15216: inst = 32'h8220000;
      15217: inst = 32'h10408000;
      15218: inst = 32'hc405132;
      15219: inst = 32'h8220000;
      15220: inst = 32'h10408000;
      15221: inst = 32'hc405133;
      15222: inst = 32'h8220000;
      15223: inst = 32'h10408000;
      15224: inst = 32'hc405181;
      15225: inst = 32'h8220000;
      15226: inst = 32'h10408000;
      15227: inst = 32'hc405182;
      15228: inst = 32'h8220000;
      15229: inst = 32'h10408000;
      15230: inst = 32'hc405183;
      15231: inst = 32'h8220000;
      15232: inst = 32'h10408000;
      15233: inst = 32'hc405184;
      15234: inst = 32'h8220000;
      15235: inst = 32'h10408000;
      15236: inst = 32'hc405185;
      15237: inst = 32'h8220000;
      15238: inst = 32'h10408000;
      15239: inst = 32'hc405186;
      15240: inst = 32'h8220000;
      15241: inst = 32'h10408000;
      15242: inst = 32'hc405187;
      15243: inst = 32'h8220000;
      15244: inst = 32'h10408000;
      15245: inst = 32'hc405188;
      15246: inst = 32'h8220000;
      15247: inst = 32'h10408000;
      15248: inst = 32'hc405189;
      15249: inst = 32'h8220000;
      15250: inst = 32'h10408000;
      15251: inst = 32'hc40518b;
      15252: inst = 32'h8220000;
      15253: inst = 32'h10408000;
      15254: inst = 32'hc40518c;
      15255: inst = 32'h8220000;
      15256: inst = 32'h10408000;
      15257: inst = 32'hc40518d;
      15258: inst = 32'h8220000;
      15259: inst = 32'h10408000;
      15260: inst = 32'hc40518e;
      15261: inst = 32'h8220000;
      15262: inst = 32'h10408000;
      15263: inst = 32'hc40518f;
      15264: inst = 32'h8220000;
      15265: inst = 32'h10408000;
      15266: inst = 32'hc405190;
      15267: inst = 32'h8220000;
      15268: inst = 32'h10408000;
      15269: inst = 32'hc405191;
      15270: inst = 32'h8220000;
      15271: inst = 32'h10408000;
      15272: inst = 32'hc405192;
      15273: inst = 32'h8220000;
      15274: inst = 32'h10408000;
      15275: inst = 32'hc405193;
      15276: inst = 32'h8220000;
      15277: inst = 32'h10408000;
      15278: inst = 32'hc4051e1;
      15279: inst = 32'h8220000;
      15280: inst = 32'h10408000;
      15281: inst = 32'hc4051e2;
      15282: inst = 32'h8220000;
      15283: inst = 32'h10408000;
      15284: inst = 32'hc4051e3;
      15285: inst = 32'h8220000;
      15286: inst = 32'h10408000;
      15287: inst = 32'hc4051e4;
      15288: inst = 32'h8220000;
      15289: inst = 32'h10408000;
      15290: inst = 32'hc4051e5;
      15291: inst = 32'h8220000;
      15292: inst = 32'h10408000;
      15293: inst = 32'hc4051e6;
      15294: inst = 32'h8220000;
      15295: inst = 32'h10408000;
      15296: inst = 32'hc4051e7;
      15297: inst = 32'h8220000;
      15298: inst = 32'h10408000;
      15299: inst = 32'hc4051e8;
      15300: inst = 32'h8220000;
      15301: inst = 32'h10408000;
      15302: inst = 32'hc4051e9;
      15303: inst = 32'h8220000;
      15304: inst = 32'h10408000;
      15305: inst = 32'hc4051eb;
      15306: inst = 32'h8220000;
      15307: inst = 32'h10408000;
      15308: inst = 32'hc4051ec;
      15309: inst = 32'h8220000;
      15310: inst = 32'h10408000;
      15311: inst = 32'hc4051ed;
      15312: inst = 32'h8220000;
      15313: inst = 32'h10408000;
      15314: inst = 32'hc4051ee;
      15315: inst = 32'h8220000;
      15316: inst = 32'h10408000;
      15317: inst = 32'hc4051ef;
      15318: inst = 32'h8220000;
      15319: inst = 32'h10408000;
      15320: inst = 32'hc4051f0;
      15321: inst = 32'h8220000;
      15322: inst = 32'h10408000;
      15323: inst = 32'hc4051f1;
      15324: inst = 32'h8220000;
      15325: inst = 32'h10408000;
      15326: inst = 32'hc4051f2;
      15327: inst = 32'h8220000;
      15328: inst = 32'h10408000;
      15329: inst = 32'hc4051f3;
      15330: inst = 32'h8220000;
      15331: inst = 32'h10408000;
      15332: inst = 32'hc405241;
      15333: inst = 32'h8220000;
      15334: inst = 32'h10408000;
      15335: inst = 32'hc405242;
      15336: inst = 32'h8220000;
      15337: inst = 32'h10408000;
      15338: inst = 32'hc405243;
      15339: inst = 32'h8220000;
      15340: inst = 32'h10408000;
      15341: inst = 32'hc405244;
      15342: inst = 32'h8220000;
      15343: inst = 32'h10408000;
      15344: inst = 32'hc405245;
      15345: inst = 32'h8220000;
      15346: inst = 32'h10408000;
      15347: inst = 32'hc405246;
      15348: inst = 32'h8220000;
      15349: inst = 32'h10408000;
      15350: inst = 32'hc405247;
      15351: inst = 32'h8220000;
      15352: inst = 32'h10408000;
      15353: inst = 32'hc405248;
      15354: inst = 32'h8220000;
      15355: inst = 32'h10408000;
      15356: inst = 32'hc405249;
      15357: inst = 32'h8220000;
      15358: inst = 32'h10408000;
      15359: inst = 32'hc40524b;
      15360: inst = 32'h8220000;
      15361: inst = 32'h10408000;
      15362: inst = 32'hc40524c;
      15363: inst = 32'h8220000;
      15364: inst = 32'h10408000;
      15365: inst = 32'hc40524d;
      15366: inst = 32'h8220000;
      15367: inst = 32'h10408000;
      15368: inst = 32'hc40524e;
      15369: inst = 32'h8220000;
      15370: inst = 32'h10408000;
      15371: inst = 32'hc40524f;
      15372: inst = 32'h8220000;
      15373: inst = 32'h10408000;
      15374: inst = 32'hc405250;
      15375: inst = 32'h8220000;
      15376: inst = 32'h10408000;
      15377: inst = 32'hc405251;
      15378: inst = 32'h8220000;
      15379: inst = 32'h10408000;
      15380: inst = 32'hc405252;
      15381: inst = 32'h8220000;
      15382: inst = 32'h10408000;
      15383: inst = 32'hc405253;
      15384: inst = 32'h8220000;
      15385: inst = 32'hc20bd73;
      15386: inst = 32'h10408000;
      15387: inst = 32'hc404e9f;
      15388: inst = 32'h8220000;
      15389: inst = 32'h10408000;
      15390: inst = 32'hc404ec0;
      15391: inst = 32'h8220000;
      15392: inst = 32'hc205aed;
      15393: inst = 32'h10408000;
      15394: inst = 32'hc404ea0;
      15395: inst = 32'h8220000;
      15396: inst = 32'h10408000;
      15397: inst = 32'hc404ea1;
      15398: inst = 32'h8220000;
      15399: inst = 32'h10408000;
      15400: inst = 32'hc404ea2;
      15401: inst = 32'h8220000;
      15402: inst = 32'h10408000;
      15403: inst = 32'hc404ea3;
      15404: inst = 32'h8220000;
      15405: inst = 32'h10408000;
      15406: inst = 32'hc404ea4;
      15407: inst = 32'h8220000;
      15408: inst = 32'h10408000;
      15409: inst = 32'hc404ebb;
      15410: inst = 32'h8220000;
      15411: inst = 32'h10408000;
      15412: inst = 32'hc404ebc;
      15413: inst = 32'h8220000;
      15414: inst = 32'h10408000;
      15415: inst = 32'hc404ebd;
      15416: inst = 32'h8220000;
      15417: inst = 32'h10408000;
      15418: inst = 32'hc404ebe;
      15419: inst = 32'h8220000;
      15420: inst = 32'h10408000;
      15421: inst = 32'hc404ebf;
      15422: inst = 32'h8220000;
      15423: inst = 32'h10408000;
      15424: inst = 32'hc404f00;
      15425: inst = 32'h8220000;
      15426: inst = 32'h10408000;
      15427: inst = 32'hc404f01;
      15428: inst = 32'h8220000;
      15429: inst = 32'h10408000;
      15430: inst = 32'hc404f02;
      15431: inst = 32'h8220000;
      15432: inst = 32'h10408000;
      15433: inst = 32'hc404f03;
      15434: inst = 32'h8220000;
      15435: inst = 32'h10408000;
      15436: inst = 32'hc404f04;
      15437: inst = 32'h8220000;
      15438: inst = 32'h10408000;
      15439: inst = 32'hc404f05;
      15440: inst = 32'h8220000;
      15441: inst = 32'h10408000;
      15442: inst = 32'hc404f1a;
      15443: inst = 32'h8220000;
      15444: inst = 32'h10408000;
      15445: inst = 32'hc404f1b;
      15446: inst = 32'h8220000;
      15447: inst = 32'h10408000;
      15448: inst = 32'hc404f1c;
      15449: inst = 32'h8220000;
      15450: inst = 32'h10408000;
      15451: inst = 32'hc404f1d;
      15452: inst = 32'h8220000;
      15453: inst = 32'h10408000;
      15454: inst = 32'hc404f1e;
      15455: inst = 32'h8220000;
      15456: inst = 32'h10408000;
      15457: inst = 32'hc404f1f;
      15458: inst = 32'h8220000;
      15459: inst = 32'h10408000;
      15460: inst = 32'hc404f60;
      15461: inst = 32'h8220000;
      15462: inst = 32'h10408000;
      15463: inst = 32'hc404f61;
      15464: inst = 32'h8220000;
      15465: inst = 32'h10408000;
      15466: inst = 32'hc404f62;
      15467: inst = 32'h8220000;
      15468: inst = 32'h10408000;
      15469: inst = 32'hc404f63;
      15470: inst = 32'h8220000;
      15471: inst = 32'h10408000;
      15472: inst = 32'hc404f64;
      15473: inst = 32'h8220000;
      15474: inst = 32'h10408000;
      15475: inst = 32'hc404f65;
      15476: inst = 32'h8220000;
      15477: inst = 32'h10408000;
      15478: inst = 32'hc404f66;
      15479: inst = 32'h8220000;
      15480: inst = 32'h10408000;
      15481: inst = 32'hc404f67;
      15482: inst = 32'h8220000;
      15483: inst = 32'h10408000;
      15484: inst = 32'hc404f78;
      15485: inst = 32'h8220000;
      15486: inst = 32'h10408000;
      15487: inst = 32'hc404f79;
      15488: inst = 32'h8220000;
      15489: inst = 32'h10408000;
      15490: inst = 32'hc404f7a;
      15491: inst = 32'h8220000;
      15492: inst = 32'h10408000;
      15493: inst = 32'hc404f7b;
      15494: inst = 32'h8220000;
      15495: inst = 32'h10408000;
      15496: inst = 32'hc404f7c;
      15497: inst = 32'h8220000;
      15498: inst = 32'h10408000;
      15499: inst = 32'hc404f7d;
      15500: inst = 32'h8220000;
      15501: inst = 32'h10408000;
      15502: inst = 32'hc404f7e;
      15503: inst = 32'h8220000;
      15504: inst = 32'h10408000;
      15505: inst = 32'hc404f7f;
      15506: inst = 32'h8220000;
      15507: inst = 32'h10408000;
      15508: inst = 32'hc404fc0;
      15509: inst = 32'h8220000;
      15510: inst = 32'h10408000;
      15511: inst = 32'hc404fc1;
      15512: inst = 32'h8220000;
      15513: inst = 32'h10408000;
      15514: inst = 32'hc404fc2;
      15515: inst = 32'h8220000;
      15516: inst = 32'h10408000;
      15517: inst = 32'hc404fc3;
      15518: inst = 32'h8220000;
      15519: inst = 32'h10408000;
      15520: inst = 32'hc404fc4;
      15521: inst = 32'h8220000;
      15522: inst = 32'h10408000;
      15523: inst = 32'hc404fc6;
      15524: inst = 32'h8220000;
      15525: inst = 32'h10408000;
      15526: inst = 32'hc404fc7;
      15527: inst = 32'h8220000;
      15528: inst = 32'h10408000;
      15529: inst = 32'hc404fd8;
      15530: inst = 32'h8220000;
      15531: inst = 32'h10408000;
      15532: inst = 32'hc404fd9;
      15533: inst = 32'h8220000;
      15534: inst = 32'h10408000;
      15535: inst = 32'hc404fdb;
      15536: inst = 32'h8220000;
      15537: inst = 32'h10408000;
      15538: inst = 32'hc404fdc;
      15539: inst = 32'h8220000;
      15540: inst = 32'h10408000;
      15541: inst = 32'hc404fdd;
      15542: inst = 32'h8220000;
      15543: inst = 32'h10408000;
      15544: inst = 32'hc404fde;
      15545: inst = 32'h8220000;
      15546: inst = 32'h10408000;
      15547: inst = 32'hc404fdf;
      15548: inst = 32'h8220000;
      15549: inst = 32'h10408000;
      15550: inst = 32'hc405020;
      15551: inst = 32'h8220000;
      15552: inst = 32'h10408000;
      15553: inst = 32'hc405021;
      15554: inst = 32'h8220000;
      15555: inst = 32'h10408000;
      15556: inst = 32'hc405022;
      15557: inst = 32'h8220000;
      15558: inst = 32'h10408000;
      15559: inst = 32'hc405023;
      15560: inst = 32'h8220000;
      15561: inst = 32'h10408000;
      15562: inst = 32'hc405026;
      15563: inst = 32'h8220000;
      15564: inst = 32'h10408000;
      15565: inst = 32'hc405027;
      15566: inst = 32'h8220000;
      15567: inst = 32'h10408000;
      15568: inst = 32'hc405038;
      15569: inst = 32'h8220000;
      15570: inst = 32'h10408000;
      15571: inst = 32'hc405039;
      15572: inst = 32'h8220000;
      15573: inst = 32'h10408000;
      15574: inst = 32'hc40503c;
      15575: inst = 32'h8220000;
      15576: inst = 32'h10408000;
      15577: inst = 32'hc40503d;
      15578: inst = 32'h8220000;
      15579: inst = 32'h10408000;
      15580: inst = 32'hc40503e;
      15581: inst = 32'h8220000;
      15582: inst = 32'h10408000;
      15583: inst = 32'hc40503f;
      15584: inst = 32'h8220000;
      15585: inst = 32'h10408000;
      15586: inst = 32'hc40507f;
      15587: inst = 32'h8220000;
      15588: inst = 32'h10408000;
      15589: inst = 32'hc405080;
      15590: inst = 32'h8220000;
      15591: inst = 32'h10408000;
      15592: inst = 32'hc405081;
      15593: inst = 32'h8220000;
      15594: inst = 32'h10408000;
      15595: inst = 32'hc405082;
      15596: inst = 32'h8220000;
      15597: inst = 32'h10408000;
      15598: inst = 32'hc405086;
      15599: inst = 32'h8220000;
      15600: inst = 32'h10408000;
      15601: inst = 32'hc405087;
      15602: inst = 32'h8220000;
      15603: inst = 32'h10408000;
      15604: inst = 32'hc405098;
      15605: inst = 32'h8220000;
      15606: inst = 32'h10408000;
      15607: inst = 32'hc405099;
      15608: inst = 32'h8220000;
      15609: inst = 32'h10408000;
      15610: inst = 32'hc40509d;
      15611: inst = 32'h8220000;
      15612: inst = 32'h10408000;
      15613: inst = 32'hc40509e;
      15614: inst = 32'h8220000;
      15615: inst = 32'h10408000;
      15616: inst = 32'hc40509f;
      15617: inst = 32'h8220000;
      15618: inst = 32'h10408000;
      15619: inst = 32'hc4050a0;
      15620: inst = 32'h8220000;
      15621: inst = 32'h10408000;
      15622: inst = 32'hc4050df;
      15623: inst = 32'h8220000;
      15624: inst = 32'h10408000;
      15625: inst = 32'hc4050e0;
      15626: inst = 32'h8220000;
      15627: inst = 32'h10408000;
      15628: inst = 32'hc4050e1;
      15629: inst = 32'h8220000;
      15630: inst = 32'h10408000;
      15631: inst = 32'hc4050e2;
      15632: inst = 32'h8220000;
      15633: inst = 32'h10408000;
      15634: inst = 32'hc4050e6;
      15635: inst = 32'h8220000;
      15636: inst = 32'h10408000;
      15637: inst = 32'hc4050e7;
      15638: inst = 32'h8220000;
      15639: inst = 32'h10408000;
      15640: inst = 32'hc4050f8;
      15641: inst = 32'h8220000;
      15642: inst = 32'h10408000;
      15643: inst = 32'hc4050f9;
      15644: inst = 32'h8220000;
      15645: inst = 32'h10408000;
      15646: inst = 32'hc4050fd;
      15647: inst = 32'h8220000;
      15648: inst = 32'h10408000;
      15649: inst = 32'hc4050fe;
      15650: inst = 32'h8220000;
      15651: inst = 32'h10408000;
      15652: inst = 32'hc4050ff;
      15653: inst = 32'h8220000;
      15654: inst = 32'h10408000;
      15655: inst = 32'hc405100;
      15656: inst = 32'h8220000;
      15657: inst = 32'h10408000;
      15658: inst = 32'hc40513f;
      15659: inst = 32'h8220000;
      15660: inst = 32'h10408000;
      15661: inst = 32'hc405140;
      15662: inst = 32'h8220000;
      15663: inst = 32'h10408000;
      15664: inst = 32'hc405141;
      15665: inst = 32'h8220000;
      15666: inst = 32'h10408000;
      15667: inst = 32'hc405146;
      15668: inst = 32'h8220000;
      15669: inst = 32'h10408000;
      15670: inst = 32'hc405147;
      15671: inst = 32'h8220000;
      15672: inst = 32'h10408000;
      15673: inst = 32'hc405158;
      15674: inst = 32'h8220000;
      15675: inst = 32'h10408000;
      15676: inst = 32'hc405159;
      15677: inst = 32'h8220000;
      15678: inst = 32'h10408000;
      15679: inst = 32'hc40515e;
      15680: inst = 32'h8220000;
      15681: inst = 32'h10408000;
      15682: inst = 32'hc40515f;
      15683: inst = 32'h8220000;
      15684: inst = 32'h10408000;
      15685: inst = 32'hc405160;
      15686: inst = 32'h8220000;
      15687: inst = 32'h10408000;
      15688: inst = 32'hc40519f;
      15689: inst = 32'h8220000;
      15690: inst = 32'h10408000;
      15691: inst = 32'hc4051a0;
      15692: inst = 32'h8220000;
      15693: inst = 32'h10408000;
      15694: inst = 32'hc4051a6;
      15695: inst = 32'h8220000;
      15696: inst = 32'h10408000;
      15697: inst = 32'hc4051a7;
      15698: inst = 32'h8220000;
      15699: inst = 32'h10408000;
      15700: inst = 32'hc4051b8;
      15701: inst = 32'h8220000;
      15702: inst = 32'h10408000;
      15703: inst = 32'hc4051b9;
      15704: inst = 32'h8220000;
      15705: inst = 32'h10408000;
      15706: inst = 32'hc4051bf;
      15707: inst = 32'h8220000;
      15708: inst = 32'h10408000;
      15709: inst = 32'hc4051c0;
      15710: inst = 32'h8220000;
      15711: inst = 32'h10408000;
      15712: inst = 32'hc4051ff;
      15713: inst = 32'h8220000;
      15714: inst = 32'h10408000;
      15715: inst = 32'hc405200;
      15716: inst = 32'h8220000;
      15717: inst = 32'h10408000;
      15718: inst = 32'hc405206;
      15719: inst = 32'h8220000;
      15720: inst = 32'h10408000;
      15721: inst = 32'hc405207;
      15722: inst = 32'h8220000;
      15723: inst = 32'h10408000;
      15724: inst = 32'hc405218;
      15725: inst = 32'h8220000;
      15726: inst = 32'h10408000;
      15727: inst = 32'hc405219;
      15728: inst = 32'h8220000;
      15729: inst = 32'h10408000;
      15730: inst = 32'hc40521f;
      15731: inst = 32'h8220000;
      15732: inst = 32'h10408000;
      15733: inst = 32'hc405220;
      15734: inst = 32'h8220000;
      15735: inst = 32'h10408000;
      15736: inst = 32'hc40525f;
      15737: inst = 32'h8220000;
      15738: inst = 32'h10408000;
      15739: inst = 32'hc405260;
      15740: inst = 32'h8220000;
      15741: inst = 32'h10408000;
      15742: inst = 32'hc405266;
      15743: inst = 32'h8220000;
      15744: inst = 32'h10408000;
      15745: inst = 32'hc405267;
      15746: inst = 32'h8220000;
      15747: inst = 32'h10408000;
      15748: inst = 32'hc405278;
      15749: inst = 32'h8220000;
      15750: inst = 32'h10408000;
      15751: inst = 32'hc405279;
      15752: inst = 32'h8220000;
      15753: inst = 32'h10408000;
      15754: inst = 32'hc40527f;
      15755: inst = 32'h8220000;
      15756: inst = 32'h10408000;
      15757: inst = 32'hc405280;
      15758: inst = 32'h8220000;
      15759: inst = 32'h10408000;
      15760: inst = 32'hc4052bf;
      15761: inst = 32'h8220000;
      15762: inst = 32'h10408000;
      15763: inst = 32'hc4052c0;
      15764: inst = 32'h8220000;
      15765: inst = 32'h10408000;
      15766: inst = 32'hc4052c6;
      15767: inst = 32'h8220000;
      15768: inst = 32'h10408000;
      15769: inst = 32'hc4052c7;
      15770: inst = 32'h8220000;
      15771: inst = 32'h10408000;
      15772: inst = 32'hc4052d8;
      15773: inst = 32'h8220000;
      15774: inst = 32'h10408000;
      15775: inst = 32'hc4052d9;
      15776: inst = 32'h8220000;
      15777: inst = 32'h10408000;
      15778: inst = 32'hc4052df;
      15779: inst = 32'h8220000;
      15780: inst = 32'h10408000;
      15781: inst = 32'hc4052e0;
      15782: inst = 32'h8220000;
      15783: inst = 32'hc207bae;
      15784: inst = 32'h10408000;
      15785: inst = 32'hc404ea5;
      15786: inst = 32'h8220000;
      15787: inst = 32'h10408000;
      15788: inst = 32'hc404eba;
      15789: inst = 32'h8220000;
      15790: inst = 32'hc20c5b4;
      15791: inst = 32'h10408000;
      15792: inst = 32'hc404ea6;
      15793: inst = 32'h8220000;
      15794: inst = 32'h10408000;
      15795: inst = 32'hc404eb9;
      15796: inst = 32'h8220000;
      15797: inst = 32'hc20d5f4;
      15798: inst = 32'h10408000;
      15799: inst = 32'hc404ea7;
      15800: inst = 32'h8220000;
      15801: inst = 32'h10408000;
      15802: inst = 32'hc404eb8;
      15803: inst = 32'h8220000;
      15804: inst = 32'hc20a4b1;
      15805: inst = 32'h10408000;
      15806: inst = 32'hc404eff;
      15807: inst = 32'h8220000;
      15808: inst = 32'h10408000;
      15809: inst = 32'hc404f20;
      15810: inst = 32'h8220000;
      15811: inst = 32'h10408000;
      15812: inst = 32'hc404fbf;
      15813: inst = 32'h8220000;
      15814: inst = 32'h10408000;
      15815: inst = 32'hc404fe0;
      15816: inst = 32'h8220000;
      15817: inst = 32'hc2062ed;
      15818: inst = 32'h10408000;
      15819: inst = 32'hc404f06;
      15820: inst = 32'h8220000;
      15821: inst = 32'h10408000;
      15822: inst = 32'hc404f19;
      15823: inst = 32'h8220000;
      15824: inst = 32'hc209450;
      15825: inst = 32'h10408000;
      15826: inst = 32'hc404f07;
      15827: inst = 32'h8220000;
      15828: inst = 32'h10408000;
      15829: inst = 32'hc404f18;
      15830: inst = 32'h8220000;
      15831: inst = 32'h10408000;
      15832: inst = 32'hc405209;
      15833: inst = 32'h8220000;
      15834: inst = 32'h10408000;
      15835: inst = 32'hc405216;
      15836: inst = 32'h8220000;
      15837: inst = 32'hc20a4d1;
      15838: inst = 32'h10408000;
      15839: inst = 32'hc404f5f;
      15840: inst = 32'h8220000;
      15841: inst = 32'h10408000;
      15842: inst = 32'hc404f80;
      15843: inst = 32'h8220000;
      15844: inst = 32'hc204a49;
      15845: inst = 32'h10408000;
      15846: inst = 32'hc404fa8;
      15847: inst = 32'h8220000;
      15848: inst = 32'h10408000;
      15849: inst = 32'hc404fac;
      15850: inst = 32'h8220000;
      15851: inst = 32'h10408000;
      15852: inst = 32'hc405008;
      15853: inst = 32'h8220000;
      15854: inst = 32'h10408000;
      15855: inst = 32'hc40500c;
      15856: inst = 32'h8220000;
      15857: inst = 32'hc205acb;
      15858: inst = 32'h10408000;
      15859: inst = 32'hc404fc5;
      15860: inst = 32'h8220000;
      15861: inst = 32'h10408000;
      15862: inst = 32'hc404fda;
      15863: inst = 32'h8220000;
      15864: inst = 32'h10408000;
      15865: inst = 32'hc405336;
      15866: inst = 32'h8220000;
      15867: inst = 32'h10408000;
      15868: inst = 32'hc405380;
      15869: inst = 32'h8220000;
      15870: inst = 32'h10408000;
      15871: inst = 32'hc40539f;
      15872: inst = 32'h8220000;
      15873: inst = 32'h10408000;
      15874: inst = 32'hc4053dd;
      15875: inst = 32'h8220000;
      15876: inst = 32'h10408000;
      15877: inst = 32'hc405402;
      15878: inst = 32'h8220000;
      15879: inst = 32'hc20630d;
      15880: inst = 32'h10408000;
      15881: inst = 32'hc40501f;
      15882: inst = 32'h8220000;
      15883: inst = 32'h10408000;
      15884: inst = 32'hc405040;
      15885: inst = 32'h8220000;
      15886: inst = 32'hc205aec;
      15887: inst = 32'h10408000;
      15888: inst = 32'hc405024;
      15889: inst = 32'h8220000;
      15890: inst = 32'h10408000;
      15891: inst = 32'hc40503b;
      15892: inst = 32'h8220000;
      15893: inst = 32'h10408000;
      15894: inst = 32'hc405083;
      15895: inst = 32'h8220000;
      15896: inst = 32'h10408000;
      15897: inst = 32'hc40509c;
      15898: inst = 32'h8220000;
      15899: inst = 32'h10408000;
      15900: inst = 32'hc4051a1;
      15901: inst = 32'h8220000;
      15902: inst = 32'h10408000;
      15903: inst = 32'hc4051be;
      15904: inst = 32'h8220000;
      15905: inst = 32'h10408000;
      15906: inst = 32'hc405329;
      15907: inst = 32'h8220000;
      15908: inst = 32'h10408000;
      15909: inst = 32'hc405568;
      15910: inst = 32'h8220000;
      15911: inst = 32'h10408000;
      15912: inst = 32'hc405577;
      15913: inst = 32'h8220000;
      15914: inst = 32'h10408000;
      15915: inst = 32'hc4057a7;
      15916: inst = 32'h8220000;
      15917: inst = 32'h10408000;
      15918: inst = 32'hc4057b8;
      15919: inst = 32'h8220000;
      15920: inst = 32'hc205269;
      15921: inst = 32'h10408000;
      15922: inst = 32'hc405025;
      15923: inst = 32'h8220000;
      15924: inst = 32'h10408000;
      15925: inst = 32'hc40503a;
      15926: inst = 32'h8220000;
      15927: inst = 32'h10408000;
      15928: inst = 32'hc40537e;
      15929: inst = 32'h8220000;
      15930: inst = 32'h10408000;
      15931: inst = 32'hc4053a1;
      15932: inst = 32'h8220000;
      15933: inst = 32'h10408000;
      15934: inst = 32'hc40549c;
      15935: inst = 32'h8220000;
      15936: inst = 32'h10408000;
      15937: inst = 32'hc4054c3;
      15938: inst = 32'h8220000;
      15939: inst = 32'hc20528a;
      15940: inst = 32'h10408000;
      15941: inst = 32'hc405084;
      15942: inst = 32'h8220000;
      15943: inst = 32'h10408000;
      15944: inst = 32'hc40509b;
      15945: inst = 32'h8220000;
      15946: inst = 32'h10408000;
      15947: inst = 32'hc4050e3;
      15948: inst = 32'h8220000;
      15949: inst = 32'h10408000;
      15950: inst = 32'hc4050fc;
      15951: inst = 32'h8220000;
      15952: inst = 32'h10408000;
      15953: inst = 32'hc4052c5;
      15954: inst = 32'h8220000;
      15955: inst = 32'h10408000;
      15956: inst = 32'hc4052da;
      15957: inst = 32'h8220000;
      15958: inst = 32'h10408000;
      15959: inst = 32'hc4053e9;
      15960: inst = 32'h8220000;
      15961: inst = 32'h10408000;
      15962: inst = 32'hc4053f6;
      15963: inst = 32'h8220000;
      15964: inst = 32'h10408000;
      15965: inst = 32'hc405449;
      15966: inst = 32'h8220000;
      15967: inst = 32'h10408000;
      15968: inst = 32'hc405456;
      15969: inst = 32'h8220000;
      15970: inst = 32'h10408000;
      15971: inst = 32'hc4054a9;
      15972: inst = 32'h8220000;
      15973: inst = 32'h10408000;
      15974: inst = 32'hc4054b6;
      15975: inst = 32'h8220000;
      15976: inst = 32'h10408000;
      15977: inst = 32'hc405509;
      15978: inst = 32'h8220000;
      15979: inst = 32'h10408000;
      15980: inst = 32'hc405516;
      15981: inst = 32'h8220000;
      15982: inst = 32'h10408000;
      15983: inst = 32'hc40555e;
      15984: inst = 32'h8220000;
      15985: inst = 32'h10408000;
      15986: inst = 32'hc405569;
      15987: inst = 32'h8220000;
      15988: inst = 32'h10408000;
      15989: inst = 32'hc405576;
      15990: inst = 32'h8220000;
      15991: inst = 32'h10408000;
      15992: inst = 32'hc405581;
      15993: inst = 32'h8220000;
      15994: inst = 32'h10408000;
      15995: inst = 32'hc4055c9;
      15996: inst = 32'h8220000;
      15997: inst = 32'h10408000;
      15998: inst = 32'hc4055d6;
      15999: inst = 32'h8220000;
      16000: inst = 32'h10408000;
      16001: inst = 32'hc405628;
      16002: inst = 32'h8220000;
      16003: inst = 32'h10408000;
      16004: inst = 32'hc405629;
      16005: inst = 32'h8220000;
      16006: inst = 32'h10408000;
      16007: inst = 32'hc405636;
      16008: inst = 32'h8220000;
      16009: inst = 32'h10408000;
      16010: inst = 32'hc405637;
      16011: inst = 32'h8220000;
      16012: inst = 32'h10408000;
      16013: inst = 32'hc40567d;
      16014: inst = 32'h8220000;
      16015: inst = 32'h10408000;
      16016: inst = 32'hc405688;
      16017: inst = 32'h8220000;
      16018: inst = 32'h10408000;
      16019: inst = 32'hc405689;
      16020: inst = 32'h8220000;
      16021: inst = 32'h10408000;
      16022: inst = 32'hc405696;
      16023: inst = 32'h8220000;
      16024: inst = 32'h10408000;
      16025: inst = 32'hc405697;
      16026: inst = 32'h8220000;
      16027: inst = 32'h10408000;
      16028: inst = 32'hc4056a2;
      16029: inst = 32'h8220000;
      16030: inst = 32'h10408000;
      16031: inst = 32'hc4056e8;
      16032: inst = 32'h8220000;
      16033: inst = 32'h10408000;
      16034: inst = 32'hc4056e9;
      16035: inst = 32'h8220000;
      16036: inst = 32'h10408000;
      16037: inst = 32'hc4056f6;
      16038: inst = 32'h8220000;
      16039: inst = 32'h10408000;
      16040: inst = 32'hc4056f7;
      16041: inst = 32'h8220000;
      16042: inst = 32'h10408000;
      16043: inst = 32'hc405748;
      16044: inst = 32'h8220000;
      16045: inst = 32'h10408000;
      16046: inst = 32'hc405749;
      16047: inst = 32'h8220000;
      16048: inst = 32'h10408000;
      16049: inst = 32'hc405756;
      16050: inst = 32'h8220000;
      16051: inst = 32'h10408000;
      16052: inst = 32'hc405757;
      16053: inst = 32'h8220000;
      16054: inst = 32'h10408000;
      16055: inst = 32'hc4057a8;
      16056: inst = 32'h8220000;
      16057: inst = 32'h10408000;
      16058: inst = 32'hc4057a9;
      16059: inst = 32'h8220000;
      16060: inst = 32'h10408000;
      16061: inst = 32'hc4057b6;
      16062: inst = 32'h8220000;
      16063: inst = 32'h10408000;
      16064: inst = 32'hc4057b7;
      16065: inst = 32'h8220000;
      16066: inst = 32'hc205aab;
      16067: inst = 32'h10408000;
      16068: inst = 32'hc405142;
      16069: inst = 32'h8220000;
      16070: inst = 32'h10408000;
      16071: inst = 32'hc40515d;
      16072: inst = 32'h8220000;
      16073: inst = 32'hc20cdd4;
      16074: inst = 32'h10408000;
      16075: inst = 32'hc40519e;
      16076: inst = 32'h8220000;
      16077: inst = 32'h10408000;
      16078: inst = 32'hc4051c1;
      16079: inst = 32'h8220000;
      16080: inst = 32'hc209471;
      16081: inst = 32'h10408000;
      16082: inst = 32'hc4051b6;
      16083: inst = 32'h8220000;
      16084: inst = 32'hc20de55;
      16085: inst = 32'h10408000;
      16086: inst = 32'hc4051fd;
      16087: inst = 32'h8220000;
      16088: inst = 32'h10408000;
      16089: inst = 32'hc405222;
      16090: inst = 32'h8220000;
      16091: inst = 32'hc209492;
      16092: inst = 32'h10408000;
      16093: inst = 32'hc4051fe;
      16094: inst = 32'h8220000;
      16095: inst = 32'h10408000;
      16096: inst = 32'hc405221;
      16097: inst = 32'h8220000;
      16098: inst = 32'hc205acc;
      16099: inst = 32'h10408000;
      16100: inst = 32'hc405201;
      16101: inst = 32'h8220000;
      16102: inst = 32'h10408000;
      16103: inst = 32'hc40521e;
      16104: inst = 32'h8220000;
      16105: inst = 32'h10408000;
      16106: inst = 32'hc405261;
      16107: inst = 32'h8220000;
      16108: inst = 32'h10408000;
      16109: inst = 32'hc40527e;
      16110: inst = 32'h8220000;
      16111: inst = 32'h10408000;
      16112: inst = 32'hc4052c1;
      16113: inst = 32'h8220000;
      16114: inst = 32'h10408000;
      16115: inst = 32'hc4052de;
      16116: inst = 32'h8220000;
      16117: inst = 32'hc20e696;
      16118: inst = 32'h10408000;
      16119: inst = 32'hc40525c;
      16120: inst = 32'h8220000;
      16121: inst = 32'h10408000;
      16122: inst = 32'hc405283;
      16123: inst = 32'h8220000;
      16124: inst = 32'hc209cb2;
      16125: inst = 32'h10408000;
      16126: inst = 32'hc40525d;
      16127: inst = 32'h8220000;
      16128: inst = 32'h10408000;
      16129: inst = 32'hc405282;
      16130: inst = 32'h8220000;
      16131: inst = 32'hc208c2f;
      16132: inst = 32'h10408000;
      16133: inst = 32'hc405269;
      16134: inst = 32'h8220000;
      16135: inst = 32'h10408000;
      16136: inst = 32'hc405276;
      16137: inst = 32'h8220000;
      16138: inst = 32'hc20ad33;
      16139: inst = 32'h10408000;
      16140: inst = 32'hc4052bc;
      16141: inst = 32'h8220000;
      16142: inst = 32'h10408000;
      16143: inst = 32'hc4052e3;
      16144: inst = 32'h8220000;
      16145: inst = 32'hc2083ee;
      16146: inst = 32'h10408000;
      16147: inst = 32'hc4052c9;
      16148: inst = 32'h8220000;
      16149: inst = 32'h10408000;
      16150: inst = 32'hc4052d6;
      16151: inst = 32'h8220000;
      16152: inst = 32'hc206b50;
      16153: inst = 32'h10408000;
      16154: inst = 32'hc405300;
      16155: inst = 32'h8220000;
      16156: inst = 32'h10408000;
      16157: inst = 32'hc405301;
      16158: inst = 32'h8220000;
      16159: inst = 32'h10408000;
      16160: inst = 32'hc405302;
      16161: inst = 32'h8220000;
      16162: inst = 32'h10408000;
      16163: inst = 32'hc405303;
      16164: inst = 32'h8220000;
      16165: inst = 32'h10408000;
      16166: inst = 32'hc405304;
      16167: inst = 32'h8220000;
      16168: inst = 32'h10408000;
      16169: inst = 32'hc405305;
      16170: inst = 32'h8220000;
      16171: inst = 32'h10408000;
      16172: inst = 32'hc405306;
      16173: inst = 32'h8220000;
      16174: inst = 32'h10408000;
      16175: inst = 32'hc405307;
      16176: inst = 32'h8220000;
      16177: inst = 32'h10408000;
      16178: inst = 32'hc405308;
      16179: inst = 32'h8220000;
      16180: inst = 32'h10408000;
      16181: inst = 32'hc405309;
      16182: inst = 32'h8220000;
      16183: inst = 32'h10408000;
      16184: inst = 32'hc40530a;
      16185: inst = 32'h8220000;
      16186: inst = 32'h10408000;
      16187: inst = 32'hc40530b;
      16188: inst = 32'h8220000;
      16189: inst = 32'h10408000;
      16190: inst = 32'hc40530c;
      16191: inst = 32'h8220000;
      16192: inst = 32'h10408000;
      16193: inst = 32'hc40530d;
      16194: inst = 32'h8220000;
      16195: inst = 32'h10408000;
      16196: inst = 32'hc40530e;
      16197: inst = 32'h8220000;
      16198: inst = 32'h10408000;
      16199: inst = 32'hc40530f;
      16200: inst = 32'h8220000;
      16201: inst = 32'h10408000;
      16202: inst = 32'hc405310;
      16203: inst = 32'h8220000;
      16204: inst = 32'h10408000;
      16205: inst = 32'hc405311;
      16206: inst = 32'h8220000;
      16207: inst = 32'h10408000;
      16208: inst = 32'hc405312;
      16209: inst = 32'h8220000;
      16210: inst = 32'h10408000;
      16211: inst = 32'hc405313;
      16212: inst = 32'h8220000;
      16213: inst = 32'h10408000;
      16214: inst = 32'hc405314;
      16215: inst = 32'h8220000;
      16216: inst = 32'h10408000;
      16217: inst = 32'hc405315;
      16218: inst = 32'h8220000;
      16219: inst = 32'h10408000;
      16220: inst = 32'hc405316;
      16221: inst = 32'h8220000;
      16222: inst = 32'h10408000;
      16223: inst = 32'hc405317;
      16224: inst = 32'h8220000;
      16225: inst = 32'h10408000;
      16226: inst = 32'hc405318;
      16227: inst = 32'h8220000;
      16228: inst = 32'h10408000;
      16229: inst = 32'hc405319;
      16230: inst = 32'h8220000;
      16231: inst = 32'h10408000;
      16232: inst = 32'hc40531a;
      16233: inst = 32'h8220000;
      16234: inst = 32'h10408000;
      16235: inst = 32'hc40532a;
      16236: inst = 32'h8220000;
      16237: inst = 32'h10408000;
      16238: inst = 32'hc40532b;
      16239: inst = 32'h8220000;
      16240: inst = 32'h10408000;
      16241: inst = 32'hc40532c;
      16242: inst = 32'h8220000;
      16243: inst = 32'h10408000;
      16244: inst = 32'hc40532d;
      16245: inst = 32'h8220000;
      16246: inst = 32'h10408000;
      16247: inst = 32'hc40532e;
      16248: inst = 32'h8220000;
      16249: inst = 32'h10408000;
      16250: inst = 32'hc40532f;
      16251: inst = 32'h8220000;
      16252: inst = 32'h10408000;
      16253: inst = 32'hc405330;
      16254: inst = 32'h8220000;
      16255: inst = 32'h10408000;
      16256: inst = 32'hc405331;
      16257: inst = 32'h8220000;
      16258: inst = 32'h10408000;
      16259: inst = 32'hc405332;
      16260: inst = 32'h8220000;
      16261: inst = 32'h10408000;
      16262: inst = 32'hc405333;
      16263: inst = 32'h8220000;
      16264: inst = 32'h10408000;
      16265: inst = 32'hc405334;
      16266: inst = 32'h8220000;
      16267: inst = 32'h10408000;
      16268: inst = 32'hc405335;
      16269: inst = 32'h8220000;
      16270: inst = 32'h10408000;
      16271: inst = 32'hc405345;
      16272: inst = 32'h8220000;
      16273: inst = 32'h10408000;
      16274: inst = 32'hc405346;
      16275: inst = 32'h8220000;
      16276: inst = 32'h10408000;
      16277: inst = 32'hc405347;
      16278: inst = 32'h8220000;
      16279: inst = 32'h10408000;
      16280: inst = 32'hc405348;
      16281: inst = 32'h8220000;
      16282: inst = 32'h10408000;
      16283: inst = 32'hc405349;
      16284: inst = 32'h8220000;
      16285: inst = 32'h10408000;
      16286: inst = 32'hc40534a;
      16287: inst = 32'h8220000;
      16288: inst = 32'h10408000;
      16289: inst = 32'hc40534b;
      16290: inst = 32'h8220000;
      16291: inst = 32'h10408000;
      16292: inst = 32'hc40534c;
      16293: inst = 32'h8220000;
      16294: inst = 32'h10408000;
      16295: inst = 32'hc40534d;
      16296: inst = 32'h8220000;
      16297: inst = 32'h10408000;
      16298: inst = 32'hc40534e;
      16299: inst = 32'h8220000;
      16300: inst = 32'h10408000;
      16301: inst = 32'hc40534f;
      16302: inst = 32'h8220000;
      16303: inst = 32'h10408000;
      16304: inst = 32'hc405350;
      16305: inst = 32'h8220000;
      16306: inst = 32'h10408000;
      16307: inst = 32'hc405351;
      16308: inst = 32'h8220000;
      16309: inst = 32'h10408000;
      16310: inst = 32'hc405352;
      16311: inst = 32'h8220000;
      16312: inst = 32'h10408000;
      16313: inst = 32'hc405353;
      16314: inst = 32'h8220000;
      16315: inst = 32'h10408000;
      16316: inst = 32'hc405354;
      16317: inst = 32'h8220000;
      16318: inst = 32'h10408000;
      16319: inst = 32'hc405355;
      16320: inst = 32'h8220000;
      16321: inst = 32'h10408000;
      16322: inst = 32'hc405356;
      16323: inst = 32'h8220000;
      16324: inst = 32'h10408000;
      16325: inst = 32'hc405357;
      16326: inst = 32'h8220000;
      16327: inst = 32'h10408000;
      16328: inst = 32'hc405358;
      16329: inst = 32'h8220000;
      16330: inst = 32'h10408000;
      16331: inst = 32'hc405359;
      16332: inst = 32'h8220000;
      16333: inst = 32'h10408000;
      16334: inst = 32'hc40535a;
      16335: inst = 32'h8220000;
      16336: inst = 32'h10408000;
      16337: inst = 32'hc40535b;
      16338: inst = 32'h8220000;
      16339: inst = 32'h10408000;
      16340: inst = 32'hc40535c;
      16341: inst = 32'h8220000;
      16342: inst = 32'h10408000;
      16343: inst = 32'hc40535d;
      16344: inst = 32'h8220000;
      16345: inst = 32'h10408000;
      16346: inst = 32'hc40535e;
      16347: inst = 32'h8220000;
      16348: inst = 32'h10408000;
      16349: inst = 32'hc40535f;
      16350: inst = 32'h8220000;
      16351: inst = 32'h10408000;
      16352: inst = 32'hc405360;
      16353: inst = 32'h8220000;
      16354: inst = 32'h10408000;
      16355: inst = 32'hc405361;
      16356: inst = 32'h8220000;
      16357: inst = 32'h10408000;
      16358: inst = 32'hc405362;
      16359: inst = 32'h8220000;
      16360: inst = 32'h10408000;
      16361: inst = 32'hc405363;
      16362: inst = 32'h8220000;
      16363: inst = 32'h10408000;
      16364: inst = 32'hc405364;
      16365: inst = 32'h8220000;
      16366: inst = 32'h10408000;
      16367: inst = 32'hc405365;
      16368: inst = 32'h8220000;
      16369: inst = 32'h10408000;
      16370: inst = 32'hc405366;
      16371: inst = 32'h8220000;
      16372: inst = 32'h10408000;
      16373: inst = 32'hc405367;
      16374: inst = 32'h8220000;
      16375: inst = 32'h10408000;
      16376: inst = 32'hc405368;
      16377: inst = 32'h8220000;
      16378: inst = 32'h10408000;
      16379: inst = 32'hc405369;
      16380: inst = 32'h8220000;
      16381: inst = 32'h10408000;
      16382: inst = 32'hc40536a;
      16383: inst = 32'h8220000;
      16384: inst = 32'h10408000;
      16385: inst = 32'hc40536b;
      16386: inst = 32'h8220000;
      16387: inst = 32'h10408000;
      16388: inst = 32'hc40536c;
      16389: inst = 32'h8220000;
      16390: inst = 32'h10408000;
      16391: inst = 32'hc40536d;
      16392: inst = 32'h8220000;
      16393: inst = 32'h10408000;
      16394: inst = 32'hc40536e;
      16395: inst = 32'h8220000;
      16396: inst = 32'h10408000;
      16397: inst = 32'hc40536f;
      16398: inst = 32'h8220000;
      16399: inst = 32'h10408000;
      16400: inst = 32'hc405370;
      16401: inst = 32'h8220000;
      16402: inst = 32'h10408000;
      16403: inst = 32'hc405371;
      16404: inst = 32'h8220000;
      16405: inst = 32'h10408000;
      16406: inst = 32'hc405372;
      16407: inst = 32'h8220000;
      16408: inst = 32'h10408000;
      16409: inst = 32'hc405373;
      16410: inst = 32'h8220000;
      16411: inst = 32'h10408000;
      16412: inst = 32'hc405374;
      16413: inst = 32'h8220000;
      16414: inst = 32'h10408000;
      16415: inst = 32'hc405375;
      16416: inst = 32'h8220000;
      16417: inst = 32'h10408000;
      16418: inst = 32'hc405376;
      16419: inst = 32'h8220000;
      16420: inst = 32'h10408000;
      16421: inst = 32'hc405377;
      16422: inst = 32'h8220000;
      16423: inst = 32'h10408000;
      16424: inst = 32'hc405378;
      16425: inst = 32'h8220000;
      16426: inst = 32'h10408000;
      16427: inst = 32'hc405379;
      16428: inst = 32'h8220000;
      16429: inst = 32'h10408000;
      16430: inst = 32'hc40538a;
      16431: inst = 32'h8220000;
      16432: inst = 32'h10408000;
      16433: inst = 32'hc40538b;
      16434: inst = 32'h8220000;
      16435: inst = 32'h10408000;
      16436: inst = 32'hc40538c;
      16437: inst = 32'h8220000;
      16438: inst = 32'h10408000;
      16439: inst = 32'hc40538d;
      16440: inst = 32'h8220000;
      16441: inst = 32'h10408000;
      16442: inst = 32'hc40538e;
      16443: inst = 32'h8220000;
      16444: inst = 32'h10408000;
      16445: inst = 32'hc40538f;
      16446: inst = 32'h8220000;
      16447: inst = 32'h10408000;
      16448: inst = 32'hc405390;
      16449: inst = 32'h8220000;
      16450: inst = 32'h10408000;
      16451: inst = 32'hc405391;
      16452: inst = 32'h8220000;
      16453: inst = 32'h10408000;
      16454: inst = 32'hc405392;
      16455: inst = 32'h8220000;
      16456: inst = 32'h10408000;
      16457: inst = 32'hc405393;
      16458: inst = 32'h8220000;
      16459: inst = 32'h10408000;
      16460: inst = 32'hc405394;
      16461: inst = 32'h8220000;
      16462: inst = 32'h10408000;
      16463: inst = 32'hc405395;
      16464: inst = 32'h8220000;
      16465: inst = 32'h10408000;
      16466: inst = 32'hc4053a6;
      16467: inst = 32'h8220000;
      16468: inst = 32'h10408000;
      16469: inst = 32'hc4053a7;
      16470: inst = 32'h8220000;
      16471: inst = 32'h10408000;
      16472: inst = 32'hc4053a8;
      16473: inst = 32'h8220000;
      16474: inst = 32'h10408000;
      16475: inst = 32'hc4053a9;
      16476: inst = 32'h8220000;
      16477: inst = 32'h10408000;
      16478: inst = 32'hc4053aa;
      16479: inst = 32'h8220000;
      16480: inst = 32'h10408000;
      16481: inst = 32'hc4053ab;
      16482: inst = 32'h8220000;
      16483: inst = 32'h10408000;
      16484: inst = 32'hc4053ac;
      16485: inst = 32'h8220000;
      16486: inst = 32'h10408000;
      16487: inst = 32'hc4053ad;
      16488: inst = 32'h8220000;
      16489: inst = 32'h10408000;
      16490: inst = 32'hc4053ae;
      16491: inst = 32'h8220000;
      16492: inst = 32'h10408000;
      16493: inst = 32'hc4053af;
      16494: inst = 32'h8220000;
      16495: inst = 32'h10408000;
      16496: inst = 32'hc4053b0;
      16497: inst = 32'h8220000;
      16498: inst = 32'h10408000;
      16499: inst = 32'hc4053b1;
      16500: inst = 32'h8220000;
      16501: inst = 32'h10408000;
      16502: inst = 32'hc4053b2;
      16503: inst = 32'h8220000;
      16504: inst = 32'h10408000;
      16505: inst = 32'hc4053b3;
      16506: inst = 32'h8220000;
      16507: inst = 32'h10408000;
      16508: inst = 32'hc4053b4;
      16509: inst = 32'h8220000;
      16510: inst = 32'h10408000;
      16511: inst = 32'hc4053b5;
      16512: inst = 32'h8220000;
      16513: inst = 32'h10408000;
      16514: inst = 32'hc4053b6;
      16515: inst = 32'h8220000;
      16516: inst = 32'h10408000;
      16517: inst = 32'hc4053b7;
      16518: inst = 32'h8220000;
      16519: inst = 32'h10408000;
      16520: inst = 32'hc4053b8;
      16521: inst = 32'h8220000;
      16522: inst = 32'h10408000;
      16523: inst = 32'hc4053b9;
      16524: inst = 32'h8220000;
      16525: inst = 32'h10408000;
      16526: inst = 32'hc4053ba;
      16527: inst = 32'h8220000;
      16528: inst = 32'h10408000;
      16529: inst = 32'hc4053bb;
      16530: inst = 32'h8220000;
      16531: inst = 32'h10408000;
      16532: inst = 32'hc4053bc;
      16533: inst = 32'h8220000;
      16534: inst = 32'h10408000;
      16535: inst = 32'hc4053bd;
      16536: inst = 32'h8220000;
      16537: inst = 32'h10408000;
      16538: inst = 32'hc4053be;
      16539: inst = 32'h8220000;
      16540: inst = 32'h10408000;
      16541: inst = 32'hc4053bf;
      16542: inst = 32'h8220000;
      16543: inst = 32'h10408000;
      16544: inst = 32'hc4053c0;
      16545: inst = 32'h8220000;
      16546: inst = 32'h10408000;
      16547: inst = 32'hc4053c1;
      16548: inst = 32'h8220000;
      16549: inst = 32'h10408000;
      16550: inst = 32'hc4053c2;
      16551: inst = 32'h8220000;
      16552: inst = 32'h10408000;
      16553: inst = 32'hc4053c3;
      16554: inst = 32'h8220000;
      16555: inst = 32'h10408000;
      16556: inst = 32'hc4053c4;
      16557: inst = 32'h8220000;
      16558: inst = 32'h10408000;
      16559: inst = 32'hc4053c5;
      16560: inst = 32'h8220000;
      16561: inst = 32'h10408000;
      16562: inst = 32'hc4053c6;
      16563: inst = 32'h8220000;
      16564: inst = 32'h10408000;
      16565: inst = 32'hc4053c7;
      16566: inst = 32'h8220000;
      16567: inst = 32'h10408000;
      16568: inst = 32'hc4053c8;
      16569: inst = 32'h8220000;
      16570: inst = 32'h10408000;
      16571: inst = 32'hc4053c9;
      16572: inst = 32'h8220000;
      16573: inst = 32'h10408000;
      16574: inst = 32'hc4053ca;
      16575: inst = 32'h8220000;
      16576: inst = 32'h10408000;
      16577: inst = 32'hc4053cb;
      16578: inst = 32'h8220000;
      16579: inst = 32'h10408000;
      16580: inst = 32'hc4053cc;
      16581: inst = 32'h8220000;
      16582: inst = 32'h10408000;
      16583: inst = 32'hc4053cd;
      16584: inst = 32'h8220000;
      16585: inst = 32'h10408000;
      16586: inst = 32'hc4053ce;
      16587: inst = 32'h8220000;
      16588: inst = 32'h10408000;
      16589: inst = 32'hc4053cf;
      16590: inst = 32'h8220000;
      16591: inst = 32'h10408000;
      16592: inst = 32'hc4053d0;
      16593: inst = 32'h8220000;
      16594: inst = 32'h10408000;
      16595: inst = 32'hc4053d1;
      16596: inst = 32'h8220000;
      16597: inst = 32'h10408000;
      16598: inst = 32'hc4053d2;
      16599: inst = 32'h8220000;
      16600: inst = 32'h10408000;
      16601: inst = 32'hc4053d3;
      16602: inst = 32'h8220000;
      16603: inst = 32'h10408000;
      16604: inst = 32'hc4053d4;
      16605: inst = 32'h8220000;
      16606: inst = 32'h10408000;
      16607: inst = 32'hc4053d5;
      16608: inst = 32'h8220000;
      16609: inst = 32'h10408000;
      16610: inst = 32'hc4053d6;
      16611: inst = 32'h8220000;
      16612: inst = 32'h10408000;
      16613: inst = 32'hc4053d7;
      16614: inst = 32'h8220000;
      16615: inst = 32'h10408000;
      16616: inst = 32'hc4053d8;
      16617: inst = 32'h8220000;
      16618: inst = 32'h10408000;
      16619: inst = 32'hc4053ea;
      16620: inst = 32'h8220000;
      16621: inst = 32'h10408000;
      16622: inst = 32'hc4053eb;
      16623: inst = 32'h8220000;
      16624: inst = 32'h10408000;
      16625: inst = 32'hc4053ec;
      16626: inst = 32'h8220000;
      16627: inst = 32'h10408000;
      16628: inst = 32'hc4053ed;
      16629: inst = 32'h8220000;
      16630: inst = 32'h10408000;
      16631: inst = 32'hc4053ee;
      16632: inst = 32'h8220000;
      16633: inst = 32'h10408000;
      16634: inst = 32'hc4053ef;
      16635: inst = 32'h8220000;
      16636: inst = 32'h10408000;
      16637: inst = 32'hc4053f0;
      16638: inst = 32'h8220000;
      16639: inst = 32'h10408000;
      16640: inst = 32'hc4053f1;
      16641: inst = 32'h8220000;
      16642: inst = 32'h10408000;
      16643: inst = 32'hc4053f2;
      16644: inst = 32'h8220000;
      16645: inst = 32'h10408000;
      16646: inst = 32'hc4053f3;
      16647: inst = 32'h8220000;
      16648: inst = 32'h10408000;
      16649: inst = 32'hc4053f4;
      16650: inst = 32'h8220000;
      16651: inst = 32'h10408000;
      16652: inst = 32'hc4053f5;
      16653: inst = 32'h8220000;
      16654: inst = 32'h10408000;
      16655: inst = 32'hc405407;
      16656: inst = 32'h8220000;
      16657: inst = 32'h10408000;
      16658: inst = 32'hc405408;
      16659: inst = 32'h8220000;
      16660: inst = 32'h10408000;
      16661: inst = 32'hc405409;
      16662: inst = 32'h8220000;
      16663: inst = 32'h10408000;
      16664: inst = 32'hc40540a;
      16665: inst = 32'h8220000;
      16666: inst = 32'h10408000;
      16667: inst = 32'hc40540b;
      16668: inst = 32'h8220000;
      16669: inst = 32'h10408000;
      16670: inst = 32'hc40540c;
      16671: inst = 32'h8220000;
      16672: inst = 32'h10408000;
      16673: inst = 32'hc40540d;
      16674: inst = 32'h8220000;
      16675: inst = 32'h10408000;
      16676: inst = 32'hc40540e;
      16677: inst = 32'h8220000;
      16678: inst = 32'h10408000;
      16679: inst = 32'hc40540f;
      16680: inst = 32'h8220000;
      16681: inst = 32'h10408000;
      16682: inst = 32'hc405410;
      16683: inst = 32'h8220000;
      16684: inst = 32'h10408000;
      16685: inst = 32'hc405411;
      16686: inst = 32'h8220000;
      16687: inst = 32'h10408000;
      16688: inst = 32'hc405412;
      16689: inst = 32'h8220000;
      16690: inst = 32'h10408000;
      16691: inst = 32'hc405413;
      16692: inst = 32'h8220000;
      16693: inst = 32'h10408000;
      16694: inst = 32'hc405414;
      16695: inst = 32'h8220000;
      16696: inst = 32'h10408000;
      16697: inst = 32'hc405415;
      16698: inst = 32'h8220000;
      16699: inst = 32'h10408000;
      16700: inst = 32'hc405416;
      16701: inst = 32'h8220000;
      16702: inst = 32'h10408000;
      16703: inst = 32'hc405417;
      16704: inst = 32'h8220000;
      16705: inst = 32'h10408000;
      16706: inst = 32'hc405418;
      16707: inst = 32'h8220000;
      16708: inst = 32'h10408000;
      16709: inst = 32'hc405419;
      16710: inst = 32'h8220000;
      16711: inst = 32'h10408000;
      16712: inst = 32'hc40541a;
      16713: inst = 32'h8220000;
      16714: inst = 32'h10408000;
      16715: inst = 32'hc40541b;
      16716: inst = 32'h8220000;
      16717: inst = 32'h10408000;
      16718: inst = 32'hc40541c;
      16719: inst = 32'h8220000;
      16720: inst = 32'h10408000;
      16721: inst = 32'hc40541d;
      16722: inst = 32'h8220000;
      16723: inst = 32'h10408000;
      16724: inst = 32'hc40541e;
      16725: inst = 32'h8220000;
      16726: inst = 32'h10408000;
      16727: inst = 32'hc40541f;
      16728: inst = 32'h8220000;
      16729: inst = 32'h10408000;
      16730: inst = 32'hc405420;
      16731: inst = 32'h8220000;
      16732: inst = 32'h10408000;
      16733: inst = 32'hc405421;
      16734: inst = 32'h8220000;
      16735: inst = 32'h10408000;
      16736: inst = 32'hc405422;
      16737: inst = 32'h8220000;
      16738: inst = 32'h10408000;
      16739: inst = 32'hc405423;
      16740: inst = 32'h8220000;
      16741: inst = 32'h10408000;
      16742: inst = 32'hc405424;
      16743: inst = 32'h8220000;
      16744: inst = 32'h10408000;
      16745: inst = 32'hc405425;
      16746: inst = 32'h8220000;
      16747: inst = 32'h10408000;
      16748: inst = 32'hc405426;
      16749: inst = 32'h8220000;
      16750: inst = 32'h10408000;
      16751: inst = 32'hc405427;
      16752: inst = 32'h8220000;
      16753: inst = 32'h10408000;
      16754: inst = 32'hc405428;
      16755: inst = 32'h8220000;
      16756: inst = 32'h10408000;
      16757: inst = 32'hc405429;
      16758: inst = 32'h8220000;
      16759: inst = 32'h10408000;
      16760: inst = 32'hc40542a;
      16761: inst = 32'h8220000;
      16762: inst = 32'h10408000;
      16763: inst = 32'hc40542b;
      16764: inst = 32'h8220000;
      16765: inst = 32'h10408000;
      16766: inst = 32'hc40542c;
      16767: inst = 32'h8220000;
      16768: inst = 32'h10408000;
      16769: inst = 32'hc40542d;
      16770: inst = 32'h8220000;
      16771: inst = 32'h10408000;
      16772: inst = 32'hc40542e;
      16773: inst = 32'h8220000;
      16774: inst = 32'h10408000;
      16775: inst = 32'hc40542f;
      16776: inst = 32'h8220000;
      16777: inst = 32'h10408000;
      16778: inst = 32'hc405430;
      16779: inst = 32'h8220000;
      16780: inst = 32'h10408000;
      16781: inst = 32'hc405431;
      16782: inst = 32'h8220000;
      16783: inst = 32'h10408000;
      16784: inst = 32'hc405432;
      16785: inst = 32'h8220000;
      16786: inst = 32'h10408000;
      16787: inst = 32'hc405433;
      16788: inst = 32'h8220000;
      16789: inst = 32'h10408000;
      16790: inst = 32'hc405434;
      16791: inst = 32'h8220000;
      16792: inst = 32'h10408000;
      16793: inst = 32'hc405435;
      16794: inst = 32'h8220000;
      16795: inst = 32'h10408000;
      16796: inst = 32'hc405436;
      16797: inst = 32'h8220000;
      16798: inst = 32'h10408000;
      16799: inst = 32'hc405437;
      16800: inst = 32'h8220000;
      16801: inst = 32'h10408000;
      16802: inst = 32'hc405438;
      16803: inst = 32'h8220000;
      16804: inst = 32'h10408000;
      16805: inst = 32'hc40544a;
      16806: inst = 32'h8220000;
      16807: inst = 32'h10408000;
      16808: inst = 32'hc40544b;
      16809: inst = 32'h8220000;
      16810: inst = 32'h10408000;
      16811: inst = 32'hc40544c;
      16812: inst = 32'h8220000;
      16813: inst = 32'h10408000;
      16814: inst = 32'hc40544d;
      16815: inst = 32'h8220000;
      16816: inst = 32'h10408000;
      16817: inst = 32'hc40544e;
      16818: inst = 32'h8220000;
      16819: inst = 32'h10408000;
      16820: inst = 32'hc40544f;
      16821: inst = 32'h8220000;
      16822: inst = 32'h10408000;
      16823: inst = 32'hc405450;
      16824: inst = 32'h8220000;
      16825: inst = 32'h10408000;
      16826: inst = 32'hc405451;
      16827: inst = 32'h8220000;
      16828: inst = 32'h10408000;
      16829: inst = 32'hc405452;
      16830: inst = 32'h8220000;
      16831: inst = 32'h10408000;
      16832: inst = 32'hc405453;
      16833: inst = 32'h8220000;
      16834: inst = 32'h10408000;
      16835: inst = 32'hc405454;
      16836: inst = 32'h8220000;
      16837: inst = 32'h10408000;
      16838: inst = 32'hc405455;
      16839: inst = 32'h8220000;
      16840: inst = 32'h10408000;
      16841: inst = 32'hc405467;
      16842: inst = 32'h8220000;
      16843: inst = 32'h10408000;
      16844: inst = 32'hc405468;
      16845: inst = 32'h8220000;
      16846: inst = 32'h10408000;
      16847: inst = 32'hc405469;
      16848: inst = 32'h8220000;
      16849: inst = 32'h10408000;
      16850: inst = 32'hc40546a;
      16851: inst = 32'h8220000;
      16852: inst = 32'h10408000;
      16853: inst = 32'hc40546b;
      16854: inst = 32'h8220000;
      16855: inst = 32'h10408000;
      16856: inst = 32'hc40546c;
      16857: inst = 32'h8220000;
      16858: inst = 32'h10408000;
      16859: inst = 32'hc40546d;
      16860: inst = 32'h8220000;
      16861: inst = 32'h10408000;
      16862: inst = 32'hc40546e;
      16863: inst = 32'h8220000;
      16864: inst = 32'h10408000;
      16865: inst = 32'hc40546f;
      16866: inst = 32'h8220000;
      16867: inst = 32'h10408000;
      16868: inst = 32'hc405470;
      16869: inst = 32'h8220000;
      16870: inst = 32'h10408000;
      16871: inst = 32'hc405471;
      16872: inst = 32'h8220000;
      16873: inst = 32'h10408000;
      16874: inst = 32'hc405472;
      16875: inst = 32'h8220000;
      16876: inst = 32'h10408000;
      16877: inst = 32'hc405473;
      16878: inst = 32'h8220000;
      16879: inst = 32'h10408000;
      16880: inst = 32'hc405474;
      16881: inst = 32'h8220000;
      16882: inst = 32'h10408000;
      16883: inst = 32'hc405475;
      16884: inst = 32'h8220000;
      16885: inst = 32'h10408000;
      16886: inst = 32'hc405476;
      16887: inst = 32'h8220000;
      16888: inst = 32'h10408000;
      16889: inst = 32'hc405477;
      16890: inst = 32'h8220000;
      16891: inst = 32'h10408000;
      16892: inst = 32'hc405478;
      16893: inst = 32'h8220000;
      16894: inst = 32'h10408000;
      16895: inst = 32'hc405479;
      16896: inst = 32'h8220000;
      16897: inst = 32'h10408000;
      16898: inst = 32'hc40547a;
      16899: inst = 32'h8220000;
      16900: inst = 32'h10408000;
      16901: inst = 32'hc40547b;
      16902: inst = 32'h8220000;
      16903: inst = 32'h10408000;
      16904: inst = 32'hc40547c;
      16905: inst = 32'h8220000;
      16906: inst = 32'h10408000;
      16907: inst = 32'hc40547d;
      16908: inst = 32'h8220000;
      16909: inst = 32'h10408000;
      16910: inst = 32'hc40547e;
      16911: inst = 32'h8220000;
      16912: inst = 32'h10408000;
      16913: inst = 32'hc40547f;
      16914: inst = 32'h8220000;
      16915: inst = 32'h10408000;
      16916: inst = 32'hc405480;
      16917: inst = 32'h8220000;
      16918: inst = 32'h10408000;
      16919: inst = 32'hc405481;
      16920: inst = 32'h8220000;
      16921: inst = 32'h10408000;
      16922: inst = 32'hc405482;
      16923: inst = 32'h8220000;
      16924: inst = 32'h10408000;
      16925: inst = 32'hc405483;
      16926: inst = 32'h8220000;
      16927: inst = 32'h10408000;
      16928: inst = 32'hc405484;
      16929: inst = 32'h8220000;
      16930: inst = 32'h10408000;
      16931: inst = 32'hc405485;
      16932: inst = 32'h8220000;
      16933: inst = 32'h10408000;
      16934: inst = 32'hc405486;
      16935: inst = 32'h8220000;
      16936: inst = 32'h10408000;
      16937: inst = 32'hc405487;
      16938: inst = 32'h8220000;
      16939: inst = 32'h10408000;
      16940: inst = 32'hc405488;
      16941: inst = 32'h8220000;
      16942: inst = 32'h10408000;
      16943: inst = 32'hc405489;
      16944: inst = 32'h8220000;
      16945: inst = 32'h10408000;
      16946: inst = 32'hc40548a;
      16947: inst = 32'h8220000;
      16948: inst = 32'h10408000;
      16949: inst = 32'hc40548b;
      16950: inst = 32'h8220000;
      16951: inst = 32'h10408000;
      16952: inst = 32'hc40548c;
      16953: inst = 32'h8220000;
      16954: inst = 32'h10408000;
      16955: inst = 32'hc40548d;
      16956: inst = 32'h8220000;
      16957: inst = 32'h10408000;
      16958: inst = 32'hc40548e;
      16959: inst = 32'h8220000;
      16960: inst = 32'h10408000;
      16961: inst = 32'hc40548f;
      16962: inst = 32'h8220000;
      16963: inst = 32'h10408000;
      16964: inst = 32'hc405490;
      16965: inst = 32'h8220000;
      16966: inst = 32'h10408000;
      16967: inst = 32'hc405491;
      16968: inst = 32'h8220000;
      16969: inst = 32'h10408000;
      16970: inst = 32'hc405492;
      16971: inst = 32'h8220000;
      16972: inst = 32'h10408000;
      16973: inst = 32'hc405493;
      16974: inst = 32'h8220000;
      16975: inst = 32'h10408000;
      16976: inst = 32'hc405494;
      16977: inst = 32'h8220000;
      16978: inst = 32'h10408000;
      16979: inst = 32'hc405495;
      16980: inst = 32'h8220000;
      16981: inst = 32'h10408000;
      16982: inst = 32'hc405496;
      16983: inst = 32'h8220000;
      16984: inst = 32'h10408000;
      16985: inst = 32'hc405497;
      16986: inst = 32'h8220000;
      16987: inst = 32'h10408000;
      16988: inst = 32'hc4054aa;
      16989: inst = 32'h8220000;
      16990: inst = 32'h10408000;
      16991: inst = 32'hc4054ab;
      16992: inst = 32'h8220000;
      16993: inst = 32'h10408000;
      16994: inst = 32'hc4054ac;
      16995: inst = 32'h8220000;
      16996: inst = 32'h10408000;
      16997: inst = 32'hc4054ad;
      16998: inst = 32'h8220000;
      16999: inst = 32'h10408000;
      17000: inst = 32'hc4054ae;
      17001: inst = 32'h8220000;
      17002: inst = 32'h10408000;
      17003: inst = 32'hc4054af;
      17004: inst = 32'h8220000;
      17005: inst = 32'h10408000;
      17006: inst = 32'hc4054b0;
      17007: inst = 32'h8220000;
      17008: inst = 32'h10408000;
      17009: inst = 32'hc4054b1;
      17010: inst = 32'h8220000;
      17011: inst = 32'h10408000;
      17012: inst = 32'hc4054b2;
      17013: inst = 32'h8220000;
      17014: inst = 32'h10408000;
      17015: inst = 32'hc4054b3;
      17016: inst = 32'h8220000;
      17017: inst = 32'h10408000;
      17018: inst = 32'hc4054b4;
      17019: inst = 32'h8220000;
      17020: inst = 32'h10408000;
      17021: inst = 32'hc4054b5;
      17022: inst = 32'h8220000;
      17023: inst = 32'h10408000;
      17024: inst = 32'hc4054c8;
      17025: inst = 32'h8220000;
      17026: inst = 32'h10408000;
      17027: inst = 32'hc4054c9;
      17028: inst = 32'h8220000;
      17029: inst = 32'h10408000;
      17030: inst = 32'hc4054ca;
      17031: inst = 32'h8220000;
      17032: inst = 32'h10408000;
      17033: inst = 32'hc4054cb;
      17034: inst = 32'h8220000;
      17035: inst = 32'h10408000;
      17036: inst = 32'hc4054cc;
      17037: inst = 32'h8220000;
      17038: inst = 32'h10408000;
      17039: inst = 32'hc4054cd;
      17040: inst = 32'h8220000;
      17041: inst = 32'h10408000;
      17042: inst = 32'hc4054ce;
      17043: inst = 32'h8220000;
      17044: inst = 32'h10408000;
      17045: inst = 32'hc4054cf;
      17046: inst = 32'h8220000;
      17047: inst = 32'h10408000;
      17048: inst = 32'hc4054d0;
      17049: inst = 32'h8220000;
      17050: inst = 32'h10408000;
      17051: inst = 32'hc4054d1;
      17052: inst = 32'h8220000;
      17053: inst = 32'h10408000;
      17054: inst = 32'hc4054d2;
      17055: inst = 32'h8220000;
      17056: inst = 32'h10408000;
      17057: inst = 32'hc4054d3;
      17058: inst = 32'h8220000;
      17059: inst = 32'h10408000;
      17060: inst = 32'hc4054d4;
      17061: inst = 32'h8220000;
      17062: inst = 32'h10408000;
      17063: inst = 32'hc4054d5;
      17064: inst = 32'h8220000;
      17065: inst = 32'h10408000;
      17066: inst = 32'hc4054d6;
      17067: inst = 32'h8220000;
      17068: inst = 32'h10408000;
      17069: inst = 32'hc4054d7;
      17070: inst = 32'h8220000;
      17071: inst = 32'h10408000;
      17072: inst = 32'hc4054d8;
      17073: inst = 32'h8220000;
      17074: inst = 32'h10408000;
      17075: inst = 32'hc4054d9;
      17076: inst = 32'h8220000;
      17077: inst = 32'h10408000;
      17078: inst = 32'hc4054da;
      17079: inst = 32'h8220000;
      17080: inst = 32'h10408000;
      17081: inst = 32'hc4054db;
      17082: inst = 32'h8220000;
      17083: inst = 32'h10408000;
      17084: inst = 32'hc4054dc;
      17085: inst = 32'h8220000;
      17086: inst = 32'h10408000;
      17087: inst = 32'hc4054dd;
      17088: inst = 32'h8220000;
      17089: inst = 32'h10408000;
      17090: inst = 32'hc4054de;
      17091: inst = 32'h8220000;
      17092: inst = 32'h10408000;
      17093: inst = 32'hc4054df;
      17094: inst = 32'h8220000;
      17095: inst = 32'h10408000;
      17096: inst = 32'hc4054e0;
      17097: inst = 32'h8220000;
      17098: inst = 32'h10408000;
      17099: inst = 32'hc4054e1;
      17100: inst = 32'h8220000;
      17101: inst = 32'h10408000;
      17102: inst = 32'hc4054e2;
      17103: inst = 32'h8220000;
      17104: inst = 32'h10408000;
      17105: inst = 32'hc4054e3;
      17106: inst = 32'h8220000;
      17107: inst = 32'h10408000;
      17108: inst = 32'hc4054e4;
      17109: inst = 32'h8220000;
      17110: inst = 32'h10408000;
      17111: inst = 32'hc4054e5;
      17112: inst = 32'h8220000;
      17113: inst = 32'h10408000;
      17114: inst = 32'hc4054e6;
      17115: inst = 32'h8220000;
      17116: inst = 32'h10408000;
      17117: inst = 32'hc4054e7;
      17118: inst = 32'h8220000;
      17119: inst = 32'h10408000;
      17120: inst = 32'hc4054e8;
      17121: inst = 32'h8220000;
      17122: inst = 32'h10408000;
      17123: inst = 32'hc4054e9;
      17124: inst = 32'h8220000;
      17125: inst = 32'h10408000;
      17126: inst = 32'hc4054ea;
      17127: inst = 32'h8220000;
      17128: inst = 32'h10408000;
      17129: inst = 32'hc4054eb;
      17130: inst = 32'h8220000;
      17131: inst = 32'h10408000;
      17132: inst = 32'hc4054ec;
      17133: inst = 32'h8220000;
      17134: inst = 32'h10408000;
      17135: inst = 32'hc4054ed;
      17136: inst = 32'h8220000;
      17137: inst = 32'h10408000;
      17138: inst = 32'hc4054ee;
      17139: inst = 32'h8220000;
      17140: inst = 32'h10408000;
      17141: inst = 32'hc4054ef;
      17142: inst = 32'h8220000;
      17143: inst = 32'h10408000;
      17144: inst = 32'hc4054f0;
      17145: inst = 32'h8220000;
      17146: inst = 32'h10408000;
      17147: inst = 32'hc4054f1;
      17148: inst = 32'h8220000;
      17149: inst = 32'h10408000;
      17150: inst = 32'hc4054f2;
      17151: inst = 32'h8220000;
      17152: inst = 32'h10408000;
      17153: inst = 32'hc4054f3;
      17154: inst = 32'h8220000;
      17155: inst = 32'h10408000;
      17156: inst = 32'hc4054f4;
      17157: inst = 32'h8220000;
      17158: inst = 32'h10408000;
      17159: inst = 32'hc4054f5;
      17160: inst = 32'h8220000;
      17161: inst = 32'h10408000;
      17162: inst = 32'hc4054f6;
      17163: inst = 32'h8220000;
      17164: inst = 32'h10408000;
      17165: inst = 32'hc40550a;
      17166: inst = 32'h8220000;
      17167: inst = 32'h10408000;
      17168: inst = 32'hc40550b;
      17169: inst = 32'h8220000;
      17170: inst = 32'h10408000;
      17171: inst = 32'hc40550c;
      17172: inst = 32'h8220000;
      17173: inst = 32'h10408000;
      17174: inst = 32'hc40550d;
      17175: inst = 32'h8220000;
      17176: inst = 32'h10408000;
      17177: inst = 32'hc40550e;
      17178: inst = 32'h8220000;
      17179: inst = 32'h10408000;
      17180: inst = 32'hc40550f;
      17181: inst = 32'h8220000;
      17182: inst = 32'h10408000;
      17183: inst = 32'hc405510;
      17184: inst = 32'h8220000;
      17185: inst = 32'h10408000;
      17186: inst = 32'hc405511;
      17187: inst = 32'h8220000;
      17188: inst = 32'h10408000;
      17189: inst = 32'hc405512;
      17190: inst = 32'h8220000;
      17191: inst = 32'h10408000;
      17192: inst = 32'hc405513;
      17193: inst = 32'h8220000;
      17194: inst = 32'h10408000;
      17195: inst = 32'hc405514;
      17196: inst = 32'h8220000;
      17197: inst = 32'h10408000;
      17198: inst = 32'hc405515;
      17199: inst = 32'h8220000;
      17200: inst = 32'h10408000;
      17201: inst = 32'hc405529;
      17202: inst = 32'h8220000;
      17203: inst = 32'h10408000;
      17204: inst = 32'hc40552a;
      17205: inst = 32'h8220000;
      17206: inst = 32'h10408000;
      17207: inst = 32'hc40552b;
      17208: inst = 32'h8220000;
      17209: inst = 32'h10408000;
      17210: inst = 32'hc40552c;
      17211: inst = 32'h8220000;
      17212: inst = 32'h10408000;
      17213: inst = 32'hc40552d;
      17214: inst = 32'h8220000;
      17215: inst = 32'h10408000;
      17216: inst = 32'hc40552e;
      17217: inst = 32'h8220000;
      17218: inst = 32'h10408000;
      17219: inst = 32'hc40552f;
      17220: inst = 32'h8220000;
      17221: inst = 32'h10408000;
      17222: inst = 32'hc405530;
      17223: inst = 32'h8220000;
      17224: inst = 32'h10408000;
      17225: inst = 32'hc405531;
      17226: inst = 32'h8220000;
      17227: inst = 32'h10408000;
      17228: inst = 32'hc405532;
      17229: inst = 32'h8220000;
      17230: inst = 32'h10408000;
      17231: inst = 32'hc405533;
      17232: inst = 32'h8220000;
      17233: inst = 32'h10408000;
      17234: inst = 32'hc405534;
      17235: inst = 32'h8220000;
      17236: inst = 32'h10408000;
      17237: inst = 32'hc405535;
      17238: inst = 32'h8220000;
      17239: inst = 32'h10408000;
      17240: inst = 32'hc405536;
      17241: inst = 32'h8220000;
      17242: inst = 32'h10408000;
      17243: inst = 32'hc405537;
      17244: inst = 32'h8220000;
      17245: inst = 32'h10408000;
      17246: inst = 32'hc405538;
      17247: inst = 32'h8220000;
      17248: inst = 32'h10408000;
      17249: inst = 32'hc405539;
      17250: inst = 32'h8220000;
      17251: inst = 32'h10408000;
      17252: inst = 32'hc40553a;
      17253: inst = 32'h8220000;
      17254: inst = 32'h10408000;
      17255: inst = 32'hc40553b;
      17256: inst = 32'h8220000;
      17257: inst = 32'h10408000;
      17258: inst = 32'hc40553c;
      17259: inst = 32'h8220000;
      17260: inst = 32'h10408000;
      17261: inst = 32'hc40553d;
      17262: inst = 32'h8220000;
      17263: inst = 32'h10408000;
      17264: inst = 32'hc40553e;
      17265: inst = 32'h8220000;
      17266: inst = 32'h10408000;
      17267: inst = 32'hc40553f;
      17268: inst = 32'h8220000;
      17269: inst = 32'h10408000;
      17270: inst = 32'hc405540;
      17271: inst = 32'h8220000;
      17272: inst = 32'h10408000;
      17273: inst = 32'hc405541;
      17274: inst = 32'h8220000;
      17275: inst = 32'h10408000;
      17276: inst = 32'hc405542;
      17277: inst = 32'h8220000;
      17278: inst = 32'h10408000;
      17279: inst = 32'hc405543;
      17280: inst = 32'h8220000;
      17281: inst = 32'h10408000;
      17282: inst = 32'hc405544;
      17283: inst = 32'h8220000;
      17284: inst = 32'h10408000;
      17285: inst = 32'hc405545;
      17286: inst = 32'h8220000;
      17287: inst = 32'h10408000;
      17288: inst = 32'hc405546;
      17289: inst = 32'h8220000;
      17290: inst = 32'h10408000;
      17291: inst = 32'hc405547;
      17292: inst = 32'h8220000;
      17293: inst = 32'h10408000;
      17294: inst = 32'hc405548;
      17295: inst = 32'h8220000;
      17296: inst = 32'h10408000;
      17297: inst = 32'hc405549;
      17298: inst = 32'h8220000;
      17299: inst = 32'h10408000;
      17300: inst = 32'hc40554a;
      17301: inst = 32'h8220000;
      17302: inst = 32'h10408000;
      17303: inst = 32'hc40554b;
      17304: inst = 32'h8220000;
      17305: inst = 32'h10408000;
      17306: inst = 32'hc40554c;
      17307: inst = 32'h8220000;
      17308: inst = 32'h10408000;
      17309: inst = 32'hc40554d;
      17310: inst = 32'h8220000;
      17311: inst = 32'h10408000;
      17312: inst = 32'hc40554e;
      17313: inst = 32'h8220000;
      17314: inst = 32'h10408000;
      17315: inst = 32'hc40554f;
      17316: inst = 32'h8220000;
      17317: inst = 32'h10408000;
      17318: inst = 32'hc405550;
      17319: inst = 32'h8220000;
      17320: inst = 32'h10408000;
      17321: inst = 32'hc405551;
      17322: inst = 32'h8220000;
      17323: inst = 32'h10408000;
      17324: inst = 32'hc405552;
      17325: inst = 32'h8220000;
      17326: inst = 32'h10408000;
      17327: inst = 32'hc405553;
      17328: inst = 32'h8220000;
      17329: inst = 32'h10408000;
      17330: inst = 32'hc405554;
      17331: inst = 32'h8220000;
      17332: inst = 32'h10408000;
      17333: inst = 32'hc405555;
      17334: inst = 32'h8220000;
      17335: inst = 32'h10408000;
      17336: inst = 32'hc40556a;
      17337: inst = 32'h8220000;
      17338: inst = 32'h10408000;
      17339: inst = 32'hc40556b;
      17340: inst = 32'h8220000;
      17341: inst = 32'h10408000;
      17342: inst = 32'hc40556c;
      17343: inst = 32'h8220000;
      17344: inst = 32'h10408000;
      17345: inst = 32'hc40556d;
      17346: inst = 32'h8220000;
      17347: inst = 32'h10408000;
      17348: inst = 32'hc40556e;
      17349: inst = 32'h8220000;
      17350: inst = 32'h10408000;
      17351: inst = 32'hc40556f;
      17352: inst = 32'h8220000;
      17353: inst = 32'h10408000;
      17354: inst = 32'hc405570;
      17355: inst = 32'h8220000;
      17356: inst = 32'h10408000;
      17357: inst = 32'hc405571;
      17358: inst = 32'h8220000;
      17359: inst = 32'h10408000;
      17360: inst = 32'hc405572;
      17361: inst = 32'h8220000;
      17362: inst = 32'h10408000;
      17363: inst = 32'hc405573;
      17364: inst = 32'h8220000;
      17365: inst = 32'h10408000;
      17366: inst = 32'hc405574;
      17367: inst = 32'h8220000;
      17368: inst = 32'h10408000;
      17369: inst = 32'hc405575;
      17370: inst = 32'h8220000;
      17371: inst = 32'h10408000;
      17372: inst = 32'hc40558a;
      17373: inst = 32'h8220000;
      17374: inst = 32'h10408000;
      17375: inst = 32'hc40558b;
      17376: inst = 32'h8220000;
      17377: inst = 32'h10408000;
      17378: inst = 32'hc40558c;
      17379: inst = 32'h8220000;
      17380: inst = 32'h10408000;
      17381: inst = 32'hc40558d;
      17382: inst = 32'h8220000;
      17383: inst = 32'h10408000;
      17384: inst = 32'hc40558e;
      17385: inst = 32'h8220000;
      17386: inst = 32'h10408000;
      17387: inst = 32'hc40558f;
      17388: inst = 32'h8220000;
      17389: inst = 32'h10408000;
      17390: inst = 32'hc405590;
      17391: inst = 32'h8220000;
      17392: inst = 32'h10408000;
      17393: inst = 32'hc405591;
      17394: inst = 32'h8220000;
      17395: inst = 32'h10408000;
      17396: inst = 32'hc405592;
      17397: inst = 32'h8220000;
      17398: inst = 32'h10408000;
      17399: inst = 32'hc405593;
      17400: inst = 32'h8220000;
      17401: inst = 32'h10408000;
      17402: inst = 32'hc405594;
      17403: inst = 32'h8220000;
      17404: inst = 32'h10408000;
      17405: inst = 32'hc405595;
      17406: inst = 32'h8220000;
      17407: inst = 32'h10408000;
      17408: inst = 32'hc405596;
      17409: inst = 32'h8220000;
      17410: inst = 32'h10408000;
      17411: inst = 32'hc405597;
      17412: inst = 32'h8220000;
      17413: inst = 32'h10408000;
      17414: inst = 32'hc405598;
      17415: inst = 32'h8220000;
      17416: inst = 32'h10408000;
      17417: inst = 32'hc405599;
      17418: inst = 32'h8220000;
      17419: inst = 32'h10408000;
      17420: inst = 32'hc40559a;
      17421: inst = 32'h8220000;
      17422: inst = 32'h10408000;
      17423: inst = 32'hc40559b;
      17424: inst = 32'h8220000;
      17425: inst = 32'h10408000;
      17426: inst = 32'hc40559c;
      17427: inst = 32'h8220000;
      17428: inst = 32'h10408000;
      17429: inst = 32'hc40559d;
      17430: inst = 32'h8220000;
      17431: inst = 32'h10408000;
      17432: inst = 32'hc40559e;
      17433: inst = 32'h8220000;
      17434: inst = 32'h10408000;
      17435: inst = 32'hc40559f;
      17436: inst = 32'h8220000;
      17437: inst = 32'h10408000;
      17438: inst = 32'hc4055a0;
      17439: inst = 32'h8220000;
      17440: inst = 32'h10408000;
      17441: inst = 32'hc4055a1;
      17442: inst = 32'h8220000;
      17443: inst = 32'h10408000;
      17444: inst = 32'hc4055a2;
      17445: inst = 32'h8220000;
      17446: inst = 32'h10408000;
      17447: inst = 32'hc4055a3;
      17448: inst = 32'h8220000;
      17449: inst = 32'h10408000;
      17450: inst = 32'hc4055a4;
      17451: inst = 32'h8220000;
      17452: inst = 32'h10408000;
      17453: inst = 32'hc4055a5;
      17454: inst = 32'h8220000;
      17455: inst = 32'h10408000;
      17456: inst = 32'hc4055a6;
      17457: inst = 32'h8220000;
      17458: inst = 32'h10408000;
      17459: inst = 32'hc4055a7;
      17460: inst = 32'h8220000;
      17461: inst = 32'h10408000;
      17462: inst = 32'hc4055a8;
      17463: inst = 32'h8220000;
      17464: inst = 32'h10408000;
      17465: inst = 32'hc4055a9;
      17466: inst = 32'h8220000;
      17467: inst = 32'h10408000;
      17468: inst = 32'hc4055aa;
      17469: inst = 32'h8220000;
      17470: inst = 32'h10408000;
      17471: inst = 32'hc4055ab;
      17472: inst = 32'h8220000;
      17473: inst = 32'h10408000;
      17474: inst = 32'hc4055ac;
      17475: inst = 32'h8220000;
      17476: inst = 32'h10408000;
      17477: inst = 32'hc4055ad;
      17478: inst = 32'h8220000;
      17479: inst = 32'h10408000;
      17480: inst = 32'hc4055ae;
      17481: inst = 32'h8220000;
      17482: inst = 32'h10408000;
      17483: inst = 32'hc4055af;
      17484: inst = 32'h8220000;
      17485: inst = 32'h10408000;
      17486: inst = 32'hc4055b0;
      17487: inst = 32'h8220000;
      17488: inst = 32'h10408000;
      17489: inst = 32'hc4055b1;
      17490: inst = 32'h8220000;
      17491: inst = 32'h10408000;
      17492: inst = 32'hc4055b2;
      17493: inst = 32'h8220000;
      17494: inst = 32'h10408000;
      17495: inst = 32'hc4055b3;
      17496: inst = 32'h8220000;
      17497: inst = 32'h10408000;
      17498: inst = 32'hc4055b4;
      17499: inst = 32'h8220000;
      17500: inst = 32'h10408000;
      17501: inst = 32'hc4055ca;
      17502: inst = 32'h8220000;
      17503: inst = 32'h10408000;
      17504: inst = 32'hc4055cb;
      17505: inst = 32'h8220000;
      17506: inst = 32'h10408000;
      17507: inst = 32'hc4055cc;
      17508: inst = 32'h8220000;
      17509: inst = 32'h10408000;
      17510: inst = 32'hc4055cd;
      17511: inst = 32'h8220000;
      17512: inst = 32'h10408000;
      17513: inst = 32'hc4055ce;
      17514: inst = 32'h8220000;
      17515: inst = 32'h10408000;
      17516: inst = 32'hc4055cf;
      17517: inst = 32'h8220000;
      17518: inst = 32'h10408000;
      17519: inst = 32'hc4055d0;
      17520: inst = 32'h8220000;
      17521: inst = 32'h10408000;
      17522: inst = 32'hc4055d1;
      17523: inst = 32'h8220000;
      17524: inst = 32'h10408000;
      17525: inst = 32'hc4055d2;
      17526: inst = 32'h8220000;
      17527: inst = 32'h10408000;
      17528: inst = 32'hc4055d3;
      17529: inst = 32'h8220000;
      17530: inst = 32'h10408000;
      17531: inst = 32'hc4055d4;
      17532: inst = 32'h8220000;
      17533: inst = 32'h10408000;
      17534: inst = 32'hc4055d5;
      17535: inst = 32'h8220000;
      17536: inst = 32'h10408000;
      17537: inst = 32'hc4055eb;
      17538: inst = 32'h8220000;
      17539: inst = 32'h10408000;
      17540: inst = 32'hc4055ec;
      17541: inst = 32'h8220000;
      17542: inst = 32'h10408000;
      17543: inst = 32'hc4055ed;
      17544: inst = 32'h8220000;
      17545: inst = 32'h10408000;
      17546: inst = 32'hc4055ee;
      17547: inst = 32'h8220000;
      17548: inst = 32'h10408000;
      17549: inst = 32'hc4055ef;
      17550: inst = 32'h8220000;
      17551: inst = 32'h10408000;
      17552: inst = 32'hc4055f0;
      17553: inst = 32'h8220000;
      17554: inst = 32'h10408000;
      17555: inst = 32'hc4055f1;
      17556: inst = 32'h8220000;
      17557: inst = 32'h10408000;
      17558: inst = 32'hc4055f2;
      17559: inst = 32'h8220000;
      17560: inst = 32'h10408000;
      17561: inst = 32'hc4055f3;
      17562: inst = 32'h8220000;
      17563: inst = 32'h10408000;
      17564: inst = 32'hc4055f4;
      17565: inst = 32'h8220000;
      17566: inst = 32'h10408000;
      17567: inst = 32'hc4055f5;
      17568: inst = 32'h8220000;
      17569: inst = 32'h10408000;
      17570: inst = 32'hc4055f6;
      17571: inst = 32'h8220000;
      17572: inst = 32'h10408000;
      17573: inst = 32'hc4055f7;
      17574: inst = 32'h8220000;
      17575: inst = 32'h10408000;
      17576: inst = 32'hc4055f8;
      17577: inst = 32'h8220000;
      17578: inst = 32'h10408000;
      17579: inst = 32'hc4055f9;
      17580: inst = 32'h8220000;
      17581: inst = 32'h10408000;
      17582: inst = 32'hc4055fa;
      17583: inst = 32'h8220000;
      17584: inst = 32'h10408000;
      17585: inst = 32'hc4055fb;
      17586: inst = 32'h8220000;
      17587: inst = 32'h10408000;
      17588: inst = 32'hc4055fc;
      17589: inst = 32'h8220000;
      17590: inst = 32'h10408000;
      17591: inst = 32'hc4055fd;
      17592: inst = 32'h8220000;
      17593: inst = 32'h10408000;
      17594: inst = 32'hc4055fe;
      17595: inst = 32'h8220000;
      17596: inst = 32'h10408000;
      17597: inst = 32'hc4055ff;
      17598: inst = 32'h8220000;
      17599: inst = 32'h10408000;
      17600: inst = 32'hc405600;
      17601: inst = 32'h8220000;
      17602: inst = 32'h10408000;
      17603: inst = 32'hc405601;
      17604: inst = 32'h8220000;
      17605: inst = 32'h10408000;
      17606: inst = 32'hc405602;
      17607: inst = 32'h8220000;
      17608: inst = 32'h10408000;
      17609: inst = 32'hc405603;
      17610: inst = 32'h8220000;
      17611: inst = 32'h10408000;
      17612: inst = 32'hc405604;
      17613: inst = 32'h8220000;
      17614: inst = 32'h10408000;
      17615: inst = 32'hc405605;
      17616: inst = 32'h8220000;
      17617: inst = 32'h10408000;
      17618: inst = 32'hc405606;
      17619: inst = 32'h8220000;
      17620: inst = 32'h10408000;
      17621: inst = 32'hc405607;
      17622: inst = 32'h8220000;
      17623: inst = 32'h10408000;
      17624: inst = 32'hc405608;
      17625: inst = 32'h8220000;
      17626: inst = 32'h10408000;
      17627: inst = 32'hc405609;
      17628: inst = 32'h8220000;
      17629: inst = 32'h10408000;
      17630: inst = 32'hc40560a;
      17631: inst = 32'h8220000;
      17632: inst = 32'h10408000;
      17633: inst = 32'hc40560b;
      17634: inst = 32'h8220000;
      17635: inst = 32'h10408000;
      17636: inst = 32'hc40560c;
      17637: inst = 32'h8220000;
      17638: inst = 32'h10408000;
      17639: inst = 32'hc40560d;
      17640: inst = 32'h8220000;
      17641: inst = 32'h10408000;
      17642: inst = 32'hc40560e;
      17643: inst = 32'h8220000;
      17644: inst = 32'h10408000;
      17645: inst = 32'hc40560f;
      17646: inst = 32'h8220000;
      17647: inst = 32'h10408000;
      17648: inst = 32'hc405610;
      17649: inst = 32'h8220000;
      17650: inst = 32'h10408000;
      17651: inst = 32'hc405611;
      17652: inst = 32'h8220000;
      17653: inst = 32'h10408000;
      17654: inst = 32'hc405612;
      17655: inst = 32'h8220000;
      17656: inst = 32'h10408000;
      17657: inst = 32'hc405613;
      17658: inst = 32'h8220000;
      17659: inst = 32'h10408000;
      17660: inst = 32'hc405614;
      17661: inst = 32'h8220000;
      17662: inst = 32'h10408000;
      17663: inst = 32'hc40562a;
      17664: inst = 32'h8220000;
      17665: inst = 32'h10408000;
      17666: inst = 32'hc40562b;
      17667: inst = 32'h8220000;
      17668: inst = 32'h10408000;
      17669: inst = 32'hc40562c;
      17670: inst = 32'h8220000;
      17671: inst = 32'h10408000;
      17672: inst = 32'hc40562d;
      17673: inst = 32'h8220000;
      17674: inst = 32'h10408000;
      17675: inst = 32'hc40562e;
      17676: inst = 32'h8220000;
      17677: inst = 32'h10408000;
      17678: inst = 32'hc40562f;
      17679: inst = 32'h8220000;
      17680: inst = 32'h10408000;
      17681: inst = 32'hc405630;
      17682: inst = 32'h8220000;
      17683: inst = 32'h10408000;
      17684: inst = 32'hc405631;
      17685: inst = 32'h8220000;
      17686: inst = 32'h10408000;
      17687: inst = 32'hc405632;
      17688: inst = 32'h8220000;
      17689: inst = 32'h10408000;
      17690: inst = 32'hc405633;
      17691: inst = 32'h8220000;
      17692: inst = 32'h10408000;
      17693: inst = 32'hc405634;
      17694: inst = 32'h8220000;
      17695: inst = 32'h10408000;
      17696: inst = 32'hc405635;
      17697: inst = 32'h8220000;
      17698: inst = 32'h10408000;
      17699: inst = 32'hc40564b;
      17700: inst = 32'h8220000;
      17701: inst = 32'h10408000;
      17702: inst = 32'hc40564c;
      17703: inst = 32'h8220000;
      17704: inst = 32'h10408000;
      17705: inst = 32'hc40564d;
      17706: inst = 32'h8220000;
      17707: inst = 32'h10408000;
      17708: inst = 32'hc40564e;
      17709: inst = 32'h8220000;
      17710: inst = 32'h10408000;
      17711: inst = 32'hc40564f;
      17712: inst = 32'h8220000;
      17713: inst = 32'h10408000;
      17714: inst = 32'hc405650;
      17715: inst = 32'h8220000;
      17716: inst = 32'h10408000;
      17717: inst = 32'hc405651;
      17718: inst = 32'h8220000;
      17719: inst = 32'h10408000;
      17720: inst = 32'hc405652;
      17721: inst = 32'h8220000;
      17722: inst = 32'h10408000;
      17723: inst = 32'hc405653;
      17724: inst = 32'h8220000;
      17725: inst = 32'h10408000;
      17726: inst = 32'hc405654;
      17727: inst = 32'h8220000;
      17728: inst = 32'h10408000;
      17729: inst = 32'hc405655;
      17730: inst = 32'h8220000;
      17731: inst = 32'h10408000;
      17732: inst = 32'hc405656;
      17733: inst = 32'h8220000;
      17734: inst = 32'h10408000;
      17735: inst = 32'hc405657;
      17736: inst = 32'h8220000;
      17737: inst = 32'h10408000;
      17738: inst = 32'hc405658;
      17739: inst = 32'h8220000;
      17740: inst = 32'h10408000;
      17741: inst = 32'hc405659;
      17742: inst = 32'h8220000;
      17743: inst = 32'h10408000;
      17744: inst = 32'hc40565a;
      17745: inst = 32'h8220000;
      17746: inst = 32'h10408000;
      17747: inst = 32'hc40565b;
      17748: inst = 32'h8220000;
      17749: inst = 32'h10408000;
      17750: inst = 32'hc40565c;
      17751: inst = 32'h8220000;
      17752: inst = 32'h10408000;
      17753: inst = 32'hc40565d;
      17754: inst = 32'h8220000;
      17755: inst = 32'h10408000;
      17756: inst = 32'hc40565e;
      17757: inst = 32'h8220000;
      17758: inst = 32'h10408000;
      17759: inst = 32'hc40565f;
      17760: inst = 32'h8220000;
      17761: inst = 32'h10408000;
      17762: inst = 32'hc405660;
      17763: inst = 32'h8220000;
      17764: inst = 32'h10408000;
      17765: inst = 32'hc405661;
      17766: inst = 32'h8220000;
      17767: inst = 32'h10408000;
      17768: inst = 32'hc405662;
      17769: inst = 32'h8220000;
      17770: inst = 32'h10408000;
      17771: inst = 32'hc405663;
      17772: inst = 32'h8220000;
      17773: inst = 32'h10408000;
      17774: inst = 32'hc405664;
      17775: inst = 32'h8220000;
      17776: inst = 32'h10408000;
      17777: inst = 32'hc405665;
      17778: inst = 32'h8220000;
      17779: inst = 32'h10408000;
      17780: inst = 32'hc405666;
      17781: inst = 32'h8220000;
      17782: inst = 32'h10408000;
      17783: inst = 32'hc405667;
      17784: inst = 32'h8220000;
      17785: inst = 32'h10408000;
      17786: inst = 32'hc405668;
      17787: inst = 32'h8220000;
      17788: inst = 32'h10408000;
      17789: inst = 32'hc405669;
      17790: inst = 32'h8220000;
      17791: inst = 32'h10408000;
      17792: inst = 32'hc40566a;
      17793: inst = 32'h8220000;
      17794: inst = 32'h10408000;
      17795: inst = 32'hc40566b;
      17796: inst = 32'h8220000;
      17797: inst = 32'h10408000;
      17798: inst = 32'hc40566c;
      17799: inst = 32'h8220000;
      17800: inst = 32'h10408000;
      17801: inst = 32'hc40566d;
      17802: inst = 32'h8220000;
      17803: inst = 32'h10408000;
      17804: inst = 32'hc40566e;
      17805: inst = 32'h8220000;
      17806: inst = 32'h10408000;
      17807: inst = 32'hc40566f;
      17808: inst = 32'h8220000;
      17809: inst = 32'h10408000;
      17810: inst = 32'hc405670;
      17811: inst = 32'h8220000;
      17812: inst = 32'h10408000;
      17813: inst = 32'hc405671;
      17814: inst = 32'h8220000;
      17815: inst = 32'h10408000;
      17816: inst = 32'hc405672;
      17817: inst = 32'h8220000;
      17818: inst = 32'h10408000;
      17819: inst = 32'hc405673;
      17820: inst = 32'h8220000;
      17821: inst = 32'h10408000;
      17822: inst = 32'hc40568a;
      17823: inst = 32'h8220000;
      17824: inst = 32'h10408000;
      17825: inst = 32'hc40568b;
      17826: inst = 32'h8220000;
      17827: inst = 32'h10408000;
      17828: inst = 32'hc40568c;
      17829: inst = 32'h8220000;
      17830: inst = 32'h10408000;
      17831: inst = 32'hc40568d;
      17832: inst = 32'h8220000;
      17833: inst = 32'h10408000;
      17834: inst = 32'hc40568e;
      17835: inst = 32'h8220000;
      17836: inst = 32'h10408000;
      17837: inst = 32'hc40568f;
      17838: inst = 32'h8220000;
      17839: inst = 32'h10408000;
      17840: inst = 32'hc405690;
      17841: inst = 32'h8220000;
      17842: inst = 32'h10408000;
      17843: inst = 32'hc405691;
      17844: inst = 32'h8220000;
      17845: inst = 32'h10408000;
      17846: inst = 32'hc405692;
      17847: inst = 32'h8220000;
      17848: inst = 32'h10408000;
      17849: inst = 32'hc405693;
      17850: inst = 32'h8220000;
      17851: inst = 32'h10408000;
      17852: inst = 32'hc405694;
      17853: inst = 32'h8220000;
      17854: inst = 32'h10408000;
      17855: inst = 32'hc405695;
      17856: inst = 32'h8220000;
      17857: inst = 32'h10408000;
      17858: inst = 32'hc4056ac;
      17859: inst = 32'h8220000;
      17860: inst = 32'h10408000;
      17861: inst = 32'hc4056ad;
      17862: inst = 32'h8220000;
      17863: inst = 32'h10408000;
      17864: inst = 32'hc4056ae;
      17865: inst = 32'h8220000;
      17866: inst = 32'h10408000;
      17867: inst = 32'hc4056af;
      17868: inst = 32'h8220000;
      17869: inst = 32'h10408000;
      17870: inst = 32'hc4056b0;
      17871: inst = 32'h8220000;
      17872: inst = 32'h10408000;
      17873: inst = 32'hc4056b1;
      17874: inst = 32'h8220000;
      17875: inst = 32'h10408000;
      17876: inst = 32'hc4056b2;
      17877: inst = 32'h8220000;
      17878: inst = 32'h10408000;
      17879: inst = 32'hc4056b3;
      17880: inst = 32'h8220000;
      17881: inst = 32'h10408000;
      17882: inst = 32'hc4056b4;
      17883: inst = 32'h8220000;
      17884: inst = 32'h10408000;
      17885: inst = 32'hc4056b5;
      17886: inst = 32'h8220000;
      17887: inst = 32'h10408000;
      17888: inst = 32'hc4056b6;
      17889: inst = 32'h8220000;
      17890: inst = 32'h10408000;
      17891: inst = 32'hc4056b7;
      17892: inst = 32'h8220000;
      17893: inst = 32'h10408000;
      17894: inst = 32'hc4056b8;
      17895: inst = 32'h8220000;
      17896: inst = 32'h10408000;
      17897: inst = 32'hc4056b9;
      17898: inst = 32'h8220000;
      17899: inst = 32'h10408000;
      17900: inst = 32'hc4056ba;
      17901: inst = 32'h8220000;
      17902: inst = 32'h10408000;
      17903: inst = 32'hc4056bb;
      17904: inst = 32'h8220000;
      17905: inst = 32'h10408000;
      17906: inst = 32'hc4056bc;
      17907: inst = 32'h8220000;
      17908: inst = 32'h10408000;
      17909: inst = 32'hc4056bd;
      17910: inst = 32'h8220000;
      17911: inst = 32'h10408000;
      17912: inst = 32'hc4056be;
      17913: inst = 32'h8220000;
      17914: inst = 32'h10408000;
      17915: inst = 32'hc4056bf;
      17916: inst = 32'h8220000;
      17917: inst = 32'h10408000;
      17918: inst = 32'hc4056c0;
      17919: inst = 32'h8220000;
      17920: inst = 32'h10408000;
      17921: inst = 32'hc4056c1;
      17922: inst = 32'h8220000;
      17923: inst = 32'h10408000;
      17924: inst = 32'hc4056c2;
      17925: inst = 32'h8220000;
      17926: inst = 32'h10408000;
      17927: inst = 32'hc4056c3;
      17928: inst = 32'h8220000;
      17929: inst = 32'h10408000;
      17930: inst = 32'hc4056c4;
      17931: inst = 32'h8220000;
      17932: inst = 32'h10408000;
      17933: inst = 32'hc4056c5;
      17934: inst = 32'h8220000;
      17935: inst = 32'h10408000;
      17936: inst = 32'hc4056c6;
      17937: inst = 32'h8220000;
      17938: inst = 32'h10408000;
      17939: inst = 32'hc4056c7;
      17940: inst = 32'h8220000;
      17941: inst = 32'h10408000;
      17942: inst = 32'hc4056c8;
      17943: inst = 32'h8220000;
      17944: inst = 32'h10408000;
      17945: inst = 32'hc4056c9;
      17946: inst = 32'h8220000;
      17947: inst = 32'h10408000;
      17948: inst = 32'hc4056ca;
      17949: inst = 32'h8220000;
      17950: inst = 32'h10408000;
      17951: inst = 32'hc4056cb;
      17952: inst = 32'h8220000;
      17953: inst = 32'h10408000;
      17954: inst = 32'hc4056cc;
      17955: inst = 32'h8220000;
      17956: inst = 32'h10408000;
      17957: inst = 32'hc4056cd;
      17958: inst = 32'h8220000;
      17959: inst = 32'h10408000;
      17960: inst = 32'hc4056ce;
      17961: inst = 32'h8220000;
      17962: inst = 32'h10408000;
      17963: inst = 32'hc4056cf;
      17964: inst = 32'h8220000;
      17965: inst = 32'h10408000;
      17966: inst = 32'hc4056d0;
      17967: inst = 32'h8220000;
      17968: inst = 32'h10408000;
      17969: inst = 32'hc4056d1;
      17970: inst = 32'h8220000;
      17971: inst = 32'h10408000;
      17972: inst = 32'hc4056d2;
      17973: inst = 32'h8220000;
      17974: inst = 32'h10408000;
      17975: inst = 32'hc4056ea;
      17976: inst = 32'h8220000;
      17977: inst = 32'h10408000;
      17978: inst = 32'hc4056eb;
      17979: inst = 32'h8220000;
      17980: inst = 32'h10408000;
      17981: inst = 32'hc4056ec;
      17982: inst = 32'h8220000;
      17983: inst = 32'h10408000;
      17984: inst = 32'hc4056ed;
      17985: inst = 32'h8220000;
      17986: inst = 32'h10408000;
      17987: inst = 32'hc4056ee;
      17988: inst = 32'h8220000;
      17989: inst = 32'h10408000;
      17990: inst = 32'hc4056ef;
      17991: inst = 32'h8220000;
      17992: inst = 32'h10408000;
      17993: inst = 32'hc4056f0;
      17994: inst = 32'h8220000;
      17995: inst = 32'h10408000;
      17996: inst = 32'hc4056f1;
      17997: inst = 32'h8220000;
      17998: inst = 32'h10408000;
      17999: inst = 32'hc4056f2;
      18000: inst = 32'h8220000;
      18001: inst = 32'h10408000;
      18002: inst = 32'hc4056f3;
      18003: inst = 32'h8220000;
      18004: inst = 32'h10408000;
      18005: inst = 32'hc4056f4;
      18006: inst = 32'h8220000;
      18007: inst = 32'h10408000;
      18008: inst = 32'hc4056f5;
      18009: inst = 32'h8220000;
      18010: inst = 32'h10408000;
      18011: inst = 32'hc40570d;
      18012: inst = 32'h8220000;
      18013: inst = 32'h10408000;
      18014: inst = 32'hc40570e;
      18015: inst = 32'h8220000;
      18016: inst = 32'h10408000;
      18017: inst = 32'hc40570f;
      18018: inst = 32'h8220000;
      18019: inst = 32'h10408000;
      18020: inst = 32'hc405710;
      18021: inst = 32'h8220000;
      18022: inst = 32'h10408000;
      18023: inst = 32'hc405711;
      18024: inst = 32'h8220000;
      18025: inst = 32'h10408000;
      18026: inst = 32'hc405712;
      18027: inst = 32'h8220000;
      18028: inst = 32'h10408000;
      18029: inst = 32'hc405713;
      18030: inst = 32'h8220000;
      18031: inst = 32'h10408000;
      18032: inst = 32'hc405714;
      18033: inst = 32'h8220000;
      18034: inst = 32'h10408000;
      18035: inst = 32'hc405715;
      18036: inst = 32'h8220000;
      18037: inst = 32'h10408000;
      18038: inst = 32'hc405716;
      18039: inst = 32'h8220000;
      18040: inst = 32'h10408000;
      18041: inst = 32'hc405717;
      18042: inst = 32'h8220000;
      18043: inst = 32'h10408000;
      18044: inst = 32'hc405718;
      18045: inst = 32'h8220000;
      18046: inst = 32'h10408000;
      18047: inst = 32'hc405719;
      18048: inst = 32'h8220000;
      18049: inst = 32'h10408000;
      18050: inst = 32'hc40571a;
      18051: inst = 32'h8220000;
      18052: inst = 32'h10408000;
      18053: inst = 32'hc40571b;
      18054: inst = 32'h8220000;
      18055: inst = 32'h10408000;
      18056: inst = 32'hc40571c;
      18057: inst = 32'h8220000;
      18058: inst = 32'h10408000;
      18059: inst = 32'hc40571d;
      18060: inst = 32'h8220000;
      18061: inst = 32'h10408000;
      18062: inst = 32'hc40571e;
      18063: inst = 32'h8220000;
      18064: inst = 32'h10408000;
      18065: inst = 32'hc40571f;
      18066: inst = 32'h8220000;
      18067: inst = 32'h10408000;
      18068: inst = 32'hc405720;
      18069: inst = 32'h8220000;
      18070: inst = 32'h10408000;
      18071: inst = 32'hc405721;
      18072: inst = 32'h8220000;
      18073: inst = 32'h10408000;
      18074: inst = 32'hc405722;
      18075: inst = 32'h8220000;
      18076: inst = 32'h10408000;
      18077: inst = 32'hc405723;
      18078: inst = 32'h8220000;
      18079: inst = 32'h10408000;
      18080: inst = 32'hc405724;
      18081: inst = 32'h8220000;
      18082: inst = 32'h10408000;
      18083: inst = 32'hc405725;
      18084: inst = 32'h8220000;
      18085: inst = 32'h10408000;
      18086: inst = 32'hc405726;
      18087: inst = 32'h8220000;
      18088: inst = 32'h10408000;
      18089: inst = 32'hc405727;
      18090: inst = 32'h8220000;
      18091: inst = 32'h10408000;
      18092: inst = 32'hc405728;
      18093: inst = 32'h8220000;
      18094: inst = 32'h10408000;
      18095: inst = 32'hc405729;
      18096: inst = 32'h8220000;
      18097: inst = 32'h10408000;
      18098: inst = 32'hc40572a;
      18099: inst = 32'h8220000;
      18100: inst = 32'h10408000;
      18101: inst = 32'hc40572b;
      18102: inst = 32'h8220000;
      18103: inst = 32'h10408000;
      18104: inst = 32'hc40572c;
      18105: inst = 32'h8220000;
      18106: inst = 32'h10408000;
      18107: inst = 32'hc40572d;
      18108: inst = 32'h8220000;
      18109: inst = 32'h10408000;
      18110: inst = 32'hc40572e;
      18111: inst = 32'h8220000;
      18112: inst = 32'h10408000;
      18113: inst = 32'hc40572f;
      18114: inst = 32'h8220000;
      18115: inst = 32'h10408000;
      18116: inst = 32'hc405730;
      18117: inst = 32'h8220000;
      18118: inst = 32'h10408000;
      18119: inst = 32'hc405731;
      18120: inst = 32'h8220000;
      18121: inst = 32'h10408000;
      18122: inst = 32'hc40574a;
      18123: inst = 32'h8220000;
      18124: inst = 32'h10408000;
      18125: inst = 32'hc40574b;
      18126: inst = 32'h8220000;
      18127: inst = 32'h10408000;
      18128: inst = 32'hc40574c;
      18129: inst = 32'h8220000;
      18130: inst = 32'h10408000;
      18131: inst = 32'hc40574d;
      18132: inst = 32'h8220000;
      18133: inst = 32'h10408000;
      18134: inst = 32'hc40574e;
      18135: inst = 32'h8220000;
      18136: inst = 32'h10408000;
      18137: inst = 32'hc40574f;
      18138: inst = 32'h8220000;
      18139: inst = 32'h10408000;
      18140: inst = 32'hc405750;
      18141: inst = 32'h8220000;
      18142: inst = 32'h10408000;
      18143: inst = 32'hc405751;
      18144: inst = 32'h8220000;
      18145: inst = 32'h10408000;
      18146: inst = 32'hc405752;
      18147: inst = 32'h8220000;
      18148: inst = 32'h10408000;
      18149: inst = 32'hc405753;
      18150: inst = 32'h8220000;
      18151: inst = 32'h10408000;
      18152: inst = 32'hc405754;
      18153: inst = 32'h8220000;
      18154: inst = 32'h10408000;
      18155: inst = 32'hc405755;
      18156: inst = 32'h8220000;
      18157: inst = 32'h10408000;
      18158: inst = 32'hc40576e;
      18159: inst = 32'h8220000;
      18160: inst = 32'h10408000;
      18161: inst = 32'hc40576f;
      18162: inst = 32'h8220000;
      18163: inst = 32'h10408000;
      18164: inst = 32'hc405770;
      18165: inst = 32'h8220000;
      18166: inst = 32'h10408000;
      18167: inst = 32'hc405771;
      18168: inst = 32'h8220000;
      18169: inst = 32'h10408000;
      18170: inst = 32'hc405772;
      18171: inst = 32'h8220000;
      18172: inst = 32'h10408000;
      18173: inst = 32'hc405773;
      18174: inst = 32'h8220000;
      18175: inst = 32'h10408000;
      18176: inst = 32'hc405774;
      18177: inst = 32'h8220000;
      18178: inst = 32'h10408000;
      18179: inst = 32'hc405775;
      18180: inst = 32'h8220000;
      18181: inst = 32'h10408000;
      18182: inst = 32'hc405776;
      18183: inst = 32'h8220000;
      18184: inst = 32'h10408000;
      18185: inst = 32'hc405777;
      18186: inst = 32'h8220000;
      18187: inst = 32'h10408000;
      18188: inst = 32'hc405778;
      18189: inst = 32'h8220000;
      18190: inst = 32'h10408000;
      18191: inst = 32'hc405779;
      18192: inst = 32'h8220000;
      18193: inst = 32'h10408000;
      18194: inst = 32'hc40577a;
      18195: inst = 32'h8220000;
      18196: inst = 32'h10408000;
      18197: inst = 32'hc40577b;
      18198: inst = 32'h8220000;
      18199: inst = 32'h10408000;
      18200: inst = 32'hc40577c;
      18201: inst = 32'h8220000;
      18202: inst = 32'h10408000;
      18203: inst = 32'hc40577d;
      18204: inst = 32'h8220000;
      18205: inst = 32'h10408000;
      18206: inst = 32'hc40577e;
      18207: inst = 32'h8220000;
      18208: inst = 32'h10408000;
      18209: inst = 32'hc40577f;
      18210: inst = 32'h8220000;
      18211: inst = 32'h10408000;
      18212: inst = 32'hc405780;
      18213: inst = 32'h8220000;
      18214: inst = 32'h10408000;
      18215: inst = 32'hc405781;
      18216: inst = 32'h8220000;
      18217: inst = 32'h10408000;
      18218: inst = 32'hc405782;
      18219: inst = 32'h8220000;
      18220: inst = 32'h10408000;
      18221: inst = 32'hc405783;
      18222: inst = 32'h8220000;
      18223: inst = 32'h10408000;
      18224: inst = 32'hc405784;
      18225: inst = 32'h8220000;
      18226: inst = 32'h10408000;
      18227: inst = 32'hc405785;
      18228: inst = 32'h8220000;
      18229: inst = 32'h10408000;
      18230: inst = 32'hc405786;
      18231: inst = 32'h8220000;
      18232: inst = 32'h10408000;
      18233: inst = 32'hc405787;
      18234: inst = 32'h8220000;
      18235: inst = 32'h10408000;
      18236: inst = 32'hc405788;
      18237: inst = 32'h8220000;
      18238: inst = 32'h10408000;
      18239: inst = 32'hc405789;
      18240: inst = 32'h8220000;
      18241: inst = 32'h10408000;
      18242: inst = 32'hc40578a;
      18243: inst = 32'h8220000;
      18244: inst = 32'h10408000;
      18245: inst = 32'hc40578b;
      18246: inst = 32'h8220000;
      18247: inst = 32'h10408000;
      18248: inst = 32'hc40578c;
      18249: inst = 32'h8220000;
      18250: inst = 32'h10408000;
      18251: inst = 32'hc40578d;
      18252: inst = 32'h8220000;
      18253: inst = 32'h10408000;
      18254: inst = 32'hc40578e;
      18255: inst = 32'h8220000;
      18256: inst = 32'h10408000;
      18257: inst = 32'hc40578f;
      18258: inst = 32'h8220000;
      18259: inst = 32'h10408000;
      18260: inst = 32'hc405790;
      18261: inst = 32'h8220000;
      18262: inst = 32'h10408000;
      18263: inst = 32'hc405791;
      18264: inst = 32'h8220000;
      18265: inst = 32'h10408000;
      18266: inst = 32'hc4057aa;
      18267: inst = 32'h8220000;
      18268: inst = 32'h10408000;
      18269: inst = 32'hc4057ab;
      18270: inst = 32'h8220000;
      18271: inst = 32'h10408000;
      18272: inst = 32'hc4057ac;
      18273: inst = 32'h8220000;
      18274: inst = 32'h10408000;
      18275: inst = 32'hc4057ad;
      18276: inst = 32'h8220000;
      18277: inst = 32'h10408000;
      18278: inst = 32'hc4057ae;
      18279: inst = 32'h8220000;
      18280: inst = 32'h10408000;
      18281: inst = 32'hc4057af;
      18282: inst = 32'h8220000;
      18283: inst = 32'h10408000;
      18284: inst = 32'hc4057b0;
      18285: inst = 32'h8220000;
      18286: inst = 32'h10408000;
      18287: inst = 32'hc4057b1;
      18288: inst = 32'h8220000;
      18289: inst = 32'h10408000;
      18290: inst = 32'hc4057b2;
      18291: inst = 32'h8220000;
      18292: inst = 32'h10408000;
      18293: inst = 32'hc4057b3;
      18294: inst = 32'h8220000;
      18295: inst = 32'h10408000;
      18296: inst = 32'hc4057b4;
      18297: inst = 32'h8220000;
      18298: inst = 32'h10408000;
      18299: inst = 32'hc4057b5;
      18300: inst = 32'h8220000;
      18301: inst = 32'h10408000;
      18302: inst = 32'hc4057ce;
      18303: inst = 32'h8220000;
      18304: inst = 32'h10408000;
      18305: inst = 32'hc4057cf;
      18306: inst = 32'h8220000;
      18307: inst = 32'h10408000;
      18308: inst = 32'hc4057d0;
      18309: inst = 32'h8220000;
      18310: inst = 32'h10408000;
      18311: inst = 32'hc4057d1;
      18312: inst = 32'h8220000;
      18313: inst = 32'h10408000;
      18314: inst = 32'hc4057d2;
      18315: inst = 32'h8220000;
      18316: inst = 32'h10408000;
      18317: inst = 32'hc4057d3;
      18318: inst = 32'h8220000;
      18319: inst = 32'h10408000;
      18320: inst = 32'hc4057d4;
      18321: inst = 32'h8220000;
      18322: inst = 32'h10408000;
      18323: inst = 32'hc4057d5;
      18324: inst = 32'h8220000;
      18325: inst = 32'h10408000;
      18326: inst = 32'hc4057d6;
      18327: inst = 32'h8220000;
      18328: inst = 32'h10408000;
      18329: inst = 32'hc4057d7;
      18330: inst = 32'h8220000;
      18331: inst = 32'h10408000;
      18332: inst = 32'hc4057d8;
      18333: inst = 32'h8220000;
      18334: inst = 32'h10408000;
      18335: inst = 32'hc4057d9;
      18336: inst = 32'h8220000;
      18337: inst = 32'h10408000;
      18338: inst = 32'hc4057da;
      18339: inst = 32'h8220000;
      18340: inst = 32'h10408000;
      18341: inst = 32'hc4057db;
      18342: inst = 32'h8220000;
      18343: inst = 32'h10408000;
      18344: inst = 32'hc4057dc;
      18345: inst = 32'h8220000;
      18346: inst = 32'h10408000;
      18347: inst = 32'hc4057dd;
      18348: inst = 32'h8220000;
      18349: inst = 32'h10408000;
      18350: inst = 32'hc4057de;
      18351: inst = 32'h8220000;
      18352: inst = 32'h10408000;
      18353: inst = 32'hc4057df;
      18354: inst = 32'h8220000;
      18355: inst = 32'hc207bd0;
      18356: inst = 32'h10408000;
      18357: inst = 32'hc40531b;
      18358: inst = 32'h8220000;
      18359: inst = 32'h10408000;
      18360: inst = 32'hc405344;
      18361: inst = 32'h8220000;
      18362: inst = 32'hc207bcf;
      18363: inst = 32'h10408000;
      18364: inst = 32'hc405321;
      18365: inst = 32'h8220000;
      18366: inst = 32'h10408000;
      18367: inst = 32'hc40533e;
      18368: inst = 32'h8220000;
      18369: inst = 32'h10408000;
      18370: inst = 32'hc405381;
      18371: inst = 32'h8220000;
      18372: inst = 32'h10408000;
      18373: inst = 32'hc40539e;
      18374: inst = 32'h8220000;
      18375: inst = 32'h10408000;
      18376: inst = 32'hc4053e1;
      18377: inst = 32'h8220000;
      18378: inst = 32'h10408000;
      18379: inst = 32'hc4053fe;
      18380: inst = 32'h8220000;
      18381: inst = 32'h10408000;
      18382: inst = 32'hc405441;
      18383: inst = 32'h8220000;
      18384: inst = 32'h10408000;
      18385: inst = 32'hc405448;
      18386: inst = 32'h8220000;
      18387: inst = 32'h10408000;
      18388: inst = 32'hc405457;
      18389: inst = 32'h8220000;
      18390: inst = 32'h10408000;
      18391: inst = 32'hc40545e;
      18392: inst = 32'h8220000;
      18393: inst = 32'h10408000;
      18394: inst = 32'hc405501;
      18395: inst = 32'h8220000;
      18396: inst = 32'h10408000;
      18397: inst = 32'hc40551e;
      18398: inst = 32'h8220000;
      18399: inst = 32'h10408000;
      18400: inst = 32'hc405561;
      18401: inst = 32'h8220000;
      18402: inst = 32'h10408000;
      18403: inst = 32'hc40557e;
      18404: inst = 32'h8220000;
      18405: inst = 32'h10408000;
      18406: inst = 32'hc4055b9;
      18407: inst = 32'h8220000;
      18408: inst = 32'h10408000;
      18409: inst = 32'hc4055c1;
      18410: inst = 32'h8220000;
      18411: inst = 32'h10408000;
      18412: inst = 32'hc4055de;
      18413: inst = 32'h8220000;
      18414: inst = 32'h10408000;
      18415: inst = 32'hc4055e6;
      18416: inst = 32'h8220000;
      18417: inst = 32'h10408000;
      18418: inst = 32'hc40561e;
      18419: inst = 32'h8220000;
      18420: inst = 32'h10408000;
      18421: inst = 32'hc405621;
      18422: inst = 32'h8220000;
      18423: inst = 32'h10408000;
      18424: inst = 32'hc40563e;
      18425: inst = 32'h8220000;
      18426: inst = 32'h10408000;
      18427: inst = 32'hc405641;
      18428: inst = 32'h8220000;
      18429: inst = 32'h10408000;
      18430: inst = 32'hc405681;
      18431: inst = 32'h8220000;
      18432: inst = 32'h10408000;
      18433: inst = 32'hc405698;
      18434: inst = 32'h8220000;
      18435: inst = 32'h10408000;
      18436: inst = 32'hc40569e;
      18437: inst = 32'h8220000;
      18438: inst = 32'h10408000;
      18439: inst = 32'hc4056e1;
      18440: inst = 32'h8220000;
      18441: inst = 32'h10408000;
      18442: inst = 32'hc4056fe;
      18443: inst = 32'h8220000;
      18444: inst = 32'hc207390;
      18445: inst = 32'h10408000;
      18446: inst = 32'hc40537a;
      18447: inst = 32'h8220000;
      18448: inst = 32'h10408000;
      18449: inst = 32'hc4053a5;
      18450: inst = 32'h8220000;
      18451: inst = 32'hc2052aa;
      18452: inst = 32'h10408000;
      18453: inst = 32'hc405389;
      18454: inst = 32'h8220000;
      18455: inst = 32'h10408000;
      18456: inst = 32'hc405396;
      18457: inst = 32'h8220000;
      18458: inst = 32'h10408000;
      18459: inst = 32'hc4054fb;
      18460: inst = 32'h8220000;
      18461: inst = 32'h10408000;
      18462: inst = 32'hc405503;
      18463: inst = 32'h8220000;
      18464: inst = 32'h10408000;
      18465: inst = 32'hc40551c;
      18466: inst = 32'h8220000;
      18467: inst = 32'h10408000;
      18468: inst = 32'hc405524;
      18469: inst = 32'h8220000;
      18470: inst = 32'h10408000;
      18471: inst = 32'hc4055c8;
      18472: inst = 32'h8220000;
      18473: inst = 32'h10408000;
      18474: inst = 32'hc4055d7;
      18475: inst = 32'h8220000;
      18476: inst = 32'h10408000;
      18477: inst = 32'hc405619;
      18478: inst = 32'h8220000;
      18479: inst = 32'h10408000;
      18480: inst = 32'hc405622;
      18481: inst = 32'h8220000;
      18482: inst = 32'h10408000;
      18483: inst = 32'hc40563d;
      18484: inst = 32'h8220000;
      18485: inst = 32'h10408000;
      18486: inst = 32'hc405646;
      18487: inst = 32'h8220000;
      18488: inst = 32'hc206b70;
      18489: inst = 32'h10408000;
      18490: inst = 32'hc4053d9;
      18491: inst = 32'h8220000;
      18492: inst = 32'h10408000;
      18493: inst = 32'hc405406;
      18494: inst = 32'h8220000;
      18495: inst = 32'h10408000;
      18496: inst = 32'hc405556;
      18497: inst = 32'h8220000;
      18498: inst = 32'h10408000;
      18499: inst = 32'hc405589;
      18500: inst = 32'h8220000;
      18501: inst = 32'h10408000;
      18502: inst = 32'hc4055b5;
      18503: inst = 32'h8220000;
      18504: inst = 32'h10408000;
      18505: inst = 32'hc4055ea;
      18506: inst = 32'h8220000;
      18507: inst = 32'h10408000;
      18508: inst = 32'hc405732;
      18509: inst = 32'h8220000;
      18510: inst = 32'h10408000;
      18511: inst = 32'hc40576d;
      18512: inst = 32'h8220000;
      18513: inst = 32'hc20736e;
      18514: inst = 32'h10408000;
      18515: inst = 32'hc4053e0;
      18516: inst = 32'h8220000;
      18517: inst = 32'h10408000;
      18518: inst = 32'hc4053ff;
      18519: inst = 32'h8220000;
      18520: inst = 32'hc205aaa;
      18521: inst = 32'h10408000;
      18522: inst = 32'hc4053e4;
      18523: inst = 32'h8220000;
      18524: inst = 32'h10408000;
      18525: inst = 32'hc4053fb;
      18526: inst = 32'h8220000;
      18527: inst = 32'hc208431;
      18528: inst = 32'h10408000;
      18529: inst = 32'hc4053e8;
      18530: inst = 32'h8220000;
      18531: inst = 32'h10408000;
      18532: inst = 32'hc4053f7;
      18533: inst = 32'h8220000;
      18534: inst = 32'h10408000;
      18535: inst = 32'hc405439;
      18536: inst = 32'h8220000;
      18537: inst = 32'h10408000;
      18538: inst = 32'hc405466;
      18539: inst = 32'h8220000;
      18540: inst = 32'h10408000;
      18541: inst = 32'hc4055b6;
      18542: inst = 32'h8220000;
      18543: inst = 32'h10408000;
      18544: inst = 32'hc4055e9;
      18545: inst = 32'h8220000;
      18546: inst = 32'h10408000;
      18547: inst = 32'hc405733;
      18548: inst = 32'h8220000;
      18549: inst = 32'h10408000;
      18550: inst = 32'hc40576c;
      18551: inst = 32'h8220000;
      18552: inst = 32'hc206b4d;
      18553: inst = 32'h10408000;
      18554: inst = 32'hc40543c;
      18555: inst = 32'h8220000;
      18556: inst = 32'h10408000;
      18557: inst = 32'hc405444;
      18558: inst = 32'h8220000;
      18559: inst = 32'h10408000;
      18560: inst = 32'hc40545b;
      18561: inst = 32'h8220000;
      18562: inst = 32'h10408000;
      18563: inst = 32'hc405463;
      18564: inst = 32'h8220000;
      18565: inst = 32'h10408000;
      18566: inst = 32'hc405563;
      18567: inst = 32'h8220000;
      18568: inst = 32'h10408000;
      18569: inst = 32'hc40557c;
      18570: inst = 32'h8220000;
      18571: inst = 32'h10408000;
      18572: inst = 32'hc405682;
      18573: inst = 32'h8220000;
      18574: inst = 32'h10408000;
      18575: inst = 32'hc40569d;
      18576: inst = 32'h8220000;
      18577: inst = 32'hc208430;
      18578: inst = 32'h10408000;
      18579: inst = 32'hc405440;
      18580: inst = 32'h8220000;
      18581: inst = 32'h10408000;
      18582: inst = 32'hc40545f;
      18583: inst = 32'h8220000;
      18584: inst = 32'hc207bf1;
      18585: inst = 32'h10408000;
      18586: inst = 32'hc405498;
      18587: inst = 32'h8220000;
      18588: inst = 32'h10408000;
      18589: inst = 32'hc4054c7;
      18590: inst = 32'h8220000;
      18591: inst = 32'h10408000;
      18592: inst = 32'hc405615;
      18593: inst = 32'h8220000;
      18594: inst = 32'h10408000;
      18595: inst = 32'hc40564a;
      18596: inst = 32'h8220000;
      18597: inst = 32'hc207bef;
      18598: inst = 32'h10408000;
      18599: inst = 32'hc40549b;
      18600: inst = 32'h8220000;
      18601: inst = 32'h10408000;
      18602: inst = 32'hc4054c4;
      18603: inst = 32'h8220000;
      18604: inst = 32'h10408000;
      18605: inst = 32'hc405687;
      18606: inst = 32'h8220000;
      18607: inst = 32'h10408000;
      18608: inst = 32'hc4056e2;
      18609: inst = 32'h8220000;
      18610: inst = 32'h10408000;
      18611: inst = 32'hc4056fd;
      18612: inst = 32'h8220000;
      18613: inst = 32'hc205aeb;
      18614: inst = 32'h10408000;
      18615: inst = 32'hc40549f;
      18616: inst = 32'h8220000;
      18617: inst = 32'h10408000;
      18618: inst = 32'hc4054c0;
      18619: inst = 32'h8220000;
      18620: inst = 32'hc206b6e;
      18621: inst = 32'h10408000;
      18622: inst = 32'hc4054a8;
      18623: inst = 32'h8220000;
      18624: inst = 32'h10408000;
      18625: inst = 32'hc4054b7;
      18626: inst = 32'h8220000;
      18627: inst = 32'h10408000;
      18628: inst = 32'hc4056e7;
      18629: inst = 32'h8220000;
      18630: inst = 32'h10408000;
      18631: inst = 32'hc4056f8;
      18632: inst = 32'h8220000;
      18633: inst = 32'hc2073b0;
      18634: inst = 32'h10408000;
      18635: inst = 32'hc4054f7;
      18636: inst = 32'h8220000;
      18637: inst = 32'h10408000;
      18638: inst = 32'hc405528;
      18639: inst = 32'h8220000;
      18640: inst = 32'h10408000;
      18641: inst = 32'hc405674;
      18642: inst = 32'h8220000;
      18643: inst = 32'h10408000;
      18644: inst = 32'hc4056ab;
      18645: inst = 32'h8220000;
      18646: inst = 32'hc2073ae;
      18647: inst = 32'h10408000;
      18648: inst = 32'hc4054ff;
      18649: inst = 32'h8220000;
      18650: inst = 32'h10408000;
      18651: inst = 32'hc405520;
      18652: inst = 32'h8220000;
      18653: inst = 32'hc20632d;
      18654: inst = 32'h10408000;
      18655: inst = 32'hc405508;
      18656: inst = 32'h8220000;
      18657: inst = 32'h10408000;
      18658: inst = 32'hc405517;
      18659: inst = 32'h8220000;
      18660: inst = 32'h10408000;
      18661: inst = 32'hc405747;
      18662: inst = 32'h8220000;
      18663: inst = 32'h10408000;
      18664: inst = 32'hc405758;
      18665: inst = 32'h8220000;
      18666: inst = 32'hc206b2d;
      18667: inst = 32'h10408000;
      18668: inst = 32'hc40555a;
      18669: inst = 32'h8220000;
      18670: inst = 32'h10408000;
      18671: inst = 32'hc405585;
      18672: inst = 32'h8220000;
      18673: inst = 32'hc20630c;
      18674: inst = 32'h10408000;
      18675: inst = 32'hc4055be;
      18676: inst = 32'h8220000;
      18677: inst = 32'h10408000;
      18678: inst = 32'hc4055e1;
      18679: inst = 32'h8220000;
      18680: inst = 32'h10408000;
      18681: inst = 32'hc405678;
      18682: inst = 32'h8220000;
      18683: inst = 32'hc20632c;
      18684: inst = 32'h10408000;
      18685: inst = 32'hc4056a7;
      18686: inst = 32'h8220000;
      18687: inst = 32'hc206b90;
      18688: inst = 32'h10408000;
      18689: inst = 32'hc4056d3;
      18690: inst = 32'h8220000;
      18691: inst = 32'h10408000;
      18692: inst = 32'hc40570c;
      18693: inst = 32'h8220000;
      18694: inst = 32'hc207c11;
      18695: inst = 32'h10408000;
      18696: inst = 32'hc405792;
      18697: inst = 32'h8220000;
      18698: inst = 32'h10408000;
      18699: inst = 32'hc4057cd;
      18700: inst = 32'h8220000;
      18701: inst = 32'h58000000;
      18702: inst = 32'hc20ea25;
      18703: inst = 32'h10408000;
      18704: inst = 32'hc40464d;
      18705: inst = 32'h8220000;
      18706: inst = 32'h10408000;
      18707: inst = 32'hc40464e;
      18708: inst = 32'h8220000;
      18709: inst = 32'h10408000;
      18710: inst = 32'hc40464f;
      18711: inst = 32'h8220000;
      18712: inst = 32'h10408000;
      18713: inst = 32'hc404650;
      18714: inst = 32'h8220000;
      18715: inst = 32'h10408000;
      18716: inst = 32'hc404651;
      18717: inst = 32'h8220000;
      18718: inst = 32'h10408000;
      18719: inst = 32'hc404652;
      18720: inst = 32'h8220000;
      18721: inst = 32'h10408000;
      18722: inst = 32'hc404653;
      18723: inst = 32'h8220000;
      18724: inst = 32'h10408000;
      18725: inst = 32'hc404654;
      18726: inst = 32'h8220000;
      18727: inst = 32'h10408000;
      18728: inst = 32'hc404655;
      18729: inst = 32'h8220000;
      18730: inst = 32'h10408000;
      18731: inst = 32'hc404659;
      18732: inst = 32'h8220000;
      18733: inst = 32'h10408000;
      18734: inst = 32'hc40465a;
      18735: inst = 32'h8220000;
      18736: inst = 32'h10408000;
      18737: inst = 32'hc40465b;
      18738: inst = 32'h8220000;
      18739: inst = 32'h10408000;
      18740: inst = 32'hc40465c;
      18741: inst = 32'h8220000;
      18742: inst = 32'h10408000;
      18743: inst = 32'hc40465d;
      18744: inst = 32'h8220000;
      18745: inst = 32'h10408000;
      18746: inst = 32'hc40465e;
      18747: inst = 32'h8220000;
      18748: inst = 32'h10408000;
      18749: inst = 32'hc40465f;
      18750: inst = 32'h8220000;
      18751: inst = 32'h10408000;
      18752: inst = 32'hc404660;
      18753: inst = 32'h8220000;
      18754: inst = 32'h10408000;
      18755: inst = 32'hc404661;
      18756: inst = 32'h8220000;
      18757: inst = 32'h10408000;
      18758: inst = 32'hc404663;
      18759: inst = 32'h8220000;
      18760: inst = 32'h10408000;
      18761: inst = 32'hc404664;
      18762: inst = 32'h8220000;
      18763: inst = 32'h10408000;
      18764: inst = 32'hc404665;
      18765: inst = 32'h8220000;
      18766: inst = 32'h10408000;
      18767: inst = 32'hc404666;
      18768: inst = 32'h8220000;
      18769: inst = 32'h10408000;
      18770: inst = 32'hc404667;
      18771: inst = 32'h8220000;
      18772: inst = 32'h10408000;
      18773: inst = 32'hc404668;
      18774: inst = 32'h8220000;
      18775: inst = 32'h10408000;
      18776: inst = 32'hc404669;
      18777: inst = 32'h8220000;
      18778: inst = 32'h10408000;
      18779: inst = 32'hc40466a;
      18780: inst = 32'h8220000;
      18781: inst = 32'h10408000;
      18782: inst = 32'hc40466b;
      18783: inst = 32'h8220000;
      18784: inst = 32'h10408000;
      18785: inst = 32'hc404671;
      18786: inst = 32'h8220000;
      18787: inst = 32'h10408000;
      18788: inst = 32'hc404672;
      18789: inst = 32'h8220000;
      18790: inst = 32'h10408000;
      18791: inst = 32'hc404673;
      18792: inst = 32'h8220000;
      18793: inst = 32'h10408000;
      18794: inst = 32'hc404674;
      18795: inst = 32'h8220000;
      18796: inst = 32'h10408000;
      18797: inst = 32'hc404675;
      18798: inst = 32'h8220000;
      18799: inst = 32'h10408000;
      18800: inst = 32'hc404676;
      18801: inst = 32'h8220000;
      18802: inst = 32'h10408000;
      18803: inst = 32'hc404677;
      18804: inst = 32'h8220000;
      18805: inst = 32'h10408000;
      18806: inst = 32'hc404678;
      18807: inst = 32'h8220000;
      18808: inst = 32'h10408000;
      18809: inst = 32'hc404679;
      18810: inst = 32'h8220000;
      18811: inst = 32'h10408000;
      18812: inst = 32'hc40467c;
      18813: inst = 32'h8220000;
      18814: inst = 32'h10408000;
      18815: inst = 32'hc40467d;
      18816: inst = 32'h8220000;
      18817: inst = 32'h10408000;
      18818: inst = 32'hc40467e;
      18819: inst = 32'h8220000;
      18820: inst = 32'h10408000;
      18821: inst = 32'hc40467f;
      18822: inst = 32'h8220000;
      18823: inst = 32'h10408000;
      18824: inst = 32'hc404680;
      18825: inst = 32'h8220000;
      18826: inst = 32'h10408000;
      18827: inst = 32'hc404681;
      18828: inst = 32'h8220000;
      18829: inst = 32'h10408000;
      18830: inst = 32'hc404682;
      18831: inst = 32'h8220000;
      18832: inst = 32'h10408000;
      18833: inst = 32'hc404683;
      18834: inst = 32'h8220000;
      18835: inst = 32'h10408000;
      18836: inst = 32'hc404684;
      18837: inst = 32'h8220000;
      18838: inst = 32'h10408000;
      18839: inst = 32'hc404685;
      18840: inst = 32'h8220000;
      18841: inst = 32'h10408000;
      18842: inst = 32'hc40468b;
      18843: inst = 32'h8220000;
      18844: inst = 32'h10408000;
      18845: inst = 32'hc40468c;
      18846: inst = 32'h8220000;
      18847: inst = 32'h10408000;
      18848: inst = 32'hc40468d;
      18849: inst = 32'h8220000;
      18850: inst = 32'h10408000;
      18851: inst = 32'hc40468e;
      18852: inst = 32'h8220000;
      18853: inst = 32'h10408000;
      18854: inst = 32'hc40468f;
      18855: inst = 32'h8220000;
      18856: inst = 32'h10408000;
      18857: inst = 32'hc404690;
      18858: inst = 32'h8220000;
      18859: inst = 32'h10408000;
      18860: inst = 32'hc404691;
      18861: inst = 32'h8220000;
      18862: inst = 32'h10408000;
      18863: inst = 32'hc404692;
      18864: inst = 32'h8220000;
      18865: inst = 32'h10408000;
      18866: inst = 32'hc404693;
      18867: inst = 32'h8220000;
      18868: inst = 32'h10408000;
      18869: inst = 32'hc4046ac;
      18870: inst = 32'h8220000;
      18871: inst = 32'h10408000;
      18872: inst = 32'hc4046ad;
      18873: inst = 32'h8220000;
      18874: inst = 32'h10408000;
      18875: inst = 32'hc4046ae;
      18876: inst = 32'h8220000;
      18877: inst = 32'h10408000;
      18878: inst = 32'hc4046af;
      18879: inst = 32'h8220000;
      18880: inst = 32'h10408000;
      18881: inst = 32'hc4046b0;
      18882: inst = 32'h8220000;
      18883: inst = 32'h10408000;
      18884: inst = 32'hc4046b1;
      18885: inst = 32'h8220000;
      18886: inst = 32'h10408000;
      18887: inst = 32'hc4046b2;
      18888: inst = 32'h8220000;
      18889: inst = 32'h10408000;
      18890: inst = 32'hc4046b3;
      18891: inst = 32'h8220000;
      18892: inst = 32'h10408000;
      18893: inst = 32'hc4046b4;
      18894: inst = 32'h8220000;
      18895: inst = 32'h10408000;
      18896: inst = 32'hc4046b5;
      18897: inst = 32'h8220000;
      18898: inst = 32'h10408000;
      18899: inst = 32'hc4046b8;
      18900: inst = 32'h8220000;
      18901: inst = 32'h10408000;
      18902: inst = 32'hc4046b9;
      18903: inst = 32'h8220000;
      18904: inst = 32'h10408000;
      18905: inst = 32'hc4046ba;
      18906: inst = 32'h8220000;
      18907: inst = 32'h10408000;
      18908: inst = 32'hc4046bb;
      18909: inst = 32'h8220000;
      18910: inst = 32'h10408000;
      18911: inst = 32'hc4046bc;
      18912: inst = 32'h8220000;
      18913: inst = 32'h10408000;
      18914: inst = 32'hc4046bd;
      18915: inst = 32'h8220000;
      18916: inst = 32'h10408000;
      18917: inst = 32'hc4046be;
      18918: inst = 32'h8220000;
      18919: inst = 32'h10408000;
      18920: inst = 32'hc4046bf;
      18921: inst = 32'h8220000;
      18922: inst = 32'h10408000;
      18923: inst = 32'hc4046c0;
      18924: inst = 32'h8220000;
      18925: inst = 32'h10408000;
      18926: inst = 32'hc4046c1;
      18927: inst = 32'h8220000;
      18928: inst = 32'h10408000;
      18929: inst = 32'hc4046c3;
      18930: inst = 32'h8220000;
      18931: inst = 32'h10408000;
      18932: inst = 32'hc4046c4;
      18933: inst = 32'h8220000;
      18934: inst = 32'h10408000;
      18935: inst = 32'hc4046c5;
      18936: inst = 32'h8220000;
      18937: inst = 32'h10408000;
      18938: inst = 32'hc4046c6;
      18939: inst = 32'h8220000;
      18940: inst = 32'h10408000;
      18941: inst = 32'hc4046c7;
      18942: inst = 32'h8220000;
      18943: inst = 32'h10408000;
      18944: inst = 32'hc4046c8;
      18945: inst = 32'h8220000;
      18946: inst = 32'h10408000;
      18947: inst = 32'hc4046c9;
      18948: inst = 32'h8220000;
      18949: inst = 32'h10408000;
      18950: inst = 32'hc4046ca;
      18951: inst = 32'h8220000;
      18952: inst = 32'h10408000;
      18953: inst = 32'hc4046cb;
      18954: inst = 32'h8220000;
      18955: inst = 32'h10408000;
      18956: inst = 32'hc4046d0;
      18957: inst = 32'h8220000;
      18958: inst = 32'h10408000;
      18959: inst = 32'hc4046d1;
      18960: inst = 32'h8220000;
      18961: inst = 32'h10408000;
      18962: inst = 32'hc4046d2;
      18963: inst = 32'h8220000;
      18964: inst = 32'h10408000;
      18965: inst = 32'hc4046d3;
      18966: inst = 32'h8220000;
      18967: inst = 32'h10408000;
      18968: inst = 32'hc4046d4;
      18969: inst = 32'h8220000;
      18970: inst = 32'h10408000;
      18971: inst = 32'hc4046d5;
      18972: inst = 32'h8220000;
      18973: inst = 32'h10408000;
      18974: inst = 32'hc4046d6;
      18975: inst = 32'h8220000;
      18976: inst = 32'h10408000;
      18977: inst = 32'hc4046d7;
      18978: inst = 32'h8220000;
      18979: inst = 32'h10408000;
      18980: inst = 32'hc4046d8;
      18981: inst = 32'h8220000;
      18982: inst = 32'h10408000;
      18983: inst = 32'hc4046da;
      18984: inst = 32'h8220000;
      18985: inst = 32'h10408000;
      18986: inst = 32'hc4046dc;
      18987: inst = 32'h8220000;
      18988: inst = 32'h10408000;
      18989: inst = 32'hc4046dd;
      18990: inst = 32'h8220000;
      18991: inst = 32'h10408000;
      18992: inst = 32'hc4046de;
      18993: inst = 32'h8220000;
      18994: inst = 32'h10408000;
      18995: inst = 32'hc4046df;
      18996: inst = 32'h8220000;
      18997: inst = 32'h10408000;
      18998: inst = 32'hc4046e0;
      18999: inst = 32'h8220000;
      19000: inst = 32'h10408000;
      19001: inst = 32'hc4046e1;
      19002: inst = 32'h8220000;
      19003: inst = 32'h10408000;
      19004: inst = 32'hc4046e2;
      19005: inst = 32'h8220000;
      19006: inst = 32'h10408000;
      19007: inst = 32'hc4046e3;
      19008: inst = 32'h8220000;
      19009: inst = 32'h10408000;
      19010: inst = 32'hc4046e4;
      19011: inst = 32'h8220000;
      19012: inst = 32'h10408000;
      19013: inst = 32'hc4046e5;
      19014: inst = 32'h8220000;
      19015: inst = 32'h10408000;
      19016: inst = 32'hc4046ea;
      19017: inst = 32'h8220000;
      19018: inst = 32'h10408000;
      19019: inst = 32'hc4046eb;
      19020: inst = 32'h8220000;
      19021: inst = 32'h10408000;
      19022: inst = 32'hc4046ec;
      19023: inst = 32'h8220000;
      19024: inst = 32'h10408000;
      19025: inst = 32'hc4046ed;
      19026: inst = 32'h8220000;
      19027: inst = 32'h10408000;
      19028: inst = 32'hc4046ee;
      19029: inst = 32'h8220000;
      19030: inst = 32'h10408000;
      19031: inst = 32'hc4046ef;
      19032: inst = 32'h8220000;
      19033: inst = 32'h10408000;
      19034: inst = 32'hc4046f0;
      19035: inst = 32'h8220000;
      19036: inst = 32'h10408000;
      19037: inst = 32'hc4046f1;
      19038: inst = 32'h8220000;
      19039: inst = 32'h10408000;
      19040: inst = 32'hc4046f2;
      19041: inst = 32'h8220000;
      19042: inst = 32'h10408000;
      19043: inst = 32'hc4046f3;
      19044: inst = 32'h8220000;
      19045: inst = 32'h10408000;
      19046: inst = 32'hc40470b;
      19047: inst = 32'h8220000;
      19048: inst = 32'h10408000;
      19049: inst = 32'hc40470c;
      19050: inst = 32'h8220000;
      19051: inst = 32'h10408000;
      19052: inst = 32'hc40470d;
      19053: inst = 32'h8220000;
      19054: inst = 32'h10408000;
      19055: inst = 32'hc404717;
      19056: inst = 32'h8220000;
      19057: inst = 32'h10408000;
      19058: inst = 32'hc404718;
      19059: inst = 32'h8220000;
      19060: inst = 32'h10408000;
      19061: inst = 32'hc404719;
      19062: inst = 32'h8220000;
      19063: inst = 32'h10408000;
      19064: inst = 32'hc404728;
      19065: inst = 32'h8220000;
      19066: inst = 32'h10408000;
      19067: inst = 32'hc404729;
      19068: inst = 32'h8220000;
      19069: inst = 32'h10408000;
      19070: inst = 32'hc40472a;
      19071: inst = 32'h8220000;
      19072: inst = 32'h10408000;
      19073: inst = 32'hc40472b;
      19074: inst = 32'h8220000;
      19075: inst = 32'h10408000;
      19076: inst = 32'hc404730;
      19077: inst = 32'h8220000;
      19078: inst = 32'h10408000;
      19079: inst = 32'hc404731;
      19080: inst = 32'h8220000;
      19081: inst = 32'h10408000;
      19082: inst = 32'hc404735;
      19083: inst = 32'h8220000;
      19084: inst = 32'h10408000;
      19085: inst = 32'hc404736;
      19086: inst = 32'h8220000;
      19087: inst = 32'h10408000;
      19088: inst = 32'hc404737;
      19089: inst = 32'h8220000;
      19090: inst = 32'h10408000;
      19091: inst = 32'hc404739;
      19092: inst = 32'h8220000;
      19093: inst = 32'h10408000;
      19094: inst = 32'hc40473a;
      19095: inst = 32'h8220000;
      19096: inst = 32'h10408000;
      19097: inst = 32'hc404742;
      19098: inst = 32'h8220000;
      19099: inst = 32'h10408000;
      19100: inst = 32'hc404743;
      19101: inst = 32'h8220000;
      19102: inst = 32'h10408000;
      19103: inst = 32'hc404744;
      19104: inst = 32'h8220000;
      19105: inst = 32'h10408000;
      19106: inst = 32'hc404745;
      19107: inst = 32'h8220000;
      19108: inst = 32'h10408000;
      19109: inst = 32'hc404749;
      19110: inst = 32'h8220000;
      19111: inst = 32'h10408000;
      19112: inst = 32'hc40474a;
      19113: inst = 32'h8220000;
      19114: inst = 32'h10408000;
      19115: inst = 32'hc40474b;
      19116: inst = 32'h8220000;
      19117: inst = 32'h10408000;
      19118: inst = 32'hc40476b;
      19119: inst = 32'h8220000;
      19120: inst = 32'h10408000;
      19121: inst = 32'hc40476c;
      19122: inst = 32'h8220000;
      19123: inst = 32'h10408000;
      19124: inst = 32'hc404777;
      19125: inst = 32'h8220000;
      19126: inst = 32'h10408000;
      19127: inst = 32'hc404778;
      19128: inst = 32'h8220000;
      19129: inst = 32'h10408000;
      19130: inst = 32'hc404788;
      19131: inst = 32'h8220000;
      19132: inst = 32'h10408000;
      19133: inst = 32'hc404789;
      19134: inst = 32'h8220000;
      19135: inst = 32'h10408000;
      19136: inst = 32'hc40478a;
      19137: inst = 32'h8220000;
      19138: inst = 32'h10408000;
      19139: inst = 32'hc404790;
      19140: inst = 32'h8220000;
      19141: inst = 32'h10408000;
      19142: inst = 32'hc404791;
      19143: inst = 32'h8220000;
      19144: inst = 32'h10408000;
      19145: inst = 32'hc404795;
      19146: inst = 32'h8220000;
      19147: inst = 32'h10408000;
      19148: inst = 32'hc404799;
      19149: inst = 32'h8220000;
      19150: inst = 32'h10408000;
      19151: inst = 32'hc40479a;
      19152: inst = 32'h8220000;
      19153: inst = 32'h10408000;
      19154: inst = 32'hc4047a2;
      19155: inst = 32'h8220000;
      19156: inst = 32'h10408000;
      19157: inst = 32'hc4047a3;
      19158: inst = 32'h8220000;
      19159: inst = 32'h10408000;
      19160: inst = 32'hc4047a4;
      19161: inst = 32'h8220000;
      19162: inst = 32'h10408000;
      19163: inst = 32'hc4047a9;
      19164: inst = 32'h8220000;
      19165: inst = 32'h10408000;
      19166: inst = 32'hc4047aa;
      19167: inst = 32'h8220000;
      19168: inst = 32'h10408000;
      19169: inst = 32'hc4047cb;
      19170: inst = 32'h8220000;
      19171: inst = 32'h10408000;
      19172: inst = 32'hc4047cc;
      19173: inst = 32'h8220000;
      19174: inst = 32'h10408000;
      19175: inst = 32'hc4047ce;
      19176: inst = 32'h8220000;
      19177: inst = 32'h10408000;
      19178: inst = 32'hc4047cf;
      19179: inst = 32'h8220000;
      19180: inst = 32'h10408000;
      19181: inst = 32'hc4047d0;
      19182: inst = 32'h8220000;
      19183: inst = 32'h10408000;
      19184: inst = 32'hc4047d1;
      19185: inst = 32'h8220000;
      19186: inst = 32'h10408000;
      19187: inst = 32'hc4047d2;
      19188: inst = 32'h8220000;
      19189: inst = 32'h10408000;
      19190: inst = 32'hc4047d7;
      19191: inst = 32'h8220000;
      19192: inst = 32'h10408000;
      19193: inst = 32'hc4047d8;
      19194: inst = 32'h8220000;
      19195: inst = 32'h10408000;
      19196: inst = 32'hc4047da;
      19197: inst = 32'h8220000;
      19198: inst = 32'h10408000;
      19199: inst = 32'hc4047db;
      19200: inst = 32'h8220000;
      19201: inst = 32'h10408000;
      19202: inst = 32'hc4047dc;
      19203: inst = 32'h8220000;
      19204: inst = 32'h10408000;
      19205: inst = 32'hc4047dd;
      19206: inst = 32'h8220000;
      19207: inst = 32'h10408000;
      19208: inst = 32'hc4047de;
      19209: inst = 32'h8220000;
      19210: inst = 32'h10408000;
      19211: inst = 32'hc4047e7;
      19212: inst = 32'h8220000;
      19213: inst = 32'h10408000;
      19214: inst = 32'hc4047e8;
      19215: inst = 32'h8220000;
      19216: inst = 32'h10408000;
      19217: inst = 32'hc4047e9;
      19218: inst = 32'h8220000;
      19219: inst = 32'h10408000;
      19220: inst = 32'hc4047f0;
      19221: inst = 32'h8220000;
      19222: inst = 32'h10408000;
      19223: inst = 32'hc4047f1;
      19224: inst = 32'h8220000;
      19225: inst = 32'h10408000;
      19226: inst = 32'hc4047f9;
      19227: inst = 32'h8220000;
      19228: inst = 32'h10408000;
      19229: inst = 32'hc4047fa;
      19230: inst = 32'h8220000;
      19231: inst = 32'h10408000;
      19232: inst = 32'hc404800;
      19233: inst = 32'h8220000;
      19234: inst = 32'h10408000;
      19235: inst = 32'hc404801;
      19236: inst = 32'h8220000;
      19237: inst = 32'h10408000;
      19238: inst = 32'hc404802;
      19239: inst = 32'h8220000;
      19240: inst = 32'h10408000;
      19241: inst = 32'hc404803;
      19242: inst = 32'h8220000;
      19243: inst = 32'h10408000;
      19244: inst = 32'hc404809;
      19245: inst = 32'h8220000;
      19246: inst = 32'h10408000;
      19247: inst = 32'hc40480a;
      19248: inst = 32'h8220000;
      19249: inst = 32'h10408000;
      19250: inst = 32'hc40480c;
      19251: inst = 32'h8220000;
      19252: inst = 32'h10408000;
      19253: inst = 32'hc40480d;
      19254: inst = 32'h8220000;
      19255: inst = 32'h10408000;
      19256: inst = 32'hc40480e;
      19257: inst = 32'h8220000;
      19258: inst = 32'h10408000;
      19259: inst = 32'hc40480f;
      19260: inst = 32'h8220000;
      19261: inst = 32'h10408000;
      19262: inst = 32'hc404810;
      19263: inst = 32'h8220000;
      19264: inst = 32'h10408000;
      19265: inst = 32'hc404811;
      19266: inst = 32'h8220000;
      19267: inst = 32'h10408000;
      19268: inst = 32'hc40482b;
      19269: inst = 32'h8220000;
      19270: inst = 32'h10408000;
      19271: inst = 32'hc40482c;
      19272: inst = 32'h8220000;
      19273: inst = 32'h10408000;
      19274: inst = 32'hc40482e;
      19275: inst = 32'h8220000;
      19276: inst = 32'h10408000;
      19277: inst = 32'hc40482f;
      19278: inst = 32'h8220000;
      19279: inst = 32'h10408000;
      19280: inst = 32'hc404830;
      19281: inst = 32'h8220000;
      19282: inst = 32'h10408000;
      19283: inst = 32'hc404831;
      19284: inst = 32'h8220000;
      19285: inst = 32'h10408000;
      19286: inst = 32'hc404832;
      19287: inst = 32'h8220000;
      19288: inst = 32'h10408000;
      19289: inst = 32'hc404837;
      19290: inst = 32'h8220000;
      19291: inst = 32'h10408000;
      19292: inst = 32'hc404838;
      19293: inst = 32'h8220000;
      19294: inst = 32'h10408000;
      19295: inst = 32'hc40483a;
      19296: inst = 32'h8220000;
      19297: inst = 32'h10408000;
      19298: inst = 32'hc40483b;
      19299: inst = 32'h8220000;
      19300: inst = 32'h10408000;
      19301: inst = 32'hc40483c;
      19302: inst = 32'h8220000;
      19303: inst = 32'h10408000;
      19304: inst = 32'hc40483d;
      19305: inst = 32'h8220000;
      19306: inst = 32'h10408000;
      19307: inst = 32'hc40483e;
      19308: inst = 32'h8220000;
      19309: inst = 32'h10408000;
      19310: inst = 32'hc404846;
      19311: inst = 32'h8220000;
      19312: inst = 32'h10408000;
      19313: inst = 32'hc404847;
      19314: inst = 32'h8220000;
      19315: inst = 32'h10408000;
      19316: inst = 32'hc404848;
      19317: inst = 32'h8220000;
      19318: inst = 32'h10408000;
      19319: inst = 32'hc404850;
      19320: inst = 32'h8220000;
      19321: inst = 32'h10408000;
      19322: inst = 32'hc404851;
      19323: inst = 32'h8220000;
      19324: inst = 32'h10408000;
      19325: inst = 32'hc404859;
      19326: inst = 32'h8220000;
      19327: inst = 32'h10408000;
      19328: inst = 32'hc40485a;
      19329: inst = 32'h8220000;
      19330: inst = 32'h10408000;
      19331: inst = 32'hc40485f;
      19332: inst = 32'h8220000;
      19333: inst = 32'h10408000;
      19334: inst = 32'hc404860;
      19335: inst = 32'h8220000;
      19336: inst = 32'h10408000;
      19337: inst = 32'hc404861;
      19338: inst = 32'h8220000;
      19339: inst = 32'h10408000;
      19340: inst = 32'hc404862;
      19341: inst = 32'h8220000;
      19342: inst = 32'h10408000;
      19343: inst = 32'hc404869;
      19344: inst = 32'h8220000;
      19345: inst = 32'h10408000;
      19346: inst = 32'hc40486a;
      19347: inst = 32'h8220000;
      19348: inst = 32'h10408000;
      19349: inst = 32'hc40486c;
      19350: inst = 32'h8220000;
      19351: inst = 32'h10408000;
      19352: inst = 32'hc40486d;
      19353: inst = 32'h8220000;
      19354: inst = 32'h10408000;
      19355: inst = 32'hc40486e;
      19356: inst = 32'h8220000;
      19357: inst = 32'h10408000;
      19358: inst = 32'hc40486f;
      19359: inst = 32'h8220000;
      19360: inst = 32'h10408000;
      19361: inst = 32'hc404870;
      19362: inst = 32'h8220000;
      19363: inst = 32'h10408000;
      19364: inst = 32'hc404871;
      19365: inst = 32'h8220000;
      19366: inst = 32'h10408000;
      19367: inst = 32'hc404872;
      19368: inst = 32'h8220000;
      19369: inst = 32'h10408000;
      19370: inst = 32'hc40488b;
      19371: inst = 32'h8220000;
      19372: inst = 32'h10408000;
      19373: inst = 32'hc40488c;
      19374: inst = 32'h8220000;
      19375: inst = 32'h10408000;
      19376: inst = 32'hc404897;
      19377: inst = 32'h8220000;
      19378: inst = 32'h10408000;
      19379: inst = 32'hc404898;
      19380: inst = 32'h8220000;
      19381: inst = 32'h10408000;
      19382: inst = 32'hc4048a6;
      19383: inst = 32'h8220000;
      19384: inst = 32'h10408000;
      19385: inst = 32'hc4048b0;
      19386: inst = 32'h8220000;
      19387: inst = 32'h10408000;
      19388: inst = 32'hc4048b1;
      19389: inst = 32'h8220000;
      19390: inst = 32'h10408000;
      19391: inst = 32'hc4048b4;
      19392: inst = 32'h8220000;
      19393: inst = 32'h10408000;
      19394: inst = 32'hc4048b5;
      19395: inst = 32'h8220000;
      19396: inst = 32'h10408000;
      19397: inst = 32'hc4048b9;
      19398: inst = 32'h8220000;
      19399: inst = 32'h10408000;
      19400: inst = 32'hc4048ba;
      19401: inst = 32'h8220000;
      19402: inst = 32'h10408000;
      19403: inst = 32'hc4048bf;
      19404: inst = 32'h8220000;
      19405: inst = 32'h10408000;
      19406: inst = 32'hc4048c9;
      19407: inst = 32'h8220000;
      19408: inst = 32'h10408000;
      19409: inst = 32'hc4048ca;
      19410: inst = 32'h8220000;
      19411: inst = 32'h10408000;
      19412: inst = 32'hc4048d1;
      19413: inst = 32'h8220000;
      19414: inst = 32'h10408000;
      19415: inst = 32'hc4048d2;
      19416: inst = 32'h8220000;
      19417: inst = 32'h10408000;
      19418: inst = 32'hc4048d3;
      19419: inst = 32'h8220000;
      19420: inst = 32'h10408000;
      19421: inst = 32'hc4048eb;
      19422: inst = 32'h8220000;
      19423: inst = 32'h10408000;
      19424: inst = 32'hc4048ec;
      19425: inst = 32'h8220000;
      19426: inst = 32'h10408000;
      19427: inst = 32'hc4048ed;
      19428: inst = 32'h8220000;
      19429: inst = 32'h10408000;
      19430: inst = 32'hc4048ee;
      19431: inst = 32'h8220000;
      19432: inst = 32'h10408000;
      19433: inst = 32'hc4048ef;
      19434: inst = 32'h8220000;
      19435: inst = 32'h10408000;
      19436: inst = 32'hc4048f0;
      19437: inst = 32'h8220000;
      19438: inst = 32'h10408000;
      19439: inst = 32'hc4048f1;
      19440: inst = 32'h8220000;
      19441: inst = 32'h10408000;
      19442: inst = 32'hc4048f2;
      19443: inst = 32'h8220000;
      19444: inst = 32'h10408000;
      19445: inst = 32'hc4048f3;
      19446: inst = 32'h8220000;
      19447: inst = 32'h10408000;
      19448: inst = 32'hc4048f4;
      19449: inst = 32'h8220000;
      19450: inst = 32'h10408000;
      19451: inst = 32'hc4048f5;
      19452: inst = 32'h8220000;
      19453: inst = 32'h10408000;
      19454: inst = 32'hc4048f7;
      19455: inst = 32'h8220000;
      19456: inst = 32'h10408000;
      19457: inst = 32'hc4048f8;
      19458: inst = 32'h8220000;
      19459: inst = 32'h10408000;
      19460: inst = 32'hc4048f9;
      19461: inst = 32'h8220000;
      19462: inst = 32'h10408000;
      19463: inst = 32'hc4048fa;
      19464: inst = 32'h8220000;
      19465: inst = 32'h10408000;
      19466: inst = 32'hc4048fb;
      19467: inst = 32'h8220000;
      19468: inst = 32'h10408000;
      19469: inst = 32'hc4048fc;
      19470: inst = 32'h8220000;
      19471: inst = 32'h10408000;
      19472: inst = 32'hc4048fd;
      19473: inst = 32'h8220000;
      19474: inst = 32'h10408000;
      19475: inst = 32'hc4048fe;
      19476: inst = 32'h8220000;
      19477: inst = 32'h10408000;
      19478: inst = 32'hc4048ff;
      19479: inst = 32'h8220000;
      19480: inst = 32'h10408000;
      19481: inst = 32'hc404900;
      19482: inst = 32'h8220000;
      19483: inst = 32'h10408000;
      19484: inst = 32'hc404901;
      19485: inst = 32'h8220000;
      19486: inst = 32'h10408000;
      19487: inst = 32'hc404904;
      19488: inst = 32'h8220000;
      19489: inst = 32'h10408000;
      19490: inst = 32'hc404905;
      19491: inst = 32'h8220000;
      19492: inst = 32'h10408000;
      19493: inst = 32'hc404906;
      19494: inst = 32'h8220000;
      19495: inst = 32'h10408000;
      19496: inst = 32'hc404907;
      19497: inst = 32'h8220000;
      19498: inst = 32'h10408000;
      19499: inst = 32'hc404908;
      19500: inst = 32'h8220000;
      19501: inst = 32'h10408000;
      19502: inst = 32'hc404909;
      19503: inst = 32'h8220000;
      19504: inst = 32'h10408000;
      19505: inst = 32'hc40490a;
      19506: inst = 32'h8220000;
      19507: inst = 32'h10408000;
      19508: inst = 32'hc40490b;
      19509: inst = 32'h8220000;
      19510: inst = 32'h10408000;
      19511: inst = 32'hc40490c;
      19512: inst = 32'h8220000;
      19513: inst = 32'h10408000;
      19514: inst = 32'hc40490d;
      19515: inst = 32'h8220000;
      19516: inst = 32'h10408000;
      19517: inst = 32'hc404910;
      19518: inst = 32'h8220000;
      19519: inst = 32'h10408000;
      19520: inst = 32'hc404911;
      19521: inst = 32'h8220000;
      19522: inst = 32'h10408000;
      19523: inst = 32'hc404912;
      19524: inst = 32'h8220000;
      19525: inst = 32'h10408000;
      19526: inst = 32'hc404913;
      19527: inst = 32'h8220000;
      19528: inst = 32'h10408000;
      19529: inst = 32'hc404914;
      19530: inst = 32'h8220000;
      19531: inst = 32'h10408000;
      19532: inst = 32'hc404915;
      19533: inst = 32'h8220000;
      19534: inst = 32'h10408000;
      19535: inst = 32'hc404916;
      19536: inst = 32'h8220000;
      19537: inst = 32'h10408000;
      19538: inst = 32'hc404917;
      19539: inst = 32'h8220000;
      19540: inst = 32'h10408000;
      19541: inst = 32'hc404918;
      19542: inst = 32'h8220000;
      19543: inst = 32'h10408000;
      19544: inst = 32'hc404919;
      19545: inst = 32'h8220000;
      19546: inst = 32'h10408000;
      19547: inst = 32'hc40491a;
      19548: inst = 32'h8220000;
      19549: inst = 32'h10408000;
      19550: inst = 32'hc40491e;
      19551: inst = 32'h8220000;
      19552: inst = 32'h10408000;
      19553: inst = 32'hc40491f;
      19554: inst = 32'h8220000;
      19555: inst = 32'h10408000;
      19556: inst = 32'hc404920;
      19557: inst = 32'h8220000;
      19558: inst = 32'h10408000;
      19559: inst = 32'hc404921;
      19560: inst = 32'h8220000;
      19561: inst = 32'h10408000;
      19562: inst = 32'hc404922;
      19563: inst = 32'h8220000;
      19564: inst = 32'h10408000;
      19565: inst = 32'hc404923;
      19566: inst = 32'h8220000;
      19567: inst = 32'h10408000;
      19568: inst = 32'hc404924;
      19569: inst = 32'h8220000;
      19570: inst = 32'h10408000;
      19571: inst = 32'hc404925;
      19572: inst = 32'h8220000;
      19573: inst = 32'h10408000;
      19574: inst = 32'hc404926;
      19575: inst = 32'h8220000;
      19576: inst = 32'h10408000;
      19577: inst = 32'hc404927;
      19578: inst = 32'h8220000;
      19579: inst = 32'h10408000;
      19580: inst = 32'hc404929;
      19581: inst = 32'h8220000;
      19582: inst = 32'h10408000;
      19583: inst = 32'hc40492a;
      19584: inst = 32'h8220000;
      19585: inst = 32'h10408000;
      19586: inst = 32'hc40492b;
      19587: inst = 32'h8220000;
      19588: inst = 32'h10408000;
      19589: inst = 32'hc40492c;
      19590: inst = 32'h8220000;
      19591: inst = 32'h10408000;
      19592: inst = 32'hc40492d;
      19593: inst = 32'h8220000;
      19594: inst = 32'h10408000;
      19595: inst = 32'hc40492e;
      19596: inst = 32'h8220000;
      19597: inst = 32'h10408000;
      19598: inst = 32'hc40492f;
      19599: inst = 32'h8220000;
      19600: inst = 32'h10408000;
      19601: inst = 32'hc404930;
      19602: inst = 32'h8220000;
      19603: inst = 32'h10408000;
      19604: inst = 32'hc404931;
      19605: inst = 32'h8220000;
      19606: inst = 32'h10408000;
      19607: inst = 32'hc404932;
      19608: inst = 32'h8220000;
      19609: inst = 32'h10408000;
      19610: inst = 32'hc404933;
      19611: inst = 32'h8220000;
      19612: inst = 32'h10408000;
      19613: inst = 32'hc40494b;
      19614: inst = 32'h8220000;
      19615: inst = 32'h10408000;
      19616: inst = 32'hc40494c;
      19617: inst = 32'h8220000;
      19618: inst = 32'h10408000;
      19619: inst = 32'hc40494d;
      19620: inst = 32'h8220000;
      19621: inst = 32'h10408000;
      19622: inst = 32'hc40494e;
      19623: inst = 32'h8220000;
      19624: inst = 32'h10408000;
      19625: inst = 32'hc40494f;
      19626: inst = 32'h8220000;
      19627: inst = 32'h10408000;
      19628: inst = 32'hc404950;
      19629: inst = 32'h8220000;
      19630: inst = 32'h10408000;
      19631: inst = 32'hc404951;
      19632: inst = 32'h8220000;
      19633: inst = 32'h10408000;
      19634: inst = 32'hc404952;
      19635: inst = 32'h8220000;
      19636: inst = 32'h10408000;
      19637: inst = 32'hc404953;
      19638: inst = 32'h8220000;
      19639: inst = 32'h10408000;
      19640: inst = 32'hc404954;
      19641: inst = 32'h8220000;
      19642: inst = 32'h10408000;
      19643: inst = 32'hc404957;
      19644: inst = 32'h8220000;
      19645: inst = 32'h10408000;
      19646: inst = 32'hc404958;
      19647: inst = 32'h8220000;
      19648: inst = 32'h10408000;
      19649: inst = 32'hc404959;
      19650: inst = 32'h8220000;
      19651: inst = 32'h10408000;
      19652: inst = 32'hc40495a;
      19653: inst = 32'h8220000;
      19654: inst = 32'h10408000;
      19655: inst = 32'hc40495b;
      19656: inst = 32'h8220000;
      19657: inst = 32'h10408000;
      19658: inst = 32'hc40495c;
      19659: inst = 32'h8220000;
      19660: inst = 32'h10408000;
      19661: inst = 32'hc40495d;
      19662: inst = 32'h8220000;
      19663: inst = 32'h10408000;
      19664: inst = 32'hc40495e;
      19665: inst = 32'h8220000;
      19666: inst = 32'h10408000;
      19667: inst = 32'hc40495f;
      19668: inst = 32'h8220000;
      19669: inst = 32'h10408000;
      19670: inst = 32'hc404960;
      19671: inst = 32'h8220000;
      19672: inst = 32'h10408000;
      19673: inst = 32'hc404961;
      19674: inst = 32'h8220000;
      19675: inst = 32'h10408000;
      19676: inst = 32'hc404963;
      19677: inst = 32'h8220000;
      19678: inst = 32'h10408000;
      19679: inst = 32'hc404964;
      19680: inst = 32'h8220000;
      19681: inst = 32'h10408000;
      19682: inst = 32'hc404965;
      19683: inst = 32'h8220000;
      19684: inst = 32'h10408000;
      19685: inst = 32'hc404966;
      19686: inst = 32'h8220000;
      19687: inst = 32'h10408000;
      19688: inst = 32'hc404967;
      19689: inst = 32'h8220000;
      19690: inst = 32'h10408000;
      19691: inst = 32'hc404968;
      19692: inst = 32'h8220000;
      19693: inst = 32'h10408000;
      19694: inst = 32'hc404969;
      19695: inst = 32'h8220000;
      19696: inst = 32'h10408000;
      19697: inst = 32'hc40496a;
      19698: inst = 32'h8220000;
      19699: inst = 32'h10408000;
      19700: inst = 32'hc40496b;
      19701: inst = 32'h8220000;
      19702: inst = 32'h10408000;
      19703: inst = 32'hc40496c;
      19704: inst = 32'h8220000;
      19705: inst = 32'h10408000;
      19706: inst = 32'hc40496d;
      19707: inst = 32'h8220000;
      19708: inst = 32'h10408000;
      19709: inst = 32'hc404970;
      19710: inst = 32'h8220000;
      19711: inst = 32'h10408000;
      19712: inst = 32'hc404971;
      19713: inst = 32'h8220000;
      19714: inst = 32'h10408000;
      19715: inst = 32'hc404972;
      19716: inst = 32'h8220000;
      19717: inst = 32'h10408000;
      19718: inst = 32'hc404973;
      19719: inst = 32'h8220000;
      19720: inst = 32'h10408000;
      19721: inst = 32'hc404974;
      19722: inst = 32'h8220000;
      19723: inst = 32'h10408000;
      19724: inst = 32'hc404975;
      19725: inst = 32'h8220000;
      19726: inst = 32'h10408000;
      19727: inst = 32'hc404976;
      19728: inst = 32'h8220000;
      19729: inst = 32'h10408000;
      19730: inst = 32'hc404977;
      19731: inst = 32'h8220000;
      19732: inst = 32'h10408000;
      19733: inst = 32'hc404978;
      19734: inst = 32'h8220000;
      19735: inst = 32'h10408000;
      19736: inst = 32'hc404979;
      19737: inst = 32'h8220000;
      19738: inst = 32'h10408000;
      19739: inst = 32'hc40497d;
      19740: inst = 32'h8220000;
      19741: inst = 32'h10408000;
      19742: inst = 32'hc40497e;
      19743: inst = 32'h8220000;
      19744: inst = 32'h10408000;
      19745: inst = 32'hc40497f;
      19746: inst = 32'h8220000;
      19747: inst = 32'h10408000;
      19748: inst = 32'hc404980;
      19749: inst = 32'h8220000;
      19750: inst = 32'h10408000;
      19751: inst = 32'hc404981;
      19752: inst = 32'h8220000;
      19753: inst = 32'h10408000;
      19754: inst = 32'hc404982;
      19755: inst = 32'h8220000;
      19756: inst = 32'h10408000;
      19757: inst = 32'hc404983;
      19758: inst = 32'h8220000;
      19759: inst = 32'h10408000;
      19760: inst = 32'hc404984;
      19761: inst = 32'h8220000;
      19762: inst = 32'h10408000;
      19763: inst = 32'hc404985;
      19764: inst = 32'h8220000;
      19765: inst = 32'h10408000;
      19766: inst = 32'hc404986;
      19767: inst = 32'h8220000;
      19768: inst = 32'h10408000;
      19769: inst = 32'hc404987;
      19770: inst = 32'h8220000;
      19771: inst = 32'h10408000;
      19772: inst = 32'hc404989;
      19773: inst = 32'h8220000;
      19774: inst = 32'h10408000;
      19775: inst = 32'hc40498a;
      19776: inst = 32'h8220000;
      19777: inst = 32'h10408000;
      19778: inst = 32'hc40498b;
      19779: inst = 32'h8220000;
      19780: inst = 32'h10408000;
      19781: inst = 32'hc40498c;
      19782: inst = 32'h8220000;
      19783: inst = 32'h10408000;
      19784: inst = 32'hc40498d;
      19785: inst = 32'h8220000;
      19786: inst = 32'h10408000;
      19787: inst = 32'hc40498e;
      19788: inst = 32'h8220000;
      19789: inst = 32'h10408000;
      19790: inst = 32'hc40498f;
      19791: inst = 32'h8220000;
      19792: inst = 32'h10408000;
      19793: inst = 32'hc404990;
      19794: inst = 32'h8220000;
      19795: inst = 32'h10408000;
      19796: inst = 32'hc404991;
      19797: inst = 32'h8220000;
      19798: inst = 32'h10408000;
      19799: inst = 32'hc404992;
      19800: inst = 32'h8220000;
      19801: inst = 32'h10408000;
      19802: inst = 32'hc404993;
      19803: inst = 32'h8220000;
      19804: inst = 32'h10408000;
      19805: inst = 32'hc404dcd;
      19806: inst = 32'h8220000;
      19807: inst = 32'h10408000;
      19808: inst = 32'hc404dce;
      19809: inst = 32'h8220000;
      19810: inst = 32'h10408000;
      19811: inst = 32'hc404dcf;
      19812: inst = 32'h8220000;
      19813: inst = 32'h10408000;
      19814: inst = 32'hc404dd0;
      19815: inst = 32'h8220000;
      19816: inst = 32'h10408000;
      19817: inst = 32'hc404dd1;
      19818: inst = 32'h8220000;
      19819: inst = 32'h10408000;
      19820: inst = 32'hc404dd2;
      19821: inst = 32'h8220000;
      19822: inst = 32'h10408000;
      19823: inst = 32'hc404dd3;
      19824: inst = 32'h8220000;
      19825: inst = 32'h10408000;
      19826: inst = 32'hc404dd4;
      19827: inst = 32'h8220000;
      19828: inst = 32'h10408000;
      19829: inst = 32'hc404dd5;
      19830: inst = 32'h8220000;
      19831: inst = 32'h10408000;
      19832: inst = 32'hc404dd7;
      19833: inst = 32'h8220000;
      19834: inst = 32'h10408000;
      19835: inst = 32'hc404dd8;
      19836: inst = 32'h8220000;
      19837: inst = 32'h10408000;
      19838: inst = 32'hc404dd9;
      19839: inst = 32'h8220000;
      19840: inst = 32'h10408000;
      19841: inst = 32'hc404dda;
      19842: inst = 32'h8220000;
      19843: inst = 32'h10408000;
      19844: inst = 32'hc404ddb;
      19845: inst = 32'h8220000;
      19846: inst = 32'h10408000;
      19847: inst = 32'hc404ddc;
      19848: inst = 32'h8220000;
      19849: inst = 32'h10408000;
      19850: inst = 32'hc404ddd;
      19851: inst = 32'h8220000;
      19852: inst = 32'h10408000;
      19853: inst = 32'hc404dde;
      19854: inst = 32'h8220000;
      19855: inst = 32'h10408000;
      19856: inst = 32'hc404ddf;
      19857: inst = 32'h8220000;
      19858: inst = 32'h10408000;
      19859: inst = 32'hc404de0;
      19860: inst = 32'h8220000;
      19861: inst = 32'h10408000;
      19862: inst = 32'hc404de1;
      19863: inst = 32'h8220000;
      19864: inst = 32'h10408000;
      19865: inst = 32'hc404de2;
      19866: inst = 32'h8220000;
      19867: inst = 32'h10408000;
      19868: inst = 32'hc404de4;
      19869: inst = 32'h8220000;
      19870: inst = 32'h10408000;
      19871: inst = 32'hc404de5;
      19872: inst = 32'h8220000;
      19873: inst = 32'h10408000;
      19874: inst = 32'hc404de6;
      19875: inst = 32'h8220000;
      19876: inst = 32'h10408000;
      19877: inst = 32'hc404de7;
      19878: inst = 32'h8220000;
      19879: inst = 32'h10408000;
      19880: inst = 32'hc404de8;
      19881: inst = 32'h8220000;
      19882: inst = 32'h10408000;
      19883: inst = 32'hc404de9;
      19884: inst = 32'h8220000;
      19885: inst = 32'h10408000;
      19886: inst = 32'hc404dea;
      19887: inst = 32'h8220000;
      19888: inst = 32'h10408000;
      19889: inst = 32'hc404deb;
      19890: inst = 32'h8220000;
      19891: inst = 32'h10408000;
      19892: inst = 32'hc404dec;
      19893: inst = 32'h8220000;
      19894: inst = 32'h10408000;
      19895: inst = 32'hc404ded;
      19896: inst = 32'h8220000;
      19897: inst = 32'h10408000;
      19898: inst = 32'hc404df0;
      19899: inst = 32'h8220000;
      19900: inst = 32'h10408000;
      19901: inst = 32'hc404df1;
      19902: inst = 32'h8220000;
      19903: inst = 32'h10408000;
      19904: inst = 32'hc404df2;
      19905: inst = 32'h8220000;
      19906: inst = 32'h10408000;
      19907: inst = 32'hc404dfc;
      19908: inst = 32'h8220000;
      19909: inst = 32'h10408000;
      19910: inst = 32'hc404dfd;
      19911: inst = 32'h8220000;
      19912: inst = 32'h10408000;
      19913: inst = 32'hc404dfe;
      19914: inst = 32'h8220000;
      19915: inst = 32'h10408000;
      19916: inst = 32'hc404dff;
      19917: inst = 32'h8220000;
      19918: inst = 32'h10408000;
      19919: inst = 32'hc404e00;
      19920: inst = 32'h8220000;
      19921: inst = 32'h10408000;
      19922: inst = 32'hc404e01;
      19923: inst = 32'h8220000;
      19924: inst = 32'h10408000;
      19925: inst = 32'hc404e02;
      19926: inst = 32'h8220000;
      19927: inst = 32'h10408000;
      19928: inst = 32'hc404e03;
      19929: inst = 32'h8220000;
      19930: inst = 32'h10408000;
      19931: inst = 32'hc404e04;
      19932: inst = 32'h8220000;
      19933: inst = 32'h10408000;
      19934: inst = 32'hc404e05;
      19935: inst = 32'h8220000;
      19936: inst = 32'h10408000;
      19937: inst = 32'hc404e06;
      19938: inst = 32'h8220000;
      19939: inst = 32'h10408000;
      19940: inst = 32'hc404e07;
      19941: inst = 32'h8220000;
      19942: inst = 32'h10408000;
      19943: inst = 32'hc404e0b;
      19944: inst = 32'h8220000;
      19945: inst = 32'h10408000;
      19946: inst = 32'hc404e0c;
      19947: inst = 32'h8220000;
      19948: inst = 32'h10408000;
      19949: inst = 32'hc404e0d;
      19950: inst = 32'h8220000;
      19951: inst = 32'h10408000;
      19952: inst = 32'hc404e0e;
      19953: inst = 32'h8220000;
      19954: inst = 32'h10408000;
      19955: inst = 32'hc404e0f;
      19956: inst = 32'h8220000;
      19957: inst = 32'h10408000;
      19958: inst = 32'hc404e10;
      19959: inst = 32'h8220000;
      19960: inst = 32'h10408000;
      19961: inst = 32'hc404e11;
      19962: inst = 32'h8220000;
      19963: inst = 32'h10408000;
      19964: inst = 32'hc404e12;
      19965: inst = 32'h8220000;
      19966: inst = 32'h10408000;
      19967: inst = 32'hc404e13;
      19968: inst = 32'h8220000;
      19969: inst = 32'h10408000;
      19970: inst = 32'hc404e2c;
      19971: inst = 32'h8220000;
      19972: inst = 32'h10408000;
      19973: inst = 32'hc404e2d;
      19974: inst = 32'h8220000;
      19975: inst = 32'h10408000;
      19976: inst = 32'hc404e2e;
      19977: inst = 32'h8220000;
      19978: inst = 32'h10408000;
      19979: inst = 32'hc404e2f;
      19980: inst = 32'h8220000;
      19981: inst = 32'h10408000;
      19982: inst = 32'hc404e30;
      19983: inst = 32'h8220000;
      19984: inst = 32'h10408000;
      19985: inst = 32'hc404e31;
      19986: inst = 32'h8220000;
      19987: inst = 32'h10408000;
      19988: inst = 32'hc404e32;
      19989: inst = 32'h8220000;
      19990: inst = 32'h10408000;
      19991: inst = 32'hc404e33;
      19992: inst = 32'h8220000;
      19993: inst = 32'h10408000;
      19994: inst = 32'hc404e34;
      19995: inst = 32'h8220000;
      19996: inst = 32'h10408000;
      19997: inst = 32'hc404e35;
      19998: inst = 32'h8220000;
      19999: inst = 32'h10408000;
      20000: inst = 32'hc404e38;
      20001: inst = 32'h8220000;
      20002: inst = 32'h10408000;
      20003: inst = 32'hc404e39;
      20004: inst = 32'h8220000;
      20005: inst = 32'h10408000;
      20006: inst = 32'hc404e3a;
      20007: inst = 32'h8220000;
      20008: inst = 32'h10408000;
      20009: inst = 32'hc404e3b;
      20010: inst = 32'h8220000;
      20011: inst = 32'h10408000;
      20012: inst = 32'hc404e3c;
      20013: inst = 32'h8220000;
      20014: inst = 32'h10408000;
      20015: inst = 32'hc404e3d;
      20016: inst = 32'h8220000;
      20017: inst = 32'h10408000;
      20018: inst = 32'hc404e3e;
      20019: inst = 32'h8220000;
      20020: inst = 32'h10408000;
      20021: inst = 32'hc404e3f;
      20022: inst = 32'h8220000;
      20023: inst = 32'h10408000;
      20024: inst = 32'hc404e40;
      20025: inst = 32'h8220000;
      20026: inst = 32'h10408000;
      20027: inst = 32'hc404e41;
      20028: inst = 32'h8220000;
      20029: inst = 32'h10408000;
      20030: inst = 32'hc404e42;
      20031: inst = 32'h8220000;
      20032: inst = 32'h10408000;
      20033: inst = 32'hc404e44;
      20034: inst = 32'h8220000;
      20035: inst = 32'h10408000;
      20036: inst = 32'hc404e45;
      20037: inst = 32'h8220000;
      20038: inst = 32'h10408000;
      20039: inst = 32'hc404e46;
      20040: inst = 32'h8220000;
      20041: inst = 32'h10408000;
      20042: inst = 32'hc404e47;
      20043: inst = 32'h8220000;
      20044: inst = 32'h10408000;
      20045: inst = 32'hc404e48;
      20046: inst = 32'h8220000;
      20047: inst = 32'h10408000;
      20048: inst = 32'hc404e49;
      20049: inst = 32'h8220000;
      20050: inst = 32'h10408000;
      20051: inst = 32'hc404e4a;
      20052: inst = 32'h8220000;
      20053: inst = 32'h10408000;
      20054: inst = 32'hc404e4b;
      20055: inst = 32'h8220000;
      20056: inst = 32'h10408000;
      20057: inst = 32'hc404e4c;
      20058: inst = 32'h8220000;
      20059: inst = 32'h10408000;
      20060: inst = 32'hc404e4d;
      20061: inst = 32'h8220000;
      20062: inst = 32'h10408000;
      20063: inst = 32'hc404e50;
      20064: inst = 32'h8220000;
      20065: inst = 32'h10408000;
      20066: inst = 32'hc404e51;
      20067: inst = 32'h8220000;
      20068: inst = 32'h10408000;
      20069: inst = 32'hc404e52;
      20070: inst = 32'h8220000;
      20071: inst = 32'h10408000;
      20072: inst = 32'hc404e53;
      20073: inst = 32'h8220000;
      20074: inst = 32'h10408000;
      20075: inst = 32'hc404e5c;
      20076: inst = 32'h8220000;
      20077: inst = 32'h10408000;
      20078: inst = 32'hc404e5d;
      20079: inst = 32'h8220000;
      20080: inst = 32'h10408000;
      20081: inst = 32'hc404e5e;
      20082: inst = 32'h8220000;
      20083: inst = 32'h10408000;
      20084: inst = 32'hc404e5f;
      20085: inst = 32'h8220000;
      20086: inst = 32'h10408000;
      20087: inst = 32'hc404e60;
      20088: inst = 32'h8220000;
      20089: inst = 32'h10408000;
      20090: inst = 32'hc404e61;
      20091: inst = 32'h8220000;
      20092: inst = 32'h10408000;
      20093: inst = 32'hc404e62;
      20094: inst = 32'h8220000;
      20095: inst = 32'h10408000;
      20096: inst = 32'hc404e63;
      20097: inst = 32'h8220000;
      20098: inst = 32'h10408000;
      20099: inst = 32'hc404e64;
      20100: inst = 32'h8220000;
      20101: inst = 32'h10408000;
      20102: inst = 32'hc404e65;
      20103: inst = 32'h8220000;
      20104: inst = 32'h10408000;
      20105: inst = 32'hc404e66;
      20106: inst = 32'h8220000;
      20107: inst = 32'h10408000;
      20108: inst = 32'hc404e6a;
      20109: inst = 32'h8220000;
      20110: inst = 32'h10408000;
      20111: inst = 32'hc404e6b;
      20112: inst = 32'h8220000;
      20113: inst = 32'h10408000;
      20114: inst = 32'hc404e6c;
      20115: inst = 32'h8220000;
      20116: inst = 32'h10408000;
      20117: inst = 32'hc404e6d;
      20118: inst = 32'h8220000;
      20119: inst = 32'h10408000;
      20120: inst = 32'hc404e6e;
      20121: inst = 32'h8220000;
      20122: inst = 32'h10408000;
      20123: inst = 32'hc404e6f;
      20124: inst = 32'h8220000;
      20125: inst = 32'h10408000;
      20126: inst = 32'hc404e70;
      20127: inst = 32'h8220000;
      20128: inst = 32'h10408000;
      20129: inst = 32'hc404e71;
      20130: inst = 32'h8220000;
      20131: inst = 32'h10408000;
      20132: inst = 32'hc404e72;
      20133: inst = 32'h8220000;
      20134: inst = 32'h10408000;
      20135: inst = 32'hc404e73;
      20136: inst = 32'h8220000;
      20137: inst = 32'h10408000;
      20138: inst = 32'hc404e8b;
      20139: inst = 32'h8220000;
      20140: inst = 32'h10408000;
      20141: inst = 32'hc404e8c;
      20142: inst = 32'h8220000;
      20143: inst = 32'h10408000;
      20144: inst = 32'hc404e8d;
      20145: inst = 32'h8220000;
      20146: inst = 32'h10408000;
      20147: inst = 32'hc404e99;
      20148: inst = 32'h8220000;
      20149: inst = 32'h10408000;
      20150: inst = 32'hc404e9a;
      20151: inst = 32'h8220000;
      20152: inst = 32'h10408000;
      20153: inst = 32'hc404e9b;
      20154: inst = 32'h8220000;
      20155: inst = 32'h10408000;
      20156: inst = 32'hc404e9c;
      20157: inst = 32'h8220000;
      20158: inst = 32'h10408000;
      20159: inst = 32'hc404ea4;
      20160: inst = 32'h8220000;
      20161: inst = 32'h10408000;
      20162: inst = 32'hc404ea5;
      20163: inst = 32'h8220000;
      20164: inst = 32'h10408000;
      20165: inst = 32'hc404eac;
      20166: inst = 32'h8220000;
      20167: inst = 32'h10408000;
      20168: inst = 32'hc404ead;
      20169: inst = 32'h8220000;
      20170: inst = 32'h10408000;
      20171: inst = 32'hc404eb0;
      20172: inst = 32'h8220000;
      20173: inst = 32'h10408000;
      20174: inst = 32'hc404eb1;
      20175: inst = 32'h8220000;
      20176: inst = 32'h10408000;
      20177: inst = 32'hc404eb2;
      20178: inst = 32'h8220000;
      20179: inst = 32'h10408000;
      20180: inst = 32'hc404eb3;
      20181: inst = 32'h8220000;
      20182: inst = 32'h10408000;
      20183: inst = 32'hc404eb4;
      20184: inst = 32'h8220000;
      20185: inst = 32'h10408000;
      20186: inst = 32'hc404ebc;
      20187: inst = 32'h8220000;
      20188: inst = 32'h10408000;
      20189: inst = 32'hc404ebd;
      20190: inst = 32'h8220000;
      20191: inst = 32'h10408000;
      20192: inst = 32'hc404ec2;
      20193: inst = 32'h8220000;
      20194: inst = 32'h10408000;
      20195: inst = 32'hc404ec3;
      20196: inst = 32'h8220000;
      20197: inst = 32'h10408000;
      20198: inst = 32'hc404ec4;
      20199: inst = 32'h8220000;
      20200: inst = 32'h10408000;
      20201: inst = 32'hc404ec5;
      20202: inst = 32'h8220000;
      20203: inst = 32'h10408000;
      20204: inst = 32'hc404ec9;
      20205: inst = 32'h8220000;
      20206: inst = 32'h10408000;
      20207: inst = 32'hc404eca;
      20208: inst = 32'h8220000;
      20209: inst = 32'h10408000;
      20210: inst = 32'hc404eeb;
      20211: inst = 32'h8220000;
      20212: inst = 32'h10408000;
      20213: inst = 32'hc404eec;
      20214: inst = 32'h8220000;
      20215: inst = 32'h10408000;
      20216: inst = 32'hc404efa;
      20217: inst = 32'h8220000;
      20218: inst = 32'h10408000;
      20219: inst = 32'hc404efb;
      20220: inst = 32'h8220000;
      20221: inst = 32'h10408000;
      20222: inst = 32'hc404efc;
      20223: inst = 32'h8220000;
      20224: inst = 32'h10408000;
      20225: inst = 32'hc404f04;
      20226: inst = 32'h8220000;
      20227: inst = 32'h10408000;
      20228: inst = 32'hc404f05;
      20229: inst = 32'h8220000;
      20230: inst = 32'h10408000;
      20231: inst = 32'hc404f0c;
      20232: inst = 32'h8220000;
      20233: inst = 32'h10408000;
      20234: inst = 32'hc404f0d;
      20235: inst = 32'h8220000;
      20236: inst = 32'h10408000;
      20237: inst = 32'hc404f10;
      20238: inst = 32'h8220000;
      20239: inst = 32'h10408000;
      20240: inst = 32'hc404f12;
      20241: inst = 32'h8220000;
      20242: inst = 32'h10408000;
      20243: inst = 32'hc404f13;
      20244: inst = 32'h8220000;
      20245: inst = 32'h10408000;
      20246: inst = 32'hc404f14;
      20247: inst = 32'h8220000;
      20248: inst = 32'h10408000;
      20249: inst = 32'hc404f15;
      20250: inst = 32'h8220000;
      20251: inst = 32'h10408000;
      20252: inst = 32'hc404f1c;
      20253: inst = 32'h8220000;
      20254: inst = 32'h10408000;
      20255: inst = 32'hc404f1d;
      20256: inst = 32'h8220000;
      20257: inst = 32'h10408000;
      20258: inst = 32'hc404f22;
      20259: inst = 32'h8220000;
      20260: inst = 32'h10408000;
      20261: inst = 32'hc404f23;
      20262: inst = 32'h8220000;
      20263: inst = 32'h10408000;
      20264: inst = 32'hc404f24;
      20265: inst = 32'h8220000;
      20266: inst = 32'h10408000;
      20267: inst = 32'hc404f29;
      20268: inst = 32'h8220000;
      20269: inst = 32'h10408000;
      20270: inst = 32'hc404f2a;
      20271: inst = 32'h8220000;
      20272: inst = 32'h10408000;
      20273: inst = 32'hc404f4b;
      20274: inst = 32'h8220000;
      20275: inst = 32'h10408000;
      20276: inst = 32'hc404f4c;
      20277: inst = 32'h8220000;
      20278: inst = 32'h10408000;
      20279: inst = 32'hc404f4e;
      20280: inst = 32'h8220000;
      20281: inst = 32'h10408000;
      20282: inst = 32'hc404f4f;
      20283: inst = 32'h8220000;
      20284: inst = 32'h10408000;
      20285: inst = 32'hc404f50;
      20286: inst = 32'h8220000;
      20287: inst = 32'h10408000;
      20288: inst = 32'hc404f51;
      20289: inst = 32'h8220000;
      20290: inst = 32'h10408000;
      20291: inst = 32'hc404f52;
      20292: inst = 32'h8220000;
      20293: inst = 32'h10408000;
      20294: inst = 32'hc404f5b;
      20295: inst = 32'h8220000;
      20296: inst = 32'h10408000;
      20297: inst = 32'hc404f5c;
      20298: inst = 32'h8220000;
      20299: inst = 32'h10408000;
      20300: inst = 32'hc404f5d;
      20301: inst = 32'h8220000;
      20302: inst = 32'h10408000;
      20303: inst = 32'hc404f64;
      20304: inst = 32'h8220000;
      20305: inst = 32'h10408000;
      20306: inst = 32'hc404f65;
      20307: inst = 32'h8220000;
      20308: inst = 32'h10408000;
      20309: inst = 32'hc404f6c;
      20310: inst = 32'h8220000;
      20311: inst = 32'h10408000;
      20312: inst = 32'hc404f70;
      20313: inst = 32'h8220000;
      20314: inst = 32'h10408000;
      20315: inst = 32'hc404f71;
      20316: inst = 32'h8220000;
      20317: inst = 32'h10408000;
      20318: inst = 32'hc404f72;
      20319: inst = 32'h8220000;
      20320: inst = 32'h10408000;
      20321: inst = 32'hc404f73;
      20322: inst = 32'h8220000;
      20323: inst = 32'h10408000;
      20324: inst = 32'hc404f74;
      20325: inst = 32'h8220000;
      20326: inst = 32'h10408000;
      20327: inst = 32'hc404f75;
      20328: inst = 32'h8220000;
      20329: inst = 32'h10408000;
      20330: inst = 32'hc404f76;
      20331: inst = 32'h8220000;
      20332: inst = 32'h10408000;
      20333: inst = 32'hc404f7c;
      20334: inst = 32'h8220000;
      20335: inst = 32'h10408000;
      20336: inst = 32'hc404f7d;
      20337: inst = 32'h8220000;
      20338: inst = 32'h10408000;
      20339: inst = 32'hc404f7f;
      20340: inst = 32'h8220000;
      20341: inst = 32'h10408000;
      20342: inst = 32'hc404f80;
      20343: inst = 32'h8220000;
      20344: inst = 32'h10408000;
      20345: inst = 32'hc404f81;
      20346: inst = 32'h8220000;
      20347: inst = 32'h10408000;
      20348: inst = 32'hc404f82;
      20349: inst = 32'h8220000;
      20350: inst = 32'h10408000;
      20351: inst = 32'hc404f83;
      20352: inst = 32'h8220000;
      20353: inst = 32'h10408000;
      20354: inst = 32'hc404f89;
      20355: inst = 32'h8220000;
      20356: inst = 32'h10408000;
      20357: inst = 32'hc404f8a;
      20358: inst = 32'h8220000;
      20359: inst = 32'h10408000;
      20360: inst = 32'hc404f8c;
      20361: inst = 32'h8220000;
      20362: inst = 32'h10408000;
      20363: inst = 32'hc404f8d;
      20364: inst = 32'h8220000;
      20365: inst = 32'h10408000;
      20366: inst = 32'hc404f8e;
      20367: inst = 32'h8220000;
      20368: inst = 32'h10408000;
      20369: inst = 32'hc404f8f;
      20370: inst = 32'h8220000;
      20371: inst = 32'h10408000;
      20372: inst = 32'hc404f90;
      20373: inst = 32'h8220000;
      20374: inst = 32'h10408000;
      20375: inst = 32'hc404fab;
      20376: inst = 32'h8220000;
      20377: inst = 32'h10408000;
      20378: inst = 32'hc404fac;
      20379: inst = 32'h8220000;
      20380: inst = 32'h10408000;
      20381: inst = 32'hc404fae;
      20382: inst = 32'h8220000;
      20383: inst = 32'h10408000;
      20384: inst = 32'hc404faf;
      20385: inst = 32'h8220000;
      20386: inst = 32'h10408000;
      20387: inst = 32'hc404fb0;
      20388: inst = 32'h8220000;
      20389: inst = 32'h10408000;
      20390: inst = 32'hc404fb1;
      20391: inst = 32'h8220000;
      20392: inst = 32'h10408000;
      20393: inst = 32'hc404fb2;
      20394: inst = 32'h8220000;
      20395: inst = 32'h10408000;
      20396: inst = 32'hc404fbc;
      20397: inst = 32'h8220000;
      20398: inst = 32'h10408000;
      20399: inst = 32'hc404fbd;
      20400: inst = 32'h8220000;
      20401: inst = 32'h10408000;
      20402: inst = 32'hc404fbe;
      20403: inst = 32'h8220000;
      20404: inst = 32'h10408000;
      20405: inst = 32'hc404fc4;
      20406: inst = 32'h8220000;
      20407: inst = 32'h10408000;
      20408: inst = 32'hc404fc5;
      20409: inst = 32'h8220000;
      20410: inst = 32'h10408000;
      20411: inst = 32'hc404fd0;
      20412: inst = 32'h8220000;
      20413: inst = 32'h10408000;
      20414: inst = 32'hc404fd1;
      20415: inst = 32'h8220000;
      20416: inst = 32'h10408000;
      20417: inst = 32'hc404fd2;
      20418: inst = 32'h8220000;
      20419: inst = 32'h10408000;
      20420: inst = 32'hc404fd4;
      20421: inst = 32'h8220000;
      20422: inst = 32'h10408000;
      20423: inst = 32'hc404fd5;
      20424: inst = 32'h8220000;
      20425: inst = 32'h10408000;
      20426: inst = 32'hc404fd6;
      20427: inst = 32'h8220000;
      20428: inst = 32'h10408000;
      20429: inst = 32'hc404fd7;
      20430: inst = 32'h8220000;
      20431: inst = 32'h10408000;
      20432: inst = 32'hc404fdc;
      20433: inst = 32'h8220000;
      20434: inst = 32'h10408000;
      20435: inst = 32'hc404fdd;
      20436: inst = 32'h8220000;
      20437: inst = 32'h10408000;
      20438: inst = 32'hc404fdf;
      20439: inst = 32'h8220000;
      20440: inst = 32'h10408000;
      20441: inst = 32'hc404fe0;
      20442: inst = 32'h8220000;
      20443: inst = 32'h10408000;
      20444: inst = 32'hc404fe1;
      20445: inst = 32'h8220000;
      20446: inst = 32'h10408000;
      20447: inst = 32'hc404fe2;
      20448: inst = 32'h8220000;
      20449: inst = 32'h10408000;
      20450: inst = 32'hc404fe9;
      20451: inst = 32'h8220000;
      20452: inst = 32'h10408000;
      20453: inst = 32'hc404fea;
      20454: inst = 32'h8220000;
      20455: inst = 32'h10408000;
      20456: inst = 32'hc404fec;
      20457: inst = 32'h8220000;
      20458: inst = 32'h10408000;
      20459: inst = 32'hc404fed;
      20460: inst = 32'h8220000;
      20461: inst = 32'h10408000;
      20462: inst = 32'hc404fee;
      20463: inst = 32'h8220000;
      20464: inst = 32'h10408000;
      20465: inst = 32'hc404fef;
      20466: inst = 32'h8220000;
      20467: inst = 32'h10408000;
      20468: inst = 32'hc404ff0;
      20469: inst = 32'h8220000;
      20470: inst = 32'h10408000;
      20471: inst = 32'hc40500b;
      20472: inst = 32'h8220000;
      20473: inst = 32'h10408000;
      20474: inst = 32'hc40500c;
      20475: inst = 32'h8220000;
      20476: inst = 32'h10408000;
      20477: inst = 32'hc40501d;
      20478: inst = 32'h8220000;
      20479: inst = 32'h10408000;
      20480: inst = 32'hc40501e;
      20481: inst = 32'h8220000;
      20482: inst = 32'h10408000;
      20483: inst = 32'hc40501f;
      20484: inst = 32'h8220000;
      20485: inst = 32'h10408000;
      20486: inst = 32'hc405024;
      20487: inst = 32'h8220000;
      20488: inst = 32'h10408000;
      20489: inst = 32'hc405025;
      20490: inst = 32'h8220000;
      20491: inst = 32'h10408000;
      20492: inst = 32'hc405030;
      20493: inst = 32'h8220000;
      20494: inst = 32'h10408000;
      20495: inst = 32'hc405031;
      20496: inst = 32'h8220000;
      20497: inst = 32'h10408000;
      20498: inst = 32'hc405032;
      20499: inst = 32'h8220000;
      20500: inst = 32'h10408000;
      20501: inst = 32'hc405033;
      20502: inst = 32'h8220000;
      20503: inst = 32'h10408000;
      20504: inst = 32'hc405034;
      20505: inst = 32'h8220000;
      20506: inst = 32'h10408000;
      20507: inst = 32'hc405035;
      20508: inst = 32'h8220000;
      20509: inst = 32'h10408000;
      20510: inst = 32'hc405036;
      20511: inst = 32'h8220000;
      20512: inst = 32'h10408000;
      20513: inst = 32'hc405037;
      20514: inst = 32'h8220000;
      20515: inst = 32'h10408000;
      20516: inst = 32'hc405038;
      20517: inst = 32'h8220000;
      20518: inst = 32'h10408000;
      20519: inst = 32'hc40503c;
      20520: inst = 32'h8220000;
      20521: inst = 32'h10408000;
      20522: inst = 32'hc40503d;
      20523: inst = 32'h8220000;
      20524: inst = 32'h10408000;
      20525: inst = 32'hc405049;
      20526: inst = 32'h8220000;
      20527: inst = 32'h10408000;
      20528: inst = 32'hc40504a;
      20529: inst = 32'h8220000;
      20530: inst = 32'h10408000;
      20531: inst = 32'hc40506b;
      20532: inst = 32'h8220000;
      20533: inst = 32'h10408000;
      20534: inst = 32'hc40506c;
      20535: inst = 32'h8220000;
      20536: inst = 32'h10408000;
      20537: inst = 32'hc40506d;
      20538: inst = 32'h8220000;
      20539: inst = 32'h10408000;
      20540: inst = 32'hc40506e;
      20541: inst = 32'h8220000;
      20542: inst = 32'h10408000;
      20543: inst = 32'hc40506f;
      20544: inst = 32'h8220000;
      20545: inst = 32'h10408000;
      20546: inst = 32'hc405070;
      20547: inst = 32'h8220000;
      20548: inst = 32'h10408000;
      20549: inst = 32'hc405071;
      20550: inst = 32'h8220000;
      20551: inst = 32'h10408000;
      20552: inst = 32'hc405072;
      20553: inst = 32'h8220000;
      20554: inst = 32'h10408000;
      20555: inst = 32'hc405073;
      20556: inst = 32'h8220000;
      20557: inst = 32'h10408000;
      20558: inst = 32'hc405074;
      20559: inst = 32'h8220000;
      20560: inst = 32'h10408000;
      20561: inst = 32'hc405075;
      20562: inst = 32'h8220000;
      20563: inst = 32'h10408000;
      20564: inst = 32'hc405077;
      20565: inst = 32'h8220000;
      20566: inst = 32'h10408000;
      20567: inst = 32'hc405078;
      20568: inst = 32'h8220000;
      20569: inst = 32'h10408000;
      20570: inst = 32'hc405079;
      20571: inst = 32'h8220000;
      20572: inst = 32'h10408000;
      20573: inst = 32'hc40507a;
      20574: inst = 32'h8220000;
      20575: inst = 32'h10408000;
      20576: inst = 32'hc40507b;
      20577: inst = 32'h8220000;
      20578: inst = 32'h10408000;
      20579: inst = 32'hc40507c;
      20580: inst = 32'h8220000;
      20581: inst = 32'h10408000;
      20582: inst = 32'hc40507d;
      20583: inst = 32'h8220000;
      20584: inst = 32'h10408000;
      20585: inst = 32'hc40507e;
      20586: inst = 32'h8220000;
      20587: inst = 32'h10408000;
      20588: inst = 32'hc40507f;
      20589: inst = 32'h8220000;
      20590: inst = 32'h10408000;
      20591: inst = 32'hc405080;
      20592: inst = 32'h8220000;
      20593: inst = 32'h10408000;
      20594: inst = 32'hc405084;
      20595: inst = 32'h8220000;
      20596: inst = 32'h10408000;
      20597: inst = 32'hc405085;
      20598: inst = 32'h8220000;
      20599: inst = 32'h10408000;
      20600: inst = 32'hc405086;
      20601: inst = 32'h8220000;
      20602: inst = 32'h10408000;
      20603: inst = 32'hc405087;
      20604: inst = 32'h8220000;
      20605: inst = 32'h10408000;
      20606: inst = 32'hc405088;
      20607: inst = 32'h8220000;
      20608: inst = 32'h10408000;
      20609: inst = 32'hc405089;
      20610: inst = 32'h8220000;
      20611: inst = 32'h10408000;
      20612: inst = 32'hc40508a;
      20613: inst = 32'h8220000;
      20614: inst = 32'h10408000;
      20615: inst = 32'hc40508b;
      20616: inst = 32'h8220000;
      20617: inst = 32'h10408000;
      20618: inst = 32'hc40508c;
      20619: inst = 32'h8220000;
      20620: inst = 32'h10408000;
      20621: inst = 32'hc40508d;
      20622: inst = 32'h8220000;
      20623: inst = 32'h10408000;
      20624: inst = 32'hc405090;
      20625: inst = 32'h8220000;
      20626: inst = 32'h10408000;
      20627: inst = 32'hc405091;
      20628: inst = 32'h8220000;
      20629: inst = 32'h10408000;
      20630: inst = 32'hc405096;
      20631: inst = 32'h8220000;
      20632: inst = 32'h10408000;
      20633: inst = 32'hc405097;
      20634: inst = 32'h8220000;
      20635: inst = 32'h10408000;
      20636: inst = 32'hc405098;
      20637: inst = 32'h8220000;
      20638: inst = 32'h10408000;
      20639: inst = 32'hc405099;
      20640: inst = 32'h8220000;
      20641: inst = 32'h10408000;
      20642: inst = 32'hc40509c;
      20643: inst = 32'h8220000;
      20644: inst = 32'h10408000;
      20645: inst = 32'hc40509d;
      20646: inst = 32'h8220000;
      20647: inst = 32'h10408000;
      20648: inst = 32'hc4050a9;
      20649: inst = 32'h8220000;
      20650: inst = 32'h10408000;
      20651: inst = 32'hc4050aa;
      20652: inst = 32'h8220000;
      20653: inst = 32'h10408000;
      20654: inst = 32'hc4050ab;
      20655: inst = 32'h8220000;
      20656: inst = 32'h10408000;
      20657: inst = 32'hc4050ac;
      20658: inst = 32'h8220000;
      20659: inst = 32'h10408000;
      20660: inst = 32'hc4050ad;
      20661: inst = 32'h8220000;
      20662: inst = 32'h10408000;
      20663: inst = 32'hc4050ae;
      20664: inst = 32'h8220000;
      20665: inst = 32'h10408000;
      20666: inst = 32'hc4050af;
      20667: inst = 32'h8220000;
      20668: inst = 32'h10408000;
      20669: inst = 32'hc4050b0;
      20670: inst = 32'h8220000;
      20671: inst = 32'h10408000;
      20672: inst = 32'hc4050b1;
      20673: inst = 32'h8220000;
      20674: inst = 32'h10408000;
      20675: inst = 32'hc4050b2;
      20676: inst = 32'h8220000;
      20677: inst = 32'h10408000;
      20678: inst = 32'hc4050b3;
      20679: inst = 32'h8220000;
      20680: inst = 32'h10408000;
      20681: inst = 32'hc4050cb;
      20682: inst = 32'h8220000;
      20683: inst = 32'h10408000;
      20684: inst = 32'hc4050cc;
      20685: inst = 32'h8220000;
      20686: inst = 32'h10408000;
      20687: inst = 32'hc4050cd;
      20688: inst = 32'h8220000;
      20689: inst = 32'h10408000;
      20690: inst = 32'hc4050ce;
      20691: inst = 32'h8220000;
      20692: inst = 32'h10408000;
      20693: inst = 32'hc4050cf;
      20694: inst = 32'h8220000;
      20695: inst = 32'h10408000;
      20696: inst = 32'hc4050d0;
      20697: inst = 32'h8220000;
      20698: inst = 32'h10408000;
      20699: inst = 32'hc4050d1;
      20700: inst = 32'h8220000;
      20701: inst = 32'h10408000;
      20702: inst = 32'hc4050d2;
      20703: inst = 32'h8220000;
      20704: inst = 32'h10408000;
      20705: inst = 32'hc4050d3;
      20706: inst = 32'h8220000;
      20707: inst = 32'h10408000;
      20708: inst = 32'hc4050d4;
      20709: inst = 32'h8220000;
      20710: inst = 32'h10408000;
      20711: inst = 32'hc4050d7;
      20712: inst = 32'h8220000;
      20713: inst = 32'h10408000;
      20714: inst = 32'hc4050d8;
      20715: inst = 32'h8220000;
      20716: inst = 32'h10408000;
      20717: inst = 32'hc4050d9;
      20718: inst = 32'h8220000;
      20719: inst = 32'h10408000;
      20720: inst = 32'hc4050da;
      20721: inst = 32'h8220000;
      20722: inst = 32'h10408000;
      20723: inst = 32'hc4050db;
      20724: inst = 32'h8220000;
      20725: inst = 32'h10408000;
      20726: inst = 32'hc4050dc;
      20727: inst = 32'h8220000;
      20728: inst = 32'h10408000;
      20729: inst = 32'hc4050dd;
      20730: inst = 32'h8220000;
      20731: inst = 32'h10408000;
      20732: inst = 32'hc4050de;
      20733: inst = 32'h8220000;
      20734: inst = 32'h10408000;
      20735: inst = 32'hc4050df;
      20736: inst = 32'h8220000;
      20737: inst = 32'h10408000;
      20738: inst = 32'hc4050e0;
      20739: inst = 32'h8220000;
      20740: inst = 32'h10408000;
      20741: inst = 32'hc4050e1;
      20742: inst = 32'h8220000;
      20743: inst = 32'h10408000;
      20744: inst = 32'hc4050e5;
      20745: inst = 32'h8220000;
      20746: inst = 32'h10408000;
      20747: inst = 32'hc4050e6;
      20748: inst = 32'h8220000;
      20749: inst = 32'h10408000;
      20750: inst = 32'hc4050e7;
      20751: inst = 32'h8220000;
      20752: inst = 32'h10408000;
      20753: inst = 32'hc4050e8;
      20754: inst = 32'h8220000;
      20755: inst = 32'h10408000;
      20756: inst = 32'hc4050e9;
      20757: inst = 32'h8220000;
      20758: inst = 32'h10408000;
      20759: inst = 32'hc4050ea;
      20760: inst = 32'h8220000;
      20761: inst = 32'h10408000;
      20762: inst = 32'hc4050eb;
      20763: inst = 32'h8220000;
      20764: inst = 32'h10408000;
      20765: inst = 32'hc4050ec;
      20766: inst = 32'h8220000;
      20767: inst = 32'h10408000;
      20768: inst = 32'hc4050ed;
      20769: inst = 32'h8220000;
      20770: inst = 32'h10408000;
      20771: inst = 32'hc4050f0;
      20772: inst = 32'h8220000;
      20773: inst = 32'h10408000;
      20774: inst = 32'hc4050f1;
      20775: inst = 32'h8220000;
      20776: inst = 32'h10408000;
      20777: inst = 32'hc4050f6;
      20778: inst = 32'h8220000;
      20779: inst = 32'h10408000;
      20780: inst = 32'hc4050f7;
      20781: inst = 32'h8220000;
      20782: inst = 32'h10408000;
      20783: inst = 32'hc4050f8;
      20784: inst = 32'h8220000;
      20785: inst = 32'h10408000;
      20786: inst = 32'hc4050f9;
      20787: inst = 32'h8220000;
      20788: inst = 32'h10408000;
      20789: inst = 32'hc4050fa;
      20790: inst = 32'h8220000;
      20791: inst = 32'h10408000;
      20792: inst = 32'hc4050fc;
      20793: inst = 32'h8220000;
      20794: inst = 32'h10408000;
      20795: inst = 32'hc4050fd;
      20796: inst = 32'h8220000;
      20797: inst = 32'h10408000;
      20798: inst = 32'hc405109;
      20799: inst = 32'h8220000;
      20800: inst = 32'h10408000;
      20801: inst = 32'hc40510a;
      20802: inst = 32'h8220000;
      20803: inst = 32'h10408000;
      20804: inst = 32'hc40510b;
      20805: inst = 32'h8220000;
      20806: inst = 32'h10408000;
      20807: inst = 32'hc40510c;
      20808: inst = 32'h8220000;
      20809: inst = 32'h10408000;
      20810: inst = 32'hc40510d;
      20811: inst = 32'h8220000;
      20812: inst = 32'h10408000;
      20813: inst = 32'hc40510e;
      20814: inst = 32'h8220000;
      20815: inst = 32'h10408000;
      20816: inst = 32'hc40510f;
      20817: inst = 32'h8220000;
      20818: inst = 32'h10408000;
      20819: inst = 32'hc405110;
      20820: inst = 32'h8220000;
      20821: inst = 32'h10408000;
      20822: inst = 32'hc405111;
      20823: inst = 32'h8220000;
      20824: inst = 32'h10408000;
      20825: inst = 32'hc405112;
      20826: inst = 32'h8220000;
      20827: inst = 32'h10408000;
      20828: inst = 32'hc405113;
      20829: inst = 32'h8220000;
      20830: inst = 32'h58000000;
      20831: inst = 32'h29c20000;
      20832: inst = 32'h29e30000;
      20833: inst = 32'h11600000;
      20834: inst = 32'hd600060;
      20835: inst = 32'h12208000;
      20836: inst = 32'he203fe0;
      20837: inst = 32'h13e00000;
      20838: inst = 32'hfe0517d;
      20839: inst = 32'h20200000;
      20840: inst = 32'h5be00000;
      20841: inst = 32'h13e00000;
      20842: inst = 32'hfe05d4c;
      20843: inst = 32'h20200001;
      20844: inst = 32'h5be00000;
      20845: inst = 32'h13e00000;
      20846: inst = 32'hfe05d4c;
      20847: inst = 32'h20200002;
      20848: inst = 32'h5be00000;
      20849: inst = 32'h13e00000;
      20850: inst = 32'hfe05972;
      20851: inst = 32'h20200003;
      20852: inst = 32'h5be00000;
      20853: inst = 32'h13e00000;
      20854: inst = 32'hfe05972;
      20855: inst = 32'h20200004;
      20856: inst = 32'h5be00000;
      20857: inst = 32'h13e00000;
      20858: inst = 32'hfe05582;
      20859: inst = 32'h20200005;
      20860: inst = 32'h5be00000;
      20861: inst = 32'hc6018c3;
      20862: inst = 32'h2a0e0000;
      20863: inst = 32'h294f0000;
      20864: inst = 32'h11200000;
      20865: inst = 32'hd205185;
      20866: inst = 32'h13e00000;
      20867: inst = 32'hfe0aa19;
      20868: inst = 32'h5be00000;
      20869: inst = 32'h244c8000;
      20870: inst = 32'h24428800;
      20871: inst = 32'h8620000;
      20872: inst = 32'h2a0e0001;
      20873: inst = 32'h294f0000;
      20874: inst = 32'h11200000;
      20875: inst = 32'hd20518f;
      20876: inst = 32'h13e00000;
      20877: inst = 32'hfe0aa19;
      20878: inst = 32'h5be00000;
      20879: inst = 32'h244c8000;
      20880: inst = 32'h24428800;
      20881: inst = 32'h8620000;
      20882: inst = 32'h2a0e0002;
      20883: inst = 32'h294f0000;
      20884: inst = 32'h11200000;
      20885: inst = 32'hd205199;
      20886: inst = 32'h13e00000;
      20887: inst = 32'hfe0aa19;
      20888: inst = 32'h5be00000;
      20889: inst = 32'h244c8000;
      20890: inst = 32'h24428800;
      20891: inst = 32'h8620000;
      20892: inst = 32'h2a0e0003;
      20893: inst = 32'h294f0000;
      20894: inst = 32'h11200000;
      20895: inst = 32'hd2051a3;
      20896: inst = 32'h13e00000;
      20897: inst = 32'hfe0aa19;
      20898: inst = 32'h5be00000;
      20899: inst = 32'h244c8000;
      20900: inst = 32'h24428800;
      20901: inst = 32'h8620000;
      20902: inst = 32'h2a0e0004;
      20903: inst = 32'h294f0000;
      20904: inst = 32'h11200000;
      20905: inst = 32'hd2051ad;
      20906: inst = 32'h13e00000;
      20907: inst = 32'hfe0aa19;
      20908: inst = 32'h5be00000;
      20909: inst = 32'h244c8000;
      20910: inst = 32'h24428800;
      20911: inst = 32'h8620000;
      20912: inst = 32'h2a0e0005;
      20913: inst = 32'h294f0000;
      20914: inst = 32'h11200000;
      20915: inst = 32'hd2051b7;
      20916: inst = 32'h13e00000;
      20917: inst = 32'hfe0aa19;
      20918: inst = 32'h5be00000;
      20919: inst = 32'h244c8000;
      20920: inst = 32'h24428800;
      20921: inst = 32'h8620000;
      20922: inst = 32'h2a0e0006;
      20923: inst = 32'h294f0000;
      20924: inst = 32'h11200000;
      20925: inst = 32'hd2051c1;
      20926: inst = 32'h13e00000;
      20927: inst = 32'hfe0aa19;
      20928: inst = 32'h5be00000;
      20929: inst = 32'h244c8000;
      20930: inst = 32'h24428800;
      20931: inst = 32'h8620000;
      20932: inst = 32'h2a0e0007;
      20933: inst = 32'h294f0000;
      20934: inst = 32'h11200000;
      20935: inst = 32'hd2051cb;
      20936: inst = 32'h13e00000;
      20937: inst = 32'hfe0aa19;
      20938: inst = 32'h5be00000;
      20939: inst = 32'h244c8000;
      20940: inst = 32'h24428800;
      20941: inst = 32'h8620000;
      20942: inst = 32'h2a0e0008;
      20943: inst = 32'h294f0000;
      20944: inst = 32'h11200000;
      20945: inst = 32'hd2051d5;
      20946: inst = 32'h13e00000;
      20947: inst = 32'hfe0aa19;
      20948: inst = 32'h5be00000;
      20949: inst = 32'h244c8000;
      20950: inst = 32'h24428800;
      20951: inst = 32'h8620000;
      20952: inst = 32'h2a0e0009;
      20953: inst = 32'h294f0000;
      20954: inst = 32'h11200000;
      20955: inst = 32'hd2051df;
      20956: inst = 32'h13e00000;
      20957: inst = 32'hfe0aa19;
      20958: inst = 32'h5be00000;
      20959: inst = 32'h244c8000;
      20960: inst = 32'h24428800;
      20961: inst = 32'h8620000;
      20962: inst = 32'h2a0e0000;
      20963: inst = 32'h294f0001;
      20964: inst = 32'h11200000;
      20965: inst = 32'hd2051e9;
      20966: inst = 32'h13e00000;
      20967: inst = 32'hfe0aa19;
      20968: inst = 32'h5be00000;
      20969: inst = 32'h244c8000;
      20970: inst = 32'h24428800;
      20971: inst = 32'h8620000;
      20972: inst = 32'h2a0e0001;
      20973: inst = 32'h294f0001;
      20974: inst = 32'h11200000;
      20975: inst = 32'hd2051f3;
      20976: inst = 32'h13e00000;
      20977: inst = 32'hfe0aa19;
      20978: inst = 32'h5be00000;
      20979: inst = 32'h244c8000;
      20980: inst = 32'h24428800;
      20981: inst = 32'h8620000;
      20982: inst = 32'h2a0e0002;
      20983: inst = 32'h294f0001;
      20984: inst = 32'h11200000;
      20985: inst = 32'hd2051fd;
      20986: inst = 32'h13e00000;
      20987: inst = 32'hfe0aa19;
      20988: inst = 32'h5be00000;
      20989: inst = 32'h244c8000;
      20990: inst = 32'h24428800;
      20991: inst = 32'h8620000;
      20992: inst = 32'h2a0e0003;
      20993: inst = 32'h294f0001;
      20994: inst = 32'h11200000;
      20995: inst = 32'hd205207;
      20996: inst = 32'h13e00000;
      20997: inst = 32'hfe0aa19;
      20998: inst = 32'h5be00000;
      20999: inst = 32'h244c8000;
      21000: inst = 32'h24428800;
      21001: inst = 32'h8620000;
      21002: inst = 32'h2a0e0004;
      21003: inst = 32'h294f0001;
      21004: inst = 32'h11200000;
      21005: inst = 32'hd205211;
      21006: inst = 32'h13e00000;
      21007: inst = 32'hfe0aa19;
      21008: inst = 32'h5be00000;
      21009: inst = 32'h244c8000;
      21010: inst = 32'h24428800;
      21011: inst = 32'h8620000;
      21012: inst = 32'h2a0e0005;
      21013: inst = 32'h294f0001;
      21014: inst = 32'h11200000;
      21015: inst = 32'hd20521b;
      21016: inst = 32'h13e00000;
      21017: inst = 32'hfe0aa19;
      21018: inst = 32'h5be00000;
      21019: inst = 32'h244c8000;
      21020: inst = 32'h24428800;
      21021: inst = 32'h8620000;
      21022: inst = 32'h2a0e0006;
      21023: inst = 32'h294f0001;
      21024: inst = 32'h11200000;
      21025: inst = 32'hd205225;
      21026: inst = 32'h13e00000;
      21027: inst = 32'hfe0aa19;
      21028: inst = 32'h5be00000;
      21029: inst = 32'h244c8000;
      21030: inst = 32'h24428800;
      21031: inst = 32'h8620000;
      21032: inst = 32'h2a0e0007;
      21033: inst = 32'h294f0001;
      21034: inst = 32'h11200000;
      21035: inst = 32'hd20522f;
      21036: inst = 32'h13e00000;
      21037: inst = 32'hfe0aa19;
      21038: inst = 32'h5be00000;
      21039: inst = 32'h244c8000;
      21040: inst = 32'h24428800;
      21041: inst = 32'h8620000;
      21042: inst = 32'h2a0e0008;
      21043: inst = 32'h294f0001;
      21044: inst = 32'h11200000;
      21045: inst = 32'hd205239;
      21046: inst = 32'h13e00000;
      21047: inst = 32'hfe0aa19;
      21048: inst = 32'h5be00000;
      21049: inst = 32'h244c8000;
      21050: inst = 32'h24428800;
      21051: inst = 32'h8620000;
      21052: inst = 32'h2a0e0009;
      21053: inst = 32'h294f0001;
      21054: inst = 32'h11200000;
      21055: inst = 32'hd205243;
      21056: inst = 32'h13e00000;
      21057: inst = 32'hfe0aa19;
      21058: inst = 32'h5be00000;
      21059: inst = 32'h244c8000;
      21060: inst = 32'h24428800;
      21061: inst = 32'h8620000;
      21062: inst = 32'h2a0e0000;
      21063: inst = 32'h294f0002;
      21064: inst = 32'h11200000;
      21065: inst = 32'hd20524d;
      21066: inst = 32'h13e00000;
      21067: inst = 32'hfe0aa19;
      21068: inst = 32'h5be00000;
      21069: inst = 32'h244c8000;
      21070: inst = 32'h24428800;
      21071: inst = 32'h8620000;
      21072: inst = 32'h2a0e0009;
      21073: inst = 32'h294f0002;
      21074: inst = 32'h11200000;
      21075: inst = 32'hd205257;
      21076: inst = 32'h13e00000;
      21077: inst = 32'hfe0aa19;
      21078: inst = 32'h5be00000;
      21079: inst = 32'h244c8000;
      21080: inst = 32'h24428800;
      21081: inst = 32'h8620000;
      21082: inst = 32'h2a0e0000;
      21083: inst = 32'h294f0003;
      21084: inst = 32'h11200000;
      21085: inst = 32'hd205261;
      21086: inst = 32'h13e00000;
      21087: inst = 32'hfe0aa19;
      21088: inst = 32'h5be00000;
      21089: inst = 32'h244c8000;
      21090: inst = 32'h24428800;
      21091: inst = 32'h8620000;
      21092: inst = 32'h2a0e0002;
      21093: inst = 32'h294f0003;
      21094: inst = 32'h11200000;
      21095: inst = 32'hd20526b;
      21096: inst = 32'h13e00000;
      21097: inst = 32'hfe0aa19;
      21098: inst = 32'h5be00000;
      21099: inst = 32'h244c8000;
      21100: inst = 32'h24428800;
      21101: inst = 32'h8620000;
      21102: inst = 32'h2a0e0007;
      21103: inst = 32'h294f0003;
      21104: inst = 32'h11200000;
      21105: inst = 32'hd205275;
      21106: inst = 32'h13e00000;
      21107: inst = 32'hfe0aa19;
      21108: inst = 32'h5be00000;
      21109: inst = 32'h244c8000;
      21110: inst = 32'h24428800;
      21111: inst = 32'h8620000;
      21112: inst = 32'h2a0e0009;
      21113: inst = 32'h294f0003;
      21114: inst = 32'h11200000;
      21115: inst = 32'hd20527f;
      21116: inst = 32'h13e00000;
      21117: inst = 32'hfe0aa19;
      21118: inst = 32'h5be00000;
      21119: inst = 32'h244c8000;
      21120: inst = 32'h24428800;
      21121: inst = 32'h8620000;
      21122: inst = 32'h2a0e0000;
      21123: inst = 32'h294f0004;
      21124: inst = 32'h11200000;
      21125: inst = 32'hd205289;
      21126: inst = 32'h13e00000;
      21127: inst = 32'hfe0aa19;
      21128: inst = 32'h5be00000;
      21129: inst = 32'h244c8000;
      21130: inst = 32'h24428800;
      21131: inst = 32'h8620000;
      21132: inst = 32'h2a0e0002;
      21133: inst = 32'h294f0004;
      21134: inst = 32'h11200000;
      21135: inst = 32'hd205293;
      21136: inst = 32'h13e00000;
      21137: inst = 32'hfe0aa19;
      21138: inst = 32'h5be00000;
      21139: inst = 32'h244c8000;
      21140: inst = 32'h24428800;
      21141: inst = 32'h8620000;
      21142: inst = 32'h2a0e0007;
      21143: inst = 32'h294f0004;
      21144: inst = 32'h11200000;
      21145: inst = 32'hd20529d;
      21146: inst = 32'h13e00000;
      21147: inst = 32'hfe0aa19;
      21148: inst = 32'h5be00000;
      21149: inst = 32'h244c8000;
      21150: inst = 32'h24428800;
      21151: inst = 32'h8620000;
      21152: inst = 32'h2a0e0009;
      21153: inst = 32'h294f0004;
      21154: inst = 32'h11200000;
      21155: inst = 32'hd2052a7;
      21156: inst = 32'h13e00000;
      21157: inst = 32'hfe0aa19;
      21158: inst = 32'h5be00000;
      21159: inst = 32'h244c8000;
      21160: inst = 32'h24428800;
      21161: inst = 32'h8620000;
      21162: inst = 32'h2a0e0000;
      21163: inst = 32'h294f0005;
      21164: inst = 32'h11200000;
      21165: inst = 32'hd2052b1;
      21166: inst = 32'h13e00000;
      21167: inst = 32'hfe0aa19;
      21168: inst = 32'h5be00000;
      21169: inst = 32'h244c8000;
      21170: inst = 32'h24428800;
      21171: inst = 32'h8620000;
      21172: inst = 32'h2a0e0009;
      21173: inst = 32'h294f0005;
      21174: inst = 32'h11200000;
      21175: inst = 32'hd2052bb;
      21176: inst = 32'h13e00000;
      21177: inst = 32'hfe0aa19;
      21178: inst = 32'h5be00000;
      21179: inst = 32'h244c8000;
      21180: inst = 32'h24428800;
      21181: inst = 32'h8620000;
      21182: inst = 32'h2a0e0000;
      21183: inst = 32'h294f0006;
      21184: inst = 32'h11200000;
      21185: inst = 32'hd2052c5;
      21186: inst = 32'h13e00000;
      21187: inst = 32'hfe0aa19;
      21188: inst = 32'h5be00000;
      21189: inst = 32'h244c8000;
      21190: inst = 32'h24428800;
      21191: inst = 32'h8620000;
      21192: inst = 32'h2a0e0009;
      21193: inst = 32'h294f0006;
      21194: inst = 32'h11200000;
      21195: inst = 32'hd2052cf;
      21196: inst = 32'h13e00000;
      21197: inst = 32'hfe0aa19;
      21198: inst = 32'h5be00000;
      21199: inst = 32'h244c8000;
      21200: inst = 32'h24428800;
      21201: inst = 32'h8620000;
      21202: inst = 32'hc60f4ce;
      21203: inst = 32'h2a0e0001;
      21204: inst = 32'h294f0002;
      21205: inst = 32'h11200000;
      21206: inst = 32'hd2052da;
      21207: inst = 32'h13e00000;
      21208: inst = 32'hfe0aa19;
      21209: inst = 32'h5be00000;
      21210: inst = 32'h244c8000;
      21211: inst = 32'h24428800;
      21212: inst = 32'h8620000;
      21213: inst = 32'h2a0e0002;
      21214: inst = 32'h294f0002;
      21215: inst = 32'h11200000;
      21216: inst = 32'hd2052e4;
      21217: inst = 32'h13e00000;
      21218: inst = 32'hfe0aa19;
      21219: inst = 32'h5be00000;
      21220: inst = 32'h244c8000;
      21221: inst = 32'h24428800;
      21222: inst = 32'h8620000;
      21223: inst = 32'h2a0e0003;
      21224: inst = 32'h294f0002;
      21225: inst = 32'h11200000;
      21226: inst = 32'hd2052ee;
      21227: inst = 32'h13e00000;
      21228: inst = 32'hfe0aa19;
      21229: inst = 32'h5be00000;
      21230: inst = 32'h244c8000;
      21231: inst = 32'h24428800;
      21232: inst = 32'h8620000;
      21233: inst = 32'h2a0e0004;
      21234: inst = 32'h294f0002;
      21235: inst = 32'h11200000;
      21236: inst = 32'hd2052f8;
      21237: inst = 32'h13e00000;
      21238: inst = 32'hfe0aa19;
      21239: inst = 32'h5be00000;
      21240: inst = 32'h244c8000;
      21241: inst = 32'h24428800;
      21242: inst = 32'h8620000;
      21243: inst = 32'h2a0e0005;
      21244: inst = 32'h294f0002;
      21245: inst = 32'h11200000;
      21246: inst = 32'hd205302;
      21247: inst = 32'h13e00000;
      21248: inst = 32'hfe0aa19;
      21249: inst = 32'h5be00000;
      21250: inst = 32'h244c8000;
      21251: inst = 32'h24428800;
      21252: inst = 32'h8620000;
      21253: inst = 32'h2a0e0006;
      21254: inst = 32'h294f0002;
      21255: inst = 32'h11200000;
      21256: inst = 32'hd20530c;
      21257: inst = 32'h13e00000;
      21258: inst = 32'hfe0aa19;
      21259: inst = 32'h5be00000;
      21260: inst = 32'h244c8000;
      21261: inst = 32'h24428800;
      21262: inst = 32'h8620000;
      21263: inst = 32'h2a0e0007;
      21264: inst = 32'h294f0002;
      21265: inst = 32'h11200000;
      21266: inst = 32'hd205316;
      21267: inst = 32'h13e00000;
      21268: inst = 32'hfe0aa19;
      21269: inst = 32'h5be00000;
      21270: inst = 32'h244c8000;
      21271: inst = 32'h24428800;
      21272: inst = 32'h8620000;
      21273: inst = 32'h2a0e0008;
      21274: inst = 32'h294f0002;
      21275: inst = 32'h11200000;
      21276: inst = 32'hd205320;
      21277: inst = 32'h13e00000;
      21278: inst = 32'hfe0aa19;
      21279: inst = 32'h5be00000;
      21280: inst = 32'h244c8000;
      21281: inst = 32'h24428800;
      21282: inst = 32'h8620000;
      21283: inst = 32'h2a0e0001;
      21284: inst = 32'h294f0003;
      21285: inst = 32'h11200000;
      21286: inst = 32'hd20532a;
      21287: inst = 32'h13e00000;
      21288: inst = 32'hfe0aa19;
      21289: inst = 32'h5be00000;
      21290: inst = 32'h244c8000;
      21291: inst = 32'h24428800;
      21292: inst = 32'h8620000;
      21293: inst = 32'h2a0e0003;
      21294: inst = 32'h294f0003;
      21295: inst = 32'h11200000;
      21296: inst = 32'hd205334;
      21297: inst = 32'h13e00000;
      21298: inst = 32'hfe0aa19;
      21299: inst = 32'h5be00000;
      21300: inst = 32'h244c8000;
      21301: inst = 32'h24428800;
      21302: inst = 32'h8620000;
      21303: inst = 32'h2a0e0004;
      21304: inst = 32'h294f0003;
      21305: inst = 32'h11200000;
      21306: inst = 32'hd20533e;
      21307: inst = 32'h13e00000;
      21308: inst = 32'hfe0aa19;
      21309: inst = 32'h5be00000;
      21310: inst = 32'h244c8000;
      21311: inst = 32'h24428800;
      21312: inst = 32'h8620000;
      21313: inst = 32'h2a0e0005;
      21314: inst = 32'h294f0003;
      21315: inst = 32'h11200000;
      21316: inst = 32'hd205348;
      21317: inst = 32'h13e00000;
      21318: inst = 32'hfe0aa19;
      21319: inst = 32'h5be00000;
      21320: inst = 32'h244c8000;
      21321: inst = 32'h24428800;
      21322: inst = 32'h8620000;
      21323: inst = 32'h2a0e0006;
      21324: inst = 32'h294f0003;
      21325: inst = 32'h11200000;
      21326: inst = 32'hd205352;
      21327: inst = 32'h13e00000;
      21328: inst = 32'hfe0aa19;
      21329: inst = 32'h5be00000;
      21330: inst = 32'h244c8000;
      21331: inst = 32'h24428800;
      21332: inst = 32'h8620000;
      21333: inst = 32'h2a0e0008;
      21334: inst = 32'h294f0003;
      21335: inst = 32'h11200000;
      21336: inst = 32'hd20535c;
      21337: inst = 32'h13e00000;
      21338: inst = 32'hfe0aa19;
      21339: inst = 32'h5be00000;
      21340: inst = 32'h244c8000;
      21341: inst = 32'h24428800;
      21342: inst = 32'h8620000;
      21343: inst = 32'h2a0e0001;
      21344: inst = 32'h294f0004;
      21345: inst = 32'h11200000;
      21346: inst = 32'hd205366;
      21347: inst = 32'h13e00000;
      21348: inst = 32'hfe0aa19;
      21349: inst = 32'h5be00000;
      21350: inst = 32'h244c8000;
      21351: inst = 32'h24428800;
      21352: inst = 32'h8620000;
      21353: inst = 32'h2a0e0003;
      21354: inst = 32'h294f0004;
      21355: inst = 32'h11200000;
      21356: inst = 32'hd205370;
      21357: inst = 32'h13e00000;
      21358: inst = 32'hfe0aa19;
      21359: inst = 32'h5be00000;
      21360: inst = 32'h244c8000;
      21361: inst = 32'h24428800;
      21362: inst = 32'h8620000;
      21363: inst = 32'h2a0e0004;
      21364: inst = 32'h294f0004;
      21365: inst = 32'h11200000;
      21366: inst = 32'hd20537a;
      21367: inst = 32'h13e00000;
      21368: inst = 32'hfe0aa19;
      21369: inst = 32'h5be00000;
      21370: inst = 32'h244c8000;
      21371: inst = 32'h24428800;
      21372: inst = 32'h8620000;
      21373: inst = 32'h2a0e0005;
      21374: inst = 32'h294f0004;
      21375: inst = 32'h11200000;
      21376: inst = 32'hd205384;
      21377: inst = 32'h13e00000;
      21378: inst = 32'hfe0aa19;
      21379: inst = 32'h5be00000;
      21380: inst = 32'h244c8000;
      21381: inst = 32'h24428800;
      21382: inst = 32'h8620000;
      21383: inst = 32'h2a0e0006;
      21384: inst = 32'h294f0004;
      21385: inst = 32'h11200000;
      21386: inst = 32'hd20538e;
      21387: inst = 32'h13e00000;
      21388: inst = 32'hfe0aa19;
      21389: inst = 32'h5be00000;
      21390: inst = 32'h244c8000;
      21391: inst = 32'h24428800;
      21392: inst = 32'h8620000;
      21393: inst = 32'h2a0e0008;
      21394: inst = 32'h294f0004;
      21395: inst = 32'h11200000;
      21396: inst = 32'hd205398;
      21397: inst = 32'h13e00000;
      21398: inst = 32'hfe0aa19;
      21399: inst = 32'h5be00000;
      21400: inst = 32'h244c8000;
      21401: inst = 32'h24428800;
      21402: inst = 32'h8620000;
      21403: inst = 32'h2a0e0001;
      21404: inst = 32'h294f0005;
      21405: inst = 32'h11200000;
      21406: inst = 32'hd2053a2;
      21407: inst = 32'h13e00000;
      21408: inst = 32'hfe0aa19;
      21409: inst = 32'h5be00000;
      21410: inst = 32'h244c8000;
      21411: inst = 32'h24428800;
      21412: inst = 32'h8620000;
      21413: inst = 32'h2a0e0002;
      21414: inst = 32'h294f0005;
      21415: inst = 32'h11200000;
      21416: inst = 32'hd2053ac;
      21417: inst = 32'h13e00000;
      21418: inst = 32'hfe0aa19;
      21419: inst = 32'h5be00000;
      21420: inst = 32'h244c8000;
      21421: inst = 32'h24428800;
      21422: inst = 32'h8620000;
      21423: inst = 32'h2a0e0003;
      21424: inst = 32'h294f0005;
      21425: inst = 32'h11200000;
      21426: inst = 32'hd2053b6;
      21427: inst = 32'h13e00000;
      21428: inst = 32'hfe0aa19;
      21429: inst = 32'h5be00000;
      21430: inst = 32'h244c8000;
      21431: inst = 32'h24428800;
      21432: inst = 32'h8620000;
      21433: inst = 32'h2a0e0004;
      21434: inst = 32'h294f0005;
      21435: inst = 32'h11200000;
      21436: inst = 32'hd2053c0;
      21437: inst = 32'h13e00000;
      21438: inst = 32'hfe0aa19;
      21439: inst = 32'h5be00000;
      21440: inst = 32'h244c8000;
      21441: inst = 32'h24428800;
      21442: inst = 32'h8620000;
      21443: inst = 32'h2a0e0005;
      21444: inst = 32'h294f0005;
      21445: inst = 32'h11200000;
      21446: inst = 32'hd2053ca;
      21447: inst = 32'h13e00000;
      21448: inst = 32'hfe0aa19;
      21449: inst = 32'h5be00000;
      21450: inst = 32'h244c8000;
      21451: inst = 32'h24428800;
      21452: inst = 32'h8620000;
      21453: inst = 32'h2a0e0006;
      21454: inst = 32'h294f0005;
      21455: inst = 32'h11200000;
      21456: inst = 32'hd2053d4;
      21457: inst = 32'h13e00000;
      21458: inst = 32'hfe0aa19;
      21459: inst = 32'h5be00000;
      21460: inst = 32'h244c8000;
      21461: inst = 32'h24428800;
      21462: inst = 32'h8620000;
      21463: inst = 32'h2a0e0007;
      21464: inst = 32'h294f0005;
      21465: inst = 32'h11200000;
      21466: inst = 32'hd2053de;
      21467: inst = 32'h13e00000;
      21468: inst = 32'hfe0aa19;
      21469: inst = 32'h5be00000;
      21470: inst = 32'h244c8000;
      21471: inst = 32'h24428800;
      21472: inst = 32'h8620000;
      21473: inst = 32'h2a0e0008;
      21474: inst = 32'h294f0005;
      21475: inst = 32'h11200000;
      21476: inst = 32'hd2053e8;
      21477: inst = 32'h13e00000;
      21478: inst = 32'hfe0aa19;
      21479: inst = 32'h5be00000;
      21480: inst = 32'h244c8000;
      21481: inst = 32'h24428800;
      21482: inst = 32'h8620000;
      21483: inst = 32'h2a0e0001;
      21484: inst = 32'h294f0006;
      21485: inst = 32'h11200000;
      21486: inst = 32'hd2053f2;
      21487: inst = 32'h13e00000;
      21488: inst = 32'hfe0aa19;
      21489: inst = 32'h5be00000;
      21490: inst = 32'h244c8000;
      21491: inst = 32'h24428800;
      21492: inst = 32'h8620000;
      21493: inst = 32'h2a0e0002;
      21494: inst = 32'h294f0006;
      21495: inst = 32'h11200000;
      21496: inst = 32'hd2053fc;
      21497: inst = 32'h13e00000;
      21498: inst = 32'hfe0aa19;
      21499: inst = 32'h5be00000;
      21500: inst = 32'h244c8000;
      21501: inst = 32'h24428800;
      21502: inst = 32'h8620000;
      21503: inst = 32'h2a0e0003;
      21504: inst = 32'h294f0006;
      21505: inst = 32'h11200000;
      21506: inst = 32'hd205406;
      21507: inst = 32'h13e00000;
      21508: inst = 32'hfe0aa19;
      21509: inst = 32'h5be00000;
      21510: inst = 32'h244c8000;
      21511: inst = 32'h24428800;
      21512: inst = 32'h8620000;
      21513: inst = 32'h2a0e0004;
      21514: inst = 32'h294f0006;
      21515: inst = 32'h11200000;
      21516: inst = 32'hd205410;
      21517: inst = 32'h13e00000;
      21518: inst = 32'hfe0aa19;
      21519: inst = 32'h5be00000;
      21520: inst = 32'h244c8000;
      21521: inst = 32'h24428800;
      21522: inst = 32'h8620000;
      21523: inst = 32'h2a0e0005;
      21524: inst = 32'h294f0006;
      21525: inst = 32'h11200000;
      21526: inst = 32'hd20541a;
      21527: inst = 32'h13e00000;
      21528: inst = 32'hfe0aa19;
      21529: inst = 32'h5be00000;
      21530: inst = 32'h244c8000;
      21531: inst = 32'h24428800;
      21532: inst = 32'h8620000;
      21533: inst = 32'h2a0e0006;
      21534: inst = 32'h294f0006;
      21535: inst = 32'h11200000;
      21536: inst = 32'hd205424;
      21537: inst = 32'h13e00000;
      21538: inst = 32'hfe0aa19;
      21539: inst = 32'h5be00000;
      21540: inst = 32'h244c8000;
      21541: inst = 32'h24428800;
      21542: inst = 32'h8620000;
      21543: inst = 32'h2a0e0007;
      21544: inst = 32'h294f0006;
      21545: inst = 32'h11200000;
      21546: inst = 32'hd20542e;
      21547: inst = 32'h13e00000;
      21548: inst = 32'hfe0aa19;
      21549: inst = 32'h5be00000;
      21550: inst = 32'h244c8000;
      21551: inst = 32'h24428800;
      21552: inst = 32'h8620000;
      21553: inst = 32'h2a0e0008;
      21554: inst = 32'h294f0006;
      21555: inst = 32'h11200000;
      21556: inst = 32'hd205438;
      21557: inst = 32'h13e00000;
      21558: inst = 32'hfe0aa19;
      21559: inst = 32'h5be00000;
      21560: inst = 32'h244c8000;
      21561: inst = 32'h24428800;
      21562: inst = 32'h8620000;
      21563: inst = 32'h2a0e0000;
      21564: inst = 32'h294f0008;
      21565: inst = 32'h11200000;
      21566: inst = 32'hd205442;
      21567: inst = 32'h13e00000;
      21568: inst = 32'hfe0aa19;
      21569: inst = 32'h5be00000;
      21570: inst = 32'h244c8000;
      21571: inst = 32'h24428800;
      21572: inst = 32'h8620000;
      21573: inst = 32'h2a0e0001;
      21574: inst = 32'h294f0008;
      21575: inst = 32'h11200000;
      21576: inst = 32'hd20544c;
      21577: inst = 32'h13e00000;
      21578: inst = 32'hfe0aa19;
      21579: inst = 32'h5be00000;
      21580: inst = 32'h244c8000;
      21581: inst = 32'h24428800;
      21582: inst = 32'h8620000;
      21583: inst = 32'h2a0e0008;
      21584: inst = 32'h294f0008;
      21585: inst = 32'h11200000;
      21586: inst = 32'hd205456;
      21587: inst = 32'h13e00000;
      21588: inst = 32'hfe0aa19;
      21589: inst = 32'h5be00000;
      21590: inst = 32'h244c8000;
      21591: inst = 32'h24428800;
      21592: inst = 32'h8620000;
      21593: inst = 32'h2a0e0009;
      21594: inst = 32'h294f0008;
      21595: inst = 32'h11200000;
      21596: inst = 32'hd205460;
      21597: inst = 32'h13e00000;
      21598: inst = 32'hfe0aa19;
      21599: inst = 32'h5be00000;
      21600: inst = 32'h244c8000;
      21601: inst = 32'h24428800;
      21602: inst = 32'h8620000;
      21603: inst = 32'h2a0e0003;
      21604: inst = 32'h294f000c;
      21605: inst = 32'h11200000;
      21606: inst = 32'hd20546a;
      21607: inst = 32'h13e00000;
      21608: inst = 32'hfe0aa19;
      21609: inst = 32'h5be00000;
      21610: inst = 32'h244c8000;
      21611: inst = 32'h24428800;
      21612: inst = 32'h8620000;
      21613: inst = 32'h2a0e0006;
      21614: inst = 32'h294f000c;
      21615: inst = 32'h11200000;
      21616: inst = 32'hd205474;
      21617: inst = 32'h13e00000;
      21618: inst = 32'hfe0aa19;
      21619: inst = 32'h5be00000;
      21620: inst = 32'h244c8000;
      21621: inst = 32'h24428800;
      21622: inst = 32'h8620000;
      21623: inst = 32'hc607800;
      21624: inst = 32'h2a0e0002;
      21625: inst = 32'h294f0007;
      21626: inst = 32'h11200000;
      21627: inst = 32'hd20547f;
      21628: inst = 32'h13e00000;
      21629: inst = 32'hfe0aa19;
      21630: inst = 32'h5be00000;
      21631: inst = 32'h244c8000;
      21632: inst = 32'h24428800;
      21633: inst = 32'h8620000;
      21634: inst = 32'h2a0e0003;
      21635: inst = 32'h294f0007;
      21636: inst = 32'h11200000;
      21637: inst = 32'hd205489;
      21638: inst = 32'h13e00000;
      21639: inst = 32'hfe0aa19;
      21640: inst = 32'h5be00000;
      21641: inst = 32'h244c8000;
      21642: inst = 32'h24428800;
      21643: inst = 32'h8620000;
      21644: inst = 32'h2a0e0006;
      21645: inst = 32'h294f0007;
      21646: inst = 32'h11200000;
      21647: inst = 32'hd205493;
      21648: inst = 32'h13e00000;
      21649: inst = 32'hfe0aa19;
      21650: inst = 32'h5be00000;
      21651: inst = 32'h244c8000;
      21652: inst = 32'h24428800;
      21653: inst = 32'h8620000;
      21654: inst = 32'h2a0e0007;
      21655: inst = 32'h294f0007;
      21656: inst = 32'h11200000;
      21657: inst = 32'hd20549d;
      21658: inst = 32'h13e00000;
      21659: inst = 32'hfe0aa19;
      21660: inst = 32'h5be00000;
      21661: inst = 32'h244c8000;
      21662: inst = 32'h24428800;
      21663: inst = 32'h8620000;
      21664: inst = 32'hc60a000;
      21665: inst = 32'h2a0e0004;
      21666: inst = 32'h294f0007;
      21667: inst = 32'h11200000;
      21668: inst = 32'hd2054a8;
      21669: inst = 32'h13e00000;
      21670: inst = 32'hfe0aa19;
      21671: inst = 32'h5be00000;
      21672: inst = 32'h244c8000;
      21673: inst = 32'h24428800;
      21674: inst = 32'h8620000;
      21675: inst = 32'h2a0e0005;
      21676: inst = 32'h294f0007;
      21677: inst = 32'h11200000;
      21678: inst = 32'hd2054b2;
      21679: inst = 32'h13e00000;
      21680: inst = 32'hfe0aa19;
      21681: inst = 32'h5be00000;
      21682: inst = 32'h244c8000;
      21683: inst = 32'h24428800;
      21684: inst = 32'h8620000;
      21685: inst = 32'h2a0e0002;
      21686: inst = 32'h294f0008;
      21687: inst = 32'h11200000;
      21688: inst = 32'hd2054bc;
      21689: inst = 32'h13e00000;
      21690: inst = 32'hfe0aa19;
      21691: inst = 32'h5be00000;
      21692: inst = 32'h244c8000;
      21693: inst = 32'h24428800;
      21694: inst = 32'h8620000;
      21695: inst = 32'h2a0e0003;
      21696: inst = 32'h294f0008;
      21697: inst = 32'h11200000;
      21698: inst = 32'hd2054c6;
      21699: inst = 32'h13e00000;
      21700: inst = 32'hfe0aa19;
      21701: inst = 32'h5be00000;
      21702: inst = 32'h244c8000;
      21703: inst = 32'h24428800;
      21704: inst = 32'h8620000;
      21705: inst = 32'h2a0e0004;
      21706: inst = 32'h294f0008;
      21707: inst = 32'h11200000;
      21708: inst = 32'hd2054d0;
      21709: inst = 32'h13e00000;
      21710: inst = 32'hfe0aa19;
      21711: inst = 32'h5be00000;
      21712: inst = 32'h244c8000;
      21713: inst = 32'h24428800;
      21714: inst = 32'h8620000;
      21715: inst = 32'h2a0e0005;
      21716: inst = 32'h294f0008;
      21717: inst = 32'h11200000;
      21718: inst = 32'hd2054da;
      21719: inst = 32'h13e00000;
      21720: inst = 32'hfe0aa19;
      21721: inst = 32'h5be00000;
      21722: inst = 32'h244c8000;
      21723: inst = 32'h24428800;
      21724: inst = 32'h8620000;
      21725: inst = 32'h2a0e0006;
      21726: inst = 32'h294f0008;
      21727: inst = 32'h11200000;
      21728: inst = 32'hd2054e4;
      21729: inst = 32'h13e00000;
      21730: inst = 32'hfe0aa19;
      21731: inst = 32'h5be00000;
      21732: inst = 32'h244c8000;
      21733: inst = 32'h24428800;
      21734: inst = 32'h8620000;
      21735: inst = 32'h2a0e0007;
      21736: inst = 32'h294f0008;
      21737: inst = 32'h11200000;
      21738: inst = 32'hd2054ee;
      21739: inst = 32'h13e00000;
      21740: inst = 32'hfe0aa19;
      21741: inst = 32'h5be00000;
      21742: inst = 32'h244c8000;
      21743: inst = 32'h24428800;
      21744: inst = 32'h8620000;
      21745: inst = 32'h2a0e0002;
      21746: inst = 32'h294f0009;
      21747: inst = 32'h11200000;
      21748: inst = 32'hd2054f8;
      21749: inst = 32'h13e00000;
      21750: inst = 32'hfe0aa19;
      21751: inst = 32'h5be00000;
      21752: inst = 32'h244c8000;
      21753: inst = 32'h24428800;
      21754: inst = 32'h8620000;
      21755: inst = 32'h2a0e0003;
      21756: inst = 32'h294f0009;
      21757: inst = 32'h11200000;
      21758: inst = 32'hd205502;
      21759: inst = 32'h13e00000;
      21760: inst = 32'hfe0aa19;
      21761: inst = 32'h5be00000;
      21762: inst = 32'h244c8000;
      21763: inst = 32'h24428800;
      21764: inst = 32'h8620000;
      21765: inst = 32'h2a0e0004;
      21766: inst = 32'h294f0009;
      21767: inst = 32'h11200000;
      21768: inst = 32'hd20550c;
      21769: inst = 32'h13e00000;
      21770: inst = 32'hfe0aa19;
      21771: inst = 32'h5be00000;
      21772: inst = 32'h244c8000;
      21773: inst = 32'h24428800;
      21774: inst = 32'h8620000;
      21775: inst = 32'h2a0e0005;
      21776: inst = 32'h294f0009;
      21777: inst = 32'h11200000;
      21778: inst = 32'hd205516;
      21779: inst = 32'h13e00000;
      21780: inst = 32'hfe0aa19;
      21781: inst = 32'h5be00000;
      21782: inst = 32'h244c8000;
      21783: inst = 32'h24428800;
      21784: inst = 32'h8620000;
      21785: inst = 32'h2a0e0006;
      21786: inst = 32'h294f0009;
      21787: inst = 32'h11200000;
      21788: inst = 32'hd205520;
      21789: inst = 32'h13e00000;
      21790: inst = 32'hfe0aa19;
      21791: inst = 32'h5be00000;
      21792: inst = 32'h244c8000;
      21793: inst = 32'h24428800;
      21794: inst = 32'h8620000;
      21795: inst = 32'h2a0e0007;
      21796: inst = 32'h294f0009;
      21797: inst = 32'h11200000;
      21798: inst = 32'hd20552a;
      21799: inst = 32'h13e00000;
      21800: inst = 32'hfe0aa19;
      21801: inst = 32'h5be00000;
      21802: inst = 32'h244c8000;
      21803: inst = 32'h24428800;
      21804: inst = 32'h8620000;
      21805: inst = 32'hc6010ac;
      21806: inst = 32'h2a0e0002;
      21807: inst = 32'h294f000a;
      21808: inst = 32'h11200000;
      21809: inst = 32'hd205535;
      21810: inst = 32'h13e00000;
      21811: inst = 32'hfe0aa19;
      21812: inst = 32'h5be00000;
      21813: inst = 32'h244c8000;
      21814: inst = 32'h24428800;
      21815: inst = 32'h8620000;
      21816: inst = 32'h2a0e0003;
      21817: inst = 32'h294f000a;
      21818: inst = 32'h11200000;
      21819: inst = 32'hd20553f;
      21820: inst = 32'h13e00000;
      21821: inst = 32'hfe0aa19;
      21822: inst = 32'h5be00000;
      21823: inst = 32'h244c8000;
      21824: inst = 32'h24428800;
      21825: inst = 32'h8620000;
      21826: inst = 32'h2a0e0004;
      21827: inst = 32'h294f000a;
      21828: inst = 32'h11200000;
      21829: inst = 32'hd205549;
      21830: inst = 32'h13e00000;
      21831: inst = 32'hfe0aa19;
      21832: inst = 32'h5be00000;
      21833: inst = 32'h244c8000;
      21834: inst = 32'h24428800;
      21835: inst = 32'h8620000;
      21836: inst = 32'h2a0e0005;
      21837: inst = 32'h294f000a;
      21838: inst = 32'h11200000;
      21839: inst = 32'hd205553;
      21840: inst = 32'h13e00000;
      21841: inst = 32'hfe0aa19;
      21842: inst = 32'h5be00000;
      21843: inst = 32'h244c8000;
      21844: inst = 32'h24428800;
      21845: inst = 32'h8620000;
      21846: inst = 32'h2a0e0006;
      21847: inst = 32'h294f000a;
      21848: inst = 32'h11200000;
      21849: inst = 32'hd20555d;
      21850: inst = 32'h13e00000;
      21851: inst = 32'hfe0aa19;
      21852: inst = 32'h5be00000;
      21853: inst = 32'h244c8000;
      21854: inst = 32'h24428800;
      21855: inst = 32'h8620000;
      21856: inst = 32'h2a0e0007;
      21857: inst = 32'h294f000a;
      21858: inst = 32'h11200000;
      21859: inst = 32'hd205567;
      21860: inst = 32'h13e00000;
      21861: inst = 32'hfe0aa19;
      21862: inst = 32'h5be00000;
      21863: inst = 32'h244c8000;
      21864: inst = 32'h24428800;
      21865: inst = 32'h8620000;
      21866: inst = 32'hc60d42c;
      21867: inst = 32'h2a0e0003;
      21868: inst = 32'h294f000b;
      21869: inst = 32'h11200000;
      21870: inst = 32'hd205572;
      21871: inst = 32'h13e00000;
      21872: inst = 32'hfe0aa19;
      21873: inst = 32'h5be00000;
      21874: inst = 32'h244c8000;
      21875: inst = 32'h24428800;
      21876: inst = 32'h8620000;
      21877: inst = 32'h2a0e0006;
      21878: inst = 32'h294f000b;
      21879: inst = 32'h11200000;
      21880: inst = 32'hd20557c;
      21881: inst = 32'h13e00000;
      21882: inst = 32'hfe0aa19;
      21883: inst = 32'h5be00000;
      21884: inst = 32'h244c8000;
      21885: inst = 32'h24428800;
      21886: inst = 32'h8620000;
      21887: inst = 32'h13e00000;
      21888: inst = 32'hfe06126;
      21889: inst = 32'h5be00000;
      21890: inst = 32'hc6018c3;
      21891: inst = 32'h2a0e0000;
      21892: inst = 32'h294f0000;
      21893: inst = 32'h11200000;
      21894: inst = 32'hd20558a;
      21895: inst = 32'h13e00000;
      21896: inst = 32'hfe0aa19;
      21897: inst = 32'h5be00000;
      21898: inst = 32'h244c8000;
      21899: inst = 32'h24428800;
      21900: inst = 32'h8620000;
      21901: inst = 32'h2a0e0001;
      21902: inst = 32'h294f0000;
      21903: inst = 32'h11200000;
      21904: inst = 32'hd205594;
      21905: inst = 32'h13e00000;
      21906: inst = 32'hfe0aa19;
      21907: inst = 32'h5be00000;
      21908: inst = 32'h244c8000;
      21909: inst = 32'h24428800;
      21910: inst = 32'h8620000;
      21911: inst = 32'h2a0e0002;
      21912: inst = 32'h294f0000;
      21913: inst = 32'h11200000;
      21914: inst = 32'hd20559e;
      21915: inst = 32'h13e00000;
      21916: inst = 32'hfe0aa19;
      21917: inst = 32'h5be00000;
      21918: inst = 32'h244c8000;
      21919: inst = 32'h24428800;
      21920: inst = 32'h8620000;
      21921: inst = 32'h2a0e0003;
      21922: inst = 32'h294f0000;
      21923: inst = 32'h11200000;
      21924: inst = 32'hd2055a8;
      21925: inst = 32'h13e00000;
      21926: inst = 32'hfe0aa19;
      21927: inst = 32'h5be00000;
      21928: inst = 32'h244c8000;
      21929: inst = 32'h24428800;
      21930: inst = 32'h8620000;
      21931: inst = 32'h2a0e0004;
      21932: inst = 32'h294f0000;
      21933: inst = 32'h11200000;
      21934: inst = 32'hd2055b2;
      21935: inst = 32'h13e00000;
      21936: inst = 32'hfe0aa19;
      21937: inst = 32'h5be00000;
      21938: inst = 32'h244c8000;
      21939: inst = 32'h24428800;
      21940: inst = 32'h8620000;
      21941: inst = 32'h2a0e0005;
      21942: inst = 32'h294f0000;
      21943: inst = 32'h11200000;
      21944: inst = 32'hd2055bc;
      21945: inst = 32'h13e00000;
      21946: inst = 32'hfe0aa19;
      21947: inst = 32'h5be00000;
      21948: inst = 32'h244c8000;
      21949: inst = 32'h24428800;
      21950: inst = 32'h8620000;
      21951: inst = 32'h2a0e0006;
      21952: inst = 32'h294f0000;
      21953: inst = 32'h11200000;
      21954: inst = 32'hd2055c6;
      21955: inst = 32'h13e00000;
      21956: inst = 32'hfe0aa19;
      21957: inst = 32'h5be00000;
      21958: inst = 32'h244c8000;
      21959: inst = 32'h24428800;
      21960: inst = 32'h8620000;
      21961: inst = 32'h2a0e0007;
      21962: inst = 32'h294f0000;
      21963: inst = 32'h11200000;
      21964: inst = 32'hd2055d0;
      21965: inst = 32'h13e00000;
      21966: inst = 32'hfe0aa19;
      21967: inst = 32'h5be00000;
      21968: inst = 32'h244c8000;
      21969: inst = 32'h24428800;
      21970: inst = 32'h8620000;
      21971: inst = 32'h2a0e0008;
      21972: inst = 32'h294f0000;
      21973: inst = 32'h11200000;
      21974: inst = 32'hd2055da;
      21975: inst = 32'h13e00000;
      21976: inst = 32'hfe0aa19;
      21977: inst = 32'h5be00000;
      21978: inst = 32'h244c8000;
      21979: inst = 32'h24428800;
      21980: inst = 32'h8620000;
      21981: inst = 32'h2a0e0009;
      21982: inst = 32'h294f0000;
      21983: inst = 32'h11200000;
      21984: inst = 32'hd2055e4;
      21985: inst = 32'h13e00000;
      21986: inst = 32'hfe0aa19;
      21987: inst = 32'h5be00000;
      21988: inst = 32'h244c8000;
      21989: inst = 32'h24428800;
      21990: inst = 32'h8620000;
      21991: inst = 32'h2a0e0000;
      21992: inst = 32'h294f0001;
      21993: inst = 32'h11200000;
      21994: inst = 32'hd2055ee;
      21995: inst = 32'h13e00000;
      21996: inst = 32'hfe0aa19;
      21997: inst = 32'h5be00000;
      21998: inst = 32'h244c8000;
      21999: inst = 32'h24428800;
      22000: inst = 32'h8620000;
      22001: inst = 32'h2a0e0001;
      22002: inst = 32'h294f0001;
      22003: inst = 32'h11200000;
      22004: inst = 32'hd2055f8;
      22005: inst = 32'h13e00000;
      22006: inst = 32'hfe0aa19;
      22007: inst = 32'h5be00000;
      22008: inst = 32'h244c8000;
      22009: inst = 32'h24428800;
      22010: inst = 32'h8620000;
      22011: inst = 32'h2a0e0002;
      22012: inst = 32'h294f0001;
      22013: inst = 32'h11200000;
      22014: inst = 32'hd205602;
      22015: inst = 32'h13e00000;
      22016: inst = 32'hfe0aa19;
      22017: inst = 32'h5be00000;
      22018: inst = 32'h244c8000;
      22019: inst = 32'h24428800;
      22020: inst = 32'h8620000;
      22021: inst = 32'h2a0e0003;
      22022: inst = 32'h294f0001;
      22023: inst = 32'h11200000;
      22024: inst = 32'hd20560c;
      22025: inst = 32'h13e00000;
      22026: inst = 32'hfe0aa19;
      22027: inst = 32'h5be00000;
      22028: inst = 32'h244c8000;
      22029: inst = 32'h24428800;
      22030: inst = 32'h8620000;
      22031: inst = 32'h2a0e0004;
      22032: inst = 32'h294f0001;
      22033: inst = 32'h11200000;
      22034: inst = 32'hd205616;
      22035: inst = 32'h13e00000;
      22036: inst = 32'hfe0aa19;
      22037: inst = 32'h5be00000;
      22038: inst = 32'h244c8000;
      22039: inst = 32'h24428800;
      22040: inst = 32'h8620000;
      22041: inst = 32'h2a0e0005;
      22042: inst = 32'h294f0001;
      22043: inst = 32'h11200000;
      22044: inst = 32'hd205620;
      22045: inst = 32'h13e00000;
      22046: inst = 32'hfe0aa19;
      22047: inst = 32'h5be00000;
      22048: inst = 32'h244c8000;
      22049: inst = 32'h24428800;
      22050: inst = 32'h8620000;
      22051: inst = 32'h2a0e0006;
      22052: inst = 32'h294f0001;
      22053: inst = 32'h11200000;
      22054: inst = 32'hd20562a;
      22055: inst = 32'h13e00000;
      22056: inst = 32'hfe0aa19;
      22057: inst = 32'h5be00000;
      22058: inst = 32'h244c8000;
      22059: inst = 32'h24428800;
      22060: inst = 32'h8620000;
      22061: inst = 32'h2a0e0007;
      22062: inst = 32'h294f0001;
      22063: inst = 32'h11200000;
      22064: inst = 32'hd205634;
      22065: inst = 32'h13e00000;
      22066: inst = 32'hfe0aa19;
      22067: inst = 32'h5be00000;
      22068: inst = 32'h244c8000;
      22069: inst = 32'h24428800;
      22070: inst = 32'h8620000;
      22071: inst = 32'h2a0e0008;
      22072: inst = 32'h294f0001;
      22073: inst = 32'h11200000;
      22074: inst = 32'hd20563e;
      22075: inst = 32'h13e00000;
      22076: inst = 32'hfe0aa19;
      22077: inst = 32'h5be00000;
      22078: inst = 32'h244c8000;
      22079: inst = 32'h24428800;
      22080: inst = 32'h8620000;
      22081: inst = 32'h2a0e0009;
      22082: inst = 32'h294f0001;
      22083: inst = 32'h11200000;
      22084: inst = 32'hd205648;
      22085: inst = 32'h13e00000;
      22086: inst = 32'hfe0aa19;
      22087: inst = 32'h5be00000;
      22088: inst = 32'h244c8000;
      22089: inst = 32'h24428800;
      22090: inst = 32'h8620000;
      22091: inst = 32'h2a0e0000;
      22092: inst = 32'h294f0002;
      22093: inst = 32'h11200000;
      22094: inst = 32'hd205652;
      22095: inst = 32'h13e00000;
      22096: inst = 32'hfe0aa19;
      22097: inst = 32'h5be00000;
      22098: inst = 32'h244c8000;
      22099: inst = 32'h24428800;
      22100: inst = 32'h8620000;
      22101: inst = 32'h2a0e0001;
      22102: inst = 32'h294f0002;
      22103: inst = 32'h11200000;
      22104: inst = 32'hd20565c;
      22105: inst = 32'h13e00000;
      22106: inst = 32'hfe0aa19;
      22107: inst = 32'h5be00000;
      22108: inst = 32'h244c8000;
      22109: inst = 32'h24428800;
      22110: inst = 32'h8620000;
      22111: inst = 32'h2a0e0002;
      22112: inst = 32'h294f0002;
      22113: inst = 32'h11200000;
      22114: inst = 32'hd205666;
      22115: inst = 32'h13e00000;
      22116: inst = 32'hfe0aa19;
      22117: inst = 32'h5be00000;
      22118: inst = 32'h244c8000;
      22119: inst = 32'h24428800;
      22120: inst = 32'h8620000;
      22121: inst = 32'h2a0e0003;
      22122: inst = 32'h294f0002;
      22123: inst = 32'h11200000;
      22124: inst = 32'hd205670;
      22125: inst = 32'h13e00000;
      22126: inst = 32'hfe0aa19;
      22127: inst = 32'h5be00000;
      22128: inst = 32'h244c8000;
      22129: inst = 32'h24428800;
      22130: inst = 32'h8620000;
      22131: inst = 32'h2a0e0004;
      22132: inst = 32'h294f0002;
      22133: inst = 32'h11200000;
      22134: inst = 32'hd20567a;
      22135: inst = 32'h13e00000;
      22136: inst = 32'hfe0aa19;
      22137: inst = 32'h5be00000;
      22138: inst = 32'h244c8000;
      22139: inst = 32'h24428800;
      22140: inst = 32'h8620000;
      22141: inst = 32'h2a0e0005;
      22142: inst = 32'h294f0002;
      22143: inst = 32'h11200000;
      22144: inst = 32'hd205684;
      22145: inst = 32'h13e00000;
      22146: inst = 32'hfe0aa19;
      22147: inst = 32'h5be00000;
      22148: inst = 32'h244c8000;
      22149: inst = 32'h24428800;
      22150: inst = 32'h8620000;
      22151: inst = 32'h2a0e0006;
      22152: inst = 32'h294f0002;
      22153: inst = 32'h11200000;
      22154: inst = 32'hd20568e;
      22155: inst = 32'h13e00000;
      22156: inst = 32'hfe0aa19;
      22157: inst = 32'h5be00000;
      22158: inst = 32'h244c8000;
      22159: inst = 32'h24428800;
      22160: inst = 32'h8620000;
      22161: inst = 32'h2a0e0007;
      22162: inst = 32'h294f0002;
      22163: inst = 32'h11200000;
      22164: inst = 32'hd205698;
      22165: inst = 32'h13e00000;
      22166: inst = 32'hfe0aa19;
      22167: inst = 32'h5be00000;
      22168: inst = 32'h244c8000;
      22169: inst = 32'h24428800;
      22170: inst = 32'h8620000;
      22171: inst = 32'h2a0e0008;
      22172: inst = 32'h294f0002;
      22173: inst = 32'h11200000;
      22174: inst = 32'hd2056a2;
      22175: inst = 32'h13e00000;
      22176: inst = 32'hfe0aa19;
      22177: inst = 32'h5be00000;
      22178: inst = 32'h244c8000;
      22179: inst = 32'h24428800;
      22180: inst = 32'h8620000;
      22181: inst = 32'h2a0e0009;
      22182: inst = 32'h294f0002;
      22183: inst = 32'h11200000;
      22184: inst = 32'hd2056ac;
      22185: inst = 32'h13e00000;
      22186: inst = 32'hfe0aa19;
      22187: inst = 32'h5be00000;
      22188: inst = 32'h244c8000;
      22189: inst = 32'h24428800;
      22190: inst = 32'h8620000;
      22191: inst = 32'h2a0e0000;
      22192: inst = 32'h294f0003;
      22193: inst = 32'h11200000;
      22194: inst = 32'hd2056b6;
      22195: inst = 32'h13e00000;
      22196: inst = 32'hfe0aa19;
      22197: inst = 32'h5be00000;
      22198: inst = 32'h244c8000;
      22199: inst = 32'h24428800;
      22200: inst = 32'h8620000;
      22201: inst = 32'h2a0e0001;
      22202: inst = 32'h294f0003;
      22203: inst = 32'h11200000;
      22204: inst = 32'hd2056c0;
      22205: inst = 32'h13e00000;
      22206: inst = 32'hfe0aa19;
      22207: inst = 32'h5be00000;
      22208: inst = 32'h244c8000;
      22209: inst = 32'h24428800;
      22210: inst = 32'h8620000;
      22211: inst = 32'h2a0e0002;
      22212: inst = 32'h294f0003;
      22213: inst = 32'h11200000;
      22214: inst = 32'hd2056ca;
      22215: inst = 32'h13e00000;
      22216: inst = 32'hfe0aa19;
      22217: inst = 32'h5be00000;
      22218: inst = 32'h244c8000;
      22219: inst = 32'h24428800;
      22220: inst = 32'h8620000;
      22221: inst = 32'h2a0e0003;
      22222: inst = 32'h294f0003;
      22223: inst = 32'h11200000;
      22224: inst = 32'hd2056d4;
      22225: inst = 32'h13e00000;
      22226: inst = 32'hfe0aa19;
      22227: inst = 32'h5be00000;
      22228: inst = 32'h244c8000;
      22229: inst = 32'h24428800;
      22230: inst = 32'h8620000;
      22231: inst = 32'h2a0e0004;
      22232: inst = 32'h294f0003;
      22233: inst = 32'h11200000;
      22234: inst = 32'hd2056de;
      22235: inst = 32'h13e00000;
      22236: inst = 32'hfe0aa19;
      22237: inst = 32'h5be00000;
      22238: inst = 32'h244c8000;
      22239: inst = 32'h24428800;
      22240: inst = 32'h8620000;
      22241: inst = 32'h2a0e0005;
      22242: inst = 32'h294f0003;
      22243: inst = 32'h11200000;
      22244: inst = 32'hd2056e8;
      22245: inst = 32'h13e00000;
      22246: inst = 32'hfe0aa19;
      22247: inst = 32'h5be00000;
      22248: inst = 32'h244c8000;
      22249: inst = 32'h24428800;
      22250: inst = 32'h8620000;
      22251: inst = 32'h2a0e0006;
      22252: inst = 32'h294f0003;
      22253: inst = 32'h11200000;
      22254: inst = 32'hd2056f2;
      22255: inst = 32'h13e00000;
      22256: inst = 32'hfe0aa19;
      22257: inst = 32'h5be00000;
      22258: inst = 32'h244c8000;
      22259: inst = 32'h24428800;
      22260: inst = 32'h8620000;
      22261: inst = 32'h2a0e0007;
      22262: inst = 32'h294f0003;
      22263: inst = 32'h11200000;
      22264: inst = 32'hd2056fc;
      22265: inst = 32'h13e00000;
      22266: inst = 32'hfe0aa19;
      22267: inst = 32'h5be00000;
      22268: inst = 32'h244c8000;
      22269: inst = 32'h24428800;
      22270: inst = 32'h8620000;
      22271: inst = 32'h2a0e0008;
      22272: inst = 32'h294f0003;
      22273: inst = 32'h11200000;
      22274: inst = 32'hd205706;
      22275: inst = 32'h13e00000;
      22276: inst = 32'hfe0aa19;
      22277: inst = 32'h5be00000;
      22278: inst = 32'h244c8000;
      22279: inst = 32'h24428800;
      22280: inst = 32'h8620000;
      22281: inst = 32'h2a0e0009;
      22282: inst = 32'h294f0003;
      22283: inst = 32'h11200000;
      22284: inst = 32'hd205710;
      22285: inst = 32'h13e00000;
      22286: inst = 32'hfe0aa19;
      22287: inst = 32'h5be00000;
      22288: inst = 32'h244c8000;
      22289: inst = 32'h24428800;
      22290: inst = 32'h8620000;
      22291: inst = 32'h2a0e0000;
      22292: inst = 32'h294f0004;
      22293: inst = 32'h11200000;
      22294: inst = 32'hd20571a;
      22295: inst = 32'h13e00000;
      22296: inst = 32'hfe0aa19;
      22297: inst = 32'h5be00000;
      22298: inst = 32'h244c8000;
      22299: inst = 32'h24428800;
      22300: inst = 32'h8620000;
      22301: inst = 32'h2a0e0001;
      22302: inst = 32'h294f0004;
      22303: inst = 32'h11200000;
      22304: inst = 32'hd205724;
      22305: inst = 32'h13e00000;
      22306: inst = 32'hfe0aa19;
      22307: inst = 32'h5be00000;
      22308: inst = 32'h244c8000;
      22309: inst = 32'h24428800;
      22310: inst = 32'h8620000;
      22311: inst = 32'h2a0e0002;
      22312: inst = 32'h294f0004;
      22313: inst = 32'h11200000;
      22314: inst = 32'hd20572e;
      22315: inst = 32'h13e00000;
      22316: inst = 32'hfe0aa19;
      22317: inst = 32'h5be00000;
      22318: inst = 32'h244c8000;
      22319: inst = 32'h24428800;
      22320: inst = 32'h8620000;
      22321: inst = 32'h2a0e0003;
      22322: inst = 32'h294f0004;
      22323: inst = 32'h11200000;
      22324: inst = 32'hd205738;
      22325: inst = 32'h13e00000;
      22326: inst = 32'hfe0aa19;
      22327: inst = 32'h5be00000;
      22328: inst = 32'h244c8000;
      22329: inst = 32'h24428800;
      22330: inst = 32'h8620000;
      22331: inst = 32'h2a0e0004;
      22332: inst = 32'h294f0004;
      22333: inst = 32'h11200000;
      22334: inst = 32'hd205742;
      22335: inst = 32'h13e00000;
      22336: inst = 32'hfe0aa19;
      22337: inst = 32'h5be00000;
      22338: inst = 32'h244c8000;
      22339: inst = 32'h24428800;
      22340: inst = 32'h8620000;
      22341: inst = 32'h2a0e0005;
      22342: inst = 32'h294f0004;
      22343: inst = 32'h11200000;
      22344: inst = 32'hd20574c;
      22345: inst = 32'h13e00000;
      22346: inst = 32'hfe0aa19;
      22347: inst = 32'h5be00000;
      22348: inst = 32'h244c8000;
      22349: inst = 32'h24428800;
      22350: inst = 32'h8620000;
      22351: inst = 32'h2a0e0006;
      22352: inst = 32'h294f0004;
      22353: inst = 32'h11200000;
      22354: inst = 32'hd205756;
      22355: inst = 32'h13e00000;
      22356: inst = 32'hfe0aa19;
      22357: inst = 32'h5be00000;
      22358: inst = 32'h244c8000;
      22359: inst = 32'h24428800;
      22360: inst = 32'h8620000;
      22361: inst = 32'h2a0e0007;
      22362: inst = 32'h294f0004;
      22363: inst = 32'h11200000;
      22364: inst = 32'hd205760;
      22365: inst = 32'h13e00000;
      22366: inst = 32'hfe0aa19;
      22367: inst = 32'h5be00000;
      22368: inst = 32'h244c8000;
      22369: inst = 32'h24428800;
      22370: inst = 32'h8620000;
      22371: inst = 32'h2a0e0008;
      22372: inst = 32'h294f0004;
      22373: inst = 32'h11200000;
      22374: inst = 32'hd20576a;
      22375: inst = 32'h13e00000;
      22376: inst = 32'hfe0aa19;
      22377: inst = 32'h5be00000;
      22378: inst = 32'h244c8000;
      22379: inst = 32'h24428800;
      22380: inst = 32'h8620000;
      22381: inst = 32'h2a0e0009;
      22382: inst = 32'h294f0004;
      22383: inst = 32'h11200000;
      22384: inst = 32'hd205774;
      22385: inst = 32'h13e00000;
      22386: inst = 32'hfe0aa19;
      22387: inst = 32'h5be00000;
      22388: inst = 32'h244c8000;
      22389: inst = 32'h24428800;
      22390: inst = 32'h8620000;
      22391: inst = 32'h2a0e0000;
      22392: inst = 32'h294f0005;
      22393: inst = 32'h11200000;
      22394: inst = 32'hd20577e;
      22395: inst = 32'h13e00000;
      22396: inst = 32'hfe0aa19;
      22397: inst = 32'h5be00000;
      22398: inst = 32'h244c8000;
      22399: inst = 32'h24428800;
      22400: inst = 32'h8620000;
      22401: inst = 32'h2a0e0001;
      22402: inst = 32'h294f0005;
      22403: inst = 32'h11200000;
      22404: inst = 32'hd205788;
      22405: inst = 32'h13e00000;
      22406: inst = 32'hfe0aa19;
      22407: inst = 32'h5be00000;
      22408: inst = 32'h244c8000;
      22409: inst = 32'h24428800;
      22410: inst = 32'h8620000;
      22411: inst = 32'h2a0e0002;
      22412: inst = 32'h294f0005;
      22413: inst = 32'h11200000;
      22414: inst = 32'hd205792;
      22415: inst = 32'h13e00000;
      22416: inst = 32'hfe0aa19;
      22417: inst = 32'h5be00000;
      22418: inst = 32'h244c8000;
      22419: inst = 32'h24428800;
      22420: inst = 32'h8620000;
      22421: inst = 32'h2a0e0003;
      22422: inst = 32'h294f0005;
      22423: inst = 32'h11200000;
      22424: inst = 32'hd20579c;
      22425: inst = 32'h13e00000;
      22426: inst = 32'hfe0aa19;
      22427: inst = 32'h5be00000;
      22428: inst = 32'h244c8000;
      22429: inst = 32'h24428800;
      22430: inst = 32'h8620000;
      22431: inst = 32'h2a0e0004;
      22432: inst = 32'h294f0005;
      22433: inst = 32'h11200000;
      22434: inst = 32'hd2057a6;
      22435: inst = 32'h13e00000;
      22436: inst = 32'hfe0aa19;
      22437: inst = 32'h5be00000;
      22438: inst = 32'h244c8000;
      22439: inst = 32'h24428800;
      22440: inst = 32'h8620000;
      22441: inst = 32'h2a0e0005;
      22442: inst = 32'h294f0005;
      22443: inst = 32'h11200000;
      22444: inst = 32'hd2057b0;
      22445: inst = 32'h13e00000;
      22446: inst = 32'hfe0aa19;
      22447: inst = 32'h5be00000;
      22448: inst = 32'h244c8000;
      22449: inst = 32'h24428800;
      22450: inst = 32'h8620000;
      22451: inst = 32'h2a0e0006;
      22452: inst = 32'h294f0005;
      22453: inst = 32'h11200000;
      22454: inst = 32'hd2057ba;
      22455: inst = 32'h13e00000;
      22456: inst = 32'hfe0aa19;
      22457: inst = 32'h5be00000;
      22458: inst = 32'h244c8000;
      22459: inst = 32'h24428800;
      22460: inst = 32'h8620000;
      22461: inst = 32'h2a0e0007;
      22462: inst = 32'h294f0005;
      22463: inst = 32'h11200000;
      22464: inst = 32'hd2057c4;
      22465: inst = 32'h13e00000;
      22466: inst = 32'hfe0aa19;
      22467: inst = 32'h5be00000;
      22468: inst = 32'h244c8000;
      22469: inst = 32'h24428800;
      22470: inst = 32'h8620000;
      22471: inst = 32'h2a0e0008;
      22472: inst = 32'h294f0005;
      22473: inst = 32'h11200000;
      22474: inst = 32'hd2057ce;
      22475: inst = 32'h13e00000;
      22476: inst = 32'hfe0aa19;
      22477: inst = 32'h5be00000;
      22478: inst = 32'h244c8000;
      22479: inst = 32'h24428800;
      22480: inst = 32'h8620000;
      22481: inst = 32'h2a0e0009;
      22482: inst = 32'h294f0005;
      22483: inst = 32'h11200000;
      22484: inst = 32'hd2057d8;
      22485: inst = 32'h13e00000;
      22486: inst = 32'hfe0aa19;
      22487: inst = 32'h5be00000;
      22488: inst = 32'h244c8000;
      22489: inst = 32'h24428800;
      22490: inst = 32'h8620000;
      22491: inst = 32'h2a0e0000;
      22492: inst = 32'h294f0006;
      22493: inst = 32'h11200000;
      22494: inst = 32'hd2057e2;
      22495: inst = 32'h13e00000;
      22496: inst = 32'hfe0aa19;
      22497: inst = 32'h5be00000;
      22498: inst = 32'h244c8000;
      22499: inst = 32'h24428800;
      22500: inst = 32'h8620000;
      22501: inst = 32'h2a0e0001;
      22502: inst = 32'h294f0006;
      22503: inst = 32'h11200000;
      22504: inst = 32'hd2057ec;
      22505: inst = 32'h13e00000;
      22506: inst = 32'hfe0aa19;
      22507: inst = 32'h5be00000;
      22508: inst = 32'h244c8000;
      22509: inst = 32'h24428800;
      22510: inst = 32'h8620000;
      22511: inst = 32'h2a0e0002;
      22512: inst = 32'h294f0006;
      22513: inst = 32'h11200000;
      22514: inst = 32'hd2057f6;
      22515: inst = 32'h13e00000;
      22516: inst = 32'hfe0aa19;
      22517: inst = 32'h5be00000;
      22518: inst = 32'h244c8000;
      22519: inst = 32'h24428800;
      22520: inst = 32'h8620000;
      22521: inst = 32'h2a0e0003;
      22522: inst = 32'h294f0006;
      22523: inst = 32'h11200000;
      22524: inst = 32'hd205800;
      22525: inst = 32'h13e00000;
      22526: inst = 32'hfe0aa19;
      22527: inst = 32'h5be00000;
      22528: inst = 32'h244c8000;
      22529: inst = 32'h24428800;
      22530: inst = 32'h8620000;
      22531: inst = 32'h2a0e0004;
      22532: inst = 32'h294f0006;
      22533: inst = 32'h11200000;
      22534: inst = 32'hd20580a;
      22535: inst = 32'h13e00000;
      22536: inst = 32'hfe0aa19;
      22537: inst = 32'h5be00000;
      22538: inst = 32'h244c8000;
      22539: inst = 32'h24428800;
      22540: inst = 32'h8620000;
      22541: inst = 32'h2a0e0005;
      22542: inst = 32'h294f0006;
      22543: inst = 32'h11200000;
      22544: inst = 32'hd205814;
      22545: inst = 32'h13e00000;
      22546: inst = 32'hfe0aa19;
      22547: inst = 32'h5be00000;
      22548: inst = 32'h244c8000;
      22549: inst = 32'h24428800;
      22550: inst = 32'h8620000;
      22551: inst = 32'h2a0e0006;
      22552: inst = 32'h294f0006;
      22553: inst = 32'h11200000;
      22554: inst = 32'hd20581e;
      22555: inst = 32'h13e00000;
      22556: inst = 32'hfe0aa19;
      22557: inst = 32'h5be00000;
      22558: inst = 32'h244c8000;
      22559: inst = 32'h24428800;
      22560: inst = 32'h8620000;
      22561: inst = 32'h2a0e0007;
      22562: inst = 32'h294f0006;
      22563: inst = 32'h11200000;
      22564: inst = 32'hd205828;
      22565: inst = 32'h13e00000;
      22566: inst = 32'hfe0aa19;
      22567: inst = 32'h5be00000;
      22568: inst = 32'h244c8000;
      22569: inst = 32'h24428800;
      22570: inst = 32'h8620000;
      22571: inst = 32'h2a0e0008;
      22572: inst = 32'h294f0006;
      22573: inst = 32'h11200000;
      22574: inst = 32'hd205832;
      22575: inst = 32'h13e00000;
      22576: inst = 32'hfe0aa19;
      22577: inst = 32'h5be00000;
      22578: inst = 32'h244c8000;
      22579: inst = 32'h24428800;
      22580: inst = 32'h8620000;
      22581: inst = 32'h2a0e0009;
      22582: inst = 32'h294f0006;
      22583: inst = 32'h11200000;
      22584: inst = 32'hd20583c;
      22585: inst = 32'h13e00000;
      22586: inst = 32'hfe0aa19;
      22587: inst = 32'h5be00000;
      22588: inst = 32'h244c8000;
      22589: inst = 32'h24428800;
      22590: inst = 32'h8620000;
      22591: inst = 32'hc60f4ce;
      22592: inst = 32'h2a0e0001;
      22593: inst = 32'h294f0007;
      22594: inst = 32'h11200000;
      22595: inst = 32'hd205847;
      22596: inst = 32'h13e00000;
      22597: inst = 32'hfe0aa19;
      22598: inst = 32'h5be00000;
      22599: inst = 32'h244c8000;
      22600: inst = 32'h24428800;
      22601: inst = 32'h8620000;
      22602: inst = 32'h2a0e0008;
      22603: inst = 32'h294f0007;
      22604: inst = 32'h11200000;
      22605: inst = 32'hd205851;
      22606: inst = 32'h13e00000;
      22607: inst = 32'hfe0aa19;
      22608: inst = 32'h5be00000;
      22609: inst = 32'h244c8000;
      22610: inst = 32'h24428800;
      22611: inst = 32'h8620000;
      22612: inst = 32'h2a0e0001;
      22613: inst = 32'h294f0008;
      22614: inst = 32'h11200000;
      22615: inst = 32'hd20585b;
      22616: inst = 32'h13e00000;
      22617: inst = 32'hfe0aa19;
      22618: inst = 32'h5be00000;
      22619: inst = 32'h244c8000;
      22620: inst = 32'h24428800;
      22621: inst = 32'h8620000;
      22622: inst = 32'h2a0e0008;
      22623: inst = 32'h294f0008;
      22624: inst = 32'h11200000;
      22625: inst = 32'hd205865;
      22626: inst = 32'h13e00000;
      22627: inst = 32'hfe0aa19;
      22628: inst = 32'h5be00000;
      22629: inst = 32'h244c8000;
      22630: inst = 32'h24428800;
      22631: inst = 32'h8620000;
      22632: inst = 32'hc607841;
      22633: inst = 32'h2a0e0002;
      22634: inst = 32'h294f0007;
      22635: inst = 32'h11200000;
      22636: inst = 32'hd205870;
      22637: inst = 32'h13e00000;
      22638: inst = 32'hfe0aa19;
      22639: inst = 32'h5be00000;
      22640: inst = 32'h244c8000;
      22641: inst = 32'h24428800;
      22642: inst = 32'h8620000;
      22643: inst = 32'h2a0e0003;
      22644: inst = 32'h294f0007;
      22645: inst = 32'h11200000;
      22646: inst = 32'hd20587a;
      22647: inst = 32'h13e00000;
      22648: inst = 32'hfe0aa19;
      22649: inst = 32'h5be00000;
      22650: inst = 32'h244c8000;
      22651: inst = 32'h24428800;
      22652: inst = 32'h8620000;
      22653: inst = 32'h2a0e0004;
      22654: inst = 32'h294f0007;
      22655: inst = 32'h11200000;
      22656: inst = 32'hd205884;
      22657: inst = 32'h13e00000;
      22658: inst = 32'hfe0aa19;
      22659: inst = 32'h5be00000;
      22660: inst = 32'h244c8000;
      22661: inst = 32'h24428800;
      22662: inst = 32'h8620000;
      22663: inst = 32'h2a0e0005;
      22664: inst = 32'h294f0007;
      22665: inst = 32'h11200000;
      22666: inst = 32'hd20588e;
      22667: inst = 32'h13e00000;
      22668: inst = 32'hfe0aa19;
      22669: inst = 32'h5be00000;
      22670: inst = 32'h244c8000;
      22671: inst = 32'h24428800;
      22672: inst = 32'h8620000;
      22673: inst = 32'h2a0e0006;
      22674: inst = 32'h294f0007;
      22675: inst = 32'h11200000;
      22676: inst = 32'hd205898;
      22677: inst = 32'h13e00000;
      22678: inst = 32'hfe0aa19;
      22679: inst = 32'h5be00000;
      22680: inst = 32'h244c8000;
      22681: inst = 32'h24428800;
      22682: inst = 32'h8620000;
      22683: inst = 32'h2a0e0007;
      22684: inst = 32'h294f0007;
      22685: inst = 32'h11200000;
      22686: inst = 32'hd2058a2;
      22687: inst = 32'h13e00000;
      22688: inst = 32'hfe0aa19;
      22689: inst = 32'h5be00000;
      22690: inst = 32'h244c8000;
      22691: inst = 32'h24428800;
      22692: inst = 32'h8620000;
      22693: inst = 32'h2a0e0002;
      22694: inst = 32'h294f0008;
      22695: inst = 32'h11200000;
      22696: inst = 32'hd2058ac;
      22697: inst = 32'h13e00000;
      22698: inst = 32'hfe0aa19;
      22699: inst = 32'h5be00000;
      22700: inst = 32'h244c8000;
      22701: inst = 32'h24428800;
      22702: inst = 32'h8620000;
      22703: inst = 32'h2a0e0003;
      22704: inst = 32'h294f0008;
      22705: inst = 32'h11200000;
      22706: inst = 32'hd2058b6;
      22707: inst = 32'h13e00000;
      22708: inst = 32'hfe0aa19;
      22709: inst = 32'h5be00000;
      22710: inst = 32'h244c8000;
      22711: inst = 32'h24428800;
      22712: inst = 32'h8620000;
      22713: inst = 32'h2a0e0004;
      22714: inst = 32'h294f0008;
      22715: inst = 32'h11200000;
      22716: inst = 32'hd2058c0;
      22717: inst = 32'h13e00000;
      22718: inst = 32'hfe0aa19;
      22719: inst = 32'h5be00000;
      22720: inst = 32'h244c8000;
      22721: inst = 32'h24428800;
      22722: inst = 32'h8620000;
      22723: inst = 32'h2a0e0005;
      22724: inst = 32'h294f0008;
      22725: inst = 32'h11200000;
      22726: inst = 32'hd2058ca;
      22727: inst = 32'h13e00000;
      22728: inst = 32'hfe0aa19;
      22729: inst = 32'h5be00000;
      22730: inst = 32'h244c8000;
      22731: inst = 32'h24428800;
      22732: inst = 32'h8620000;
      22733: inst = 32'h2a0e0006;
      22734: inst = 32'h294f0008;
      22735: inst = 32'h11200000;
      22736: inst = 32'hd2058d4;
      22737: inst = 32'h13e00000;
      22738: inst = 32'hfe0aa19;
      22739: inst = 32'h5be00000;
      22740: inst = 32'h244c8000;
      22741: inst = 32'h24428800;
      22742: inst = 32'h8620000;
      22743: inst = 32'h2a0e0007;
      22744: inst = 32'h294f0008;
      22745: inst = 32'h11200000;
      22746: inst = 32'hd2058de;
      22747: inst = 32'h13e00000;
      22748: inst = 32'hfe0aa19;
      22749: inst = 32'h5be00000;
      22750: inst = 32'h244c8000;
      22751: inst = 32'h24428800;
      22752: inst = 32'h8620000;
      22753: inst = 32'h2a0e0002;
      22754: inst = 32'h294f0009;
      22755: inst = 32'h11200000;
      22756: inst = 32'hd2058e8;
      22757: inst = 32'h13e00000;
      22758: inst = 32'hfe0aa19;
      22759: inst = 32'h5be00000;
      22760: inst = 32'h244c8000;
      22761: inst = 32'h24428800;
      22762: inst = 32'h8620000;
      22763: inst = 32'h2a0e0003;
      22764: inst = 32'h294f0009;
      22765: inst = 32'h11200000;
      22766: inst = 32'hd2058f2;
      22767: inst = 32'h13e00000;
      22768: inst = 32'hfe0aa19;
      22769: inst = 32'h5be00000;
      22770: inst = 32'h244c8000;
      22771: inst = 32'h24428800;
      22772: inst = 32'h8620000;
      22773: inst = 32'h2a0e0004;
      22774: inst = 32'h294f0009;
      22775: inst = 32'h11200000;
      22776: inst = 32'hd2058fc;
      22777: inst = 32'h13e00000;
      22778: inst = 32'hfe0aa19;
      22779: inst = 32'h5be00000;
      22780: inst = 32'h244c8000;
      22781: inst = 32'h24428800;
      22782: inst = 32'h8620000;
      22783: inst = 32'h2a0e0005;
      22784: inst = 32'h294f0009;
      22785: inst = 32'h11200000;
      22786: inst = 32'hd205906;
      22787: inst = 32'h13e00000;
      22788: inst = 32'hfe0aa19;
      22789: inst = 32'h5be00000;
      22790: inst = 32'h244c8000;
      22791: inst = 32'h24428800;
      22792: inst = 32'h8620000;
      22793: inst = 32'h2a0e0006;
      22794: inst = 32'h294f0009;
      22795: inst = 32'h11200000;
      22796: inst = 32'hd205910;
      22797: inst = 32'h13e00000;
      22798: inst = 32'hfe0aa19;
      22799: inst = 32'h5be00000;
      22800: inst = 32'h244c8000;
      22801: inst = 32'h24428800;
      22802: inst = 32'h8620000;
      22803: inst = 32'h2a0e0007;
      22804: inst = 32'h294f0009;
      22805: inst = 32'h11200000;
      22806: inst = 32'hd20591a;
      22807: inst = 32'h13e00000;
      22808: inst = 32'hfe0aa19;
      22809: inst = 32'h5be00000;
      22810: inst = 32'h244c8000;
      22811: inst = 32'h24428800;
      22812: inst = 32'h8620000;
      22813: inst = 32'hc6010ac;
      22814: inst = 32'h2a0e0002;
      22815: inst = 32'h294f000a;
      22816: inst = 32'h11200000;
      22817: inst = 32'hd205925;
      22818: inst = 32'h13e00000;
      22819: inst = 32'hfe0aa19;
      22820: inst = 32'h5be00000;
      22821: inst = 32'h244c8000;
      22822: inst = 32'h24428800;
      22823: inst = 32'h8620000;
      22824: inst = 32'h2a0e0003;
      22825: inst = 32'h294f000a;
      22826: inst = 32'h11200000;
      22827: inst = 32'hd20592f;
      22828: inst = 32'h13e00000;
      22829: inst = 32'hfe0aa19;
      22830: inst = 32'h5be00000;
      22831: inst = 32'h244c8000;
      22832: inst = 32'h24428800;
      22833: inst = 32'h8620000;
      22834: inst = 32'h2a0e0004;
      22835: inst = 32'h294f000a;
      22836: inst = 32'h11200000;
      22837: inst = 32'hd205939;
      22838: inst = 32'h13e00000;
      22839: inst = 32'hfe0aa19;
      22840: inst = 32'h5be00000;
      22841: inst = 32'h244c8000;
      22842: inst = 32'h24428800;
      22843: inst = 32'h8620000;
      22844: inst = 32'h2a0e0005;
      22845: inst = 32'h294f000a;
      22846: inst = 32'h11200000;
      22847: inst = 32'hd205943;
      22848: inst = 32'h13e00000;
      22849: inst = 32'hfe0aa19;
      22850: inst = 32'h5be00000;
      22851: inst = 32'h244c8000;
      22852: inst = 32'h24428800;
      22853: inst = 32'h8620000;
      22854: inst = 32'h2a0e0006;
      22855: inst = 32'h294f000a;
      22856: inst = 32'h11200000;
      22857: inst = 32'hd20594d;
      22858: inst = 32'h13e00000;
      22859: inst = 32'hfe0aa19;
      22860: inst = 32'h5be00000;
      22861: inst = 32'h244c8000;
      22862: inst = 32'h24428800;
      22863: inst = 32'h8620000;
      22864: inst = 32'h2a0e0007;
      22865: inst = 32'h294f000a;
      22866: inst = 32'h11200000;
      22867: inst = 32'hd205957;
      22868: inst = 32'h13e00000;
      22869: inst = 32'hfe0aa19;
      22870: inst = 32'h5be00000;
      22871: inst = 32'h244c8000;
      22872: inst = 32'h24428800;
      22873: inst = 32'h8620000;
      22874: inst = 32'hc60d42c;
      22875: inst = 32'h2a0e0003;
      22876: inst = 32'h294f000b;
      22877: inst = 32'h11200000;
      22878: inst = 32'hd205962;
      22879: inst = 32'h13e00000;
      22880: inst = 32'hfe0aa19;
      22881: inst = 32'h5be00000;
      22882: inst = 32'h244c8000;
      22883: inst = 32'h24428800;
      22884: inst = 32'h8620000;
      22885: inst = 32'h2a0e0006;
      22886: inst = 32'h294f000b;
      22887: inst = 32'h11200000;
      22888: inst = 32'hd20596c;
      22889: inst = 32'h13e00000;
      22890: inst = 32'hfe0aa19;
      22891: inst = 32'h5be00000;
      22892: inst = 32'h244c8000;
      22893: inst = 32'h24428800;
      22894: inst = 32'h8620000;
      22895: inst = 32'h13e00000;
      22896: inst = 32'hfe06126;
      22897: inst = 32'h5be00000;
      22898: inst = 32'hc6018c3;
      22899: inst = 32'h2a0e0000;
      22900: inst = 32'h294f0000;
      22901: inst = 32'h11200000;
      22902: inst = 32'hd20597a;
      22903: inst = 32'h13e00000;
      22904: inst = 32'hfe0aa19;
      22905: inst = 32'h5be00000;
      22906: inst = 32'h244c8000;
      22907: inst = 32'h24428800;
      22908: inst = 32'h8620000;
      22909: inst = 32'h2a0e0001;
      22910: inst = 32'h294f0000;
      22911: inst = 32'h11200000;
      22912: inst = 32'hd205984;
      22913: inst = 32'h13e00000;
      22914: inst = 32'hfe0aa19;
      22915: inst = 32'h5be00000;
      22916: inst = 32'h244c8000;
      22917: inst = 32'h24428800;
      22918: inst = 32'h8620000;
      22919: inst = 32'h2a0e0002;
      22920: inst = 32'h294f0000;
      22921: inst = 32'h11200000;
      22922: inst = 32'hd20598e;
      22923: inst = 32'h13e00000;
      22924: inst = 32'hfe0aa19;
      22925: inst = 32'h5be00000;
      22926: inst = 32'h244c8000;
      22927: inst = 32'h24428800;
      22928: inst = 32'h8620000;
      22929: inst = 32'h2a0e0003;
      22930: inst = 32'h294f0000;
      22931: inst = 32'h11200000;
      22932: inst = 32'hd205998;
      22933: inst = 32'h13e00000;
      22934: inst = 32'hfe0aa19;
      22935: inst = 32'h5be00000;
      22936: inst = 32'h244c8000;
      22937: inst = 32'h24428800;
      22938: inst = 32'h8620000;
      22939: inst = 32'h2a0e0004;
      22940: inst = 32'h294f0000;
      22941: inst = 32'h11200000;
      22942: inst = 32'hd2059a2;
      22943: inst = 32'h13e00000;
      22944: inst = 32'hfe0aa19;
      22945: inst = 32'h5be00000;
      22946: inst = 32'h244c8000;
      22947: inst = 32'h24428800;
      22948: inst = 32'h8620000;
      22949: inst = 32'h2a0e0005;
      22950: inst = 32'h294f0000;
      22951: inst = 32'h11200000;
      22952: inst = 32'hd2059ac;
      22953: inst = 32'h13e00000;
      22954: inst = 32'hfe0aa19;
      22955: inst = 32'h5be00000;
      22956: inst = 32'h244c8000;
      22957: inst = 32'h24428800;
      22958: inst = 32'h8620000;
      22959: inst = 32'h2a0e0006;
      22960: inst = 32'h294f0000;
      22961: inst = 32'h11200000;
      22962: inst = 32'hd2059b6;
      22963: inst = 32'h13e00000;
      22964: inst = 32'hfe0aa19;
      22965: inst = 32'h5be00000;
      22966: inst = 32'h244c8000;
      22967: inst = 32'h24428800;
      22968: inst = 32'h8620000;
      22969: inst = 32'h2a0e0007;
      22970: inst = 32'h294f0000;
      22971: inst = 32'h11200000;
      22972: inst = 32'hd2059c0;
      22973: inst = 32'h13e00000;
      22974: inst = 32'hfe0aa19;
      22975: inst = 32'h5be00000;
      22976: inst = 32'h244c8000;
      22977: inst = 32'h24428800;
      22978: inst = 32'h8620000;
      22979: inst = 32'h2a0e0008;
      22980: inst = 32'h294f0000;
      22981: inst = 32'h11200000;
      22982: inst = 32'hd2059ca;
      22983: inst = 32'h13e00000;
      22984: inst = 32'hfe0aa19;
      22985: inst = 32'h5be00000;
      22986: inst = 32'h244c8000;
      22987: inst = 32'h24428800;
      22988: inst = 32'h8620000;
      22989: inst = 32'h2a0e0009;
      22990: inst = 32'h294f0000;
      22991: inst = 32'h11200000;
      22992: inst = 32'hd2059d4;
      22993: inst = 32'h13e00000;
      22994: inst = 32'hfe0aa19;
      22995: inst = 32'h5be00000;
      22996: inst = 32'h244c8000;
      22997: inst = 32'h24428800;
      22998: inst = 32'h8620000;
      22999: inst = 32'h2a0e0000;
      23000: inst = 32'h294f0001;
      23001: inst = 32'h11200000;
      23002: inst = 32'hd2059de;
      23003: inst = 32'h13e00000;
      23004: inst = 32'hfe0aa19;
      23005: inst = 32'h5be00000;
      23006: inst = 32'h244c8000;
      23007: inst = 32'h24428800;
      23008: inst = 32'h8620000;
      23009: inst = 32'h2a0e0001;
      23010: inst = 32'h294f0001;
      23011: inst = 32'h11200000;
      23012: inst = 32'hd2059e8;
      23013: inst = 32'h13e00000;
      23014: inst = 32'hfe0aa19;
      23015: inst = 32'h5be00000;
      23016: inst = 32'h244c8000;
      23017: inst = 32'h24428800;
      23018: inst = 32'h8620000;
      23019: inst = 32'h2a0e0002;
      23020: inst = 32'h294f0001;
      23021: inst = 32'h11200000;
      23022: inst = 32'hd2059f2;
      23023: inst = 32'h13e00000;
      23024: inst = 32'hfe0aa19;
      23025: inst = 32'h5be00000;
      23026: inst = 32'h244c8000;
      23027: inst = 32'h24428800;
      23028: inst = 32'h8620000;
      23029: inst = 32'h2a0e0003;
      23030: inst = 32'h294f0001;
      23031: inst = 32'h11200000;
      23032: inst = 32'hd2059fc;
      23033: inst = 32'h13e00000;
      23034: inst = 32'hfe0aa19;
      23035: inst = 32'h5be00000;
      23036: inst = 32'h244c8000;
      23037: inst = 32'h24428800;
      23038: inst = 32'h8620000;
      23039: inst = 32'h2a0e0004;
      23040: inst = 32'h294f0001;
      23041: inst = 32'h11200000;
      23042: inst = 32'hd205a06;
      23043: inst = 32'h13e00000;
      23044: inst = 32'hfe0aa19;
      23045: inst = 32'h5be00000;
      23046: inst = 32'h244c8000;
      23047: inst = 32'h24428800;
      23048: inst = 32'h8620000;
      23049: inst = 32'h2a0e0005;
      23050: inst = 32'h294f0001;
      23051: inst = 32'h11200000;
      23052: inst = 32'hd205a10;
      23053: inst = 32'h13e00000;
      23054: inst = 32'hfe0aa19;
      23055: inst = 32'h5be00000;
      23056: inst = 32'h244c8000;
      23057: inst = 32'h24428800;
      23058: inst = 32'h8620000;
      23059: inst = 32'h2a0e0006;
      23060: inst = 32'h294f0001;
      23061: inst = 32'h11200000;
      23062: inst = 32'hd205a1a;
      23063: inst = 32'h13e00000;
      23064: inst = 32'hfe0aa19;
      23065: inst = 32'h5be00000;
      23066: inst = 32'h244c8000;
      23067: inst = 32'h24428800;
      23068: inst = 32'h8620000;
      23069: inst = 32'h2a0e0007;
      23070: inst = 32'h294f0001;
      23071: inst = 32'h11200000;
      23072: inst = 32'hd205a24;
      23073: inst = 32'h13e00000;
      23074: inst = 32'hfe0aa19;
      23075: inst = 32'h5be00000;
      23076: inst = 32'h244c8000;
      23077: inst = 32'h24428800;
      23078: inst = 32'h8620000;
      23079: inst = 32'h2a0e0008;
      23080: inst = 32'h294f0001;
      23081: inst = 32'h11200000;
      23082: inst = 32'hd205a2e;
      23083: inst = 32'h13e00000;
      23084: inst = 32'hfe0aa19;
      23085: inst = 32'h5be00000;
      23086: inst = 32'h244c8000;
      23087: inst = 32'h24428800;
      23088: inst = 32'h8620000;
      23089: inst = 32'h2a0e0009;
      23090: inst = 32'h294f0001;
      23091: inst = 32'h11200000;
      23092: inst = 32'hd205a38;
      23093: inst = 32'h13e00000;
      23094: inst = 32'hfe0aa19;
      23095: inst = 32'h5be00000;
      23096: inst = 32'h244c8000;
      23097: inst = 32'h24428800;
      23098: inst = 32'h8620000;
      23099: inst = 32'h2a0e0000;
      23100: inst = 32'h294f0002;
      23101: inst = 32'h11200000;
      23102: inst = 32'hd205a42;
      23103: inst = 32'h13e00000;
      23104: inst = 32'hfe0aa19;
      23105: inst = 32'h5be00000;
      23106: inst = 32'h244c8000;
      23107: inst = 32'h24428800;
      23108: inst = 32'h8620000;
      23109: inst = 32'h2a0e0001;
      23110: inst = 32'h294f0002;
      23111: inst = 32'h11200000;
      23112: inst = 32'hd205a4c;
      23113: inst = 32'h13e00000;
      23114: inst = 32'hfe0aa19;
      23115: inst = 32'h5be00000;
      23116: inst = 32'h244c8000;
      23117: inst = 32'h24428800;
      23118: inst = 32'h8620000;
      23119: inst = 32'h2a0e0000;
      23120: inst = 32'h294f0003;
      23121: inst = 32'h11200000;
      23122: inst = 32'hd205a56;
      23123: inst = 32'h13e00000;
      23124: inst = 32'hfe0aa19;
      23125: inst = 32'h5be00000;
      23126: inst = 32'h244c8000;
      23127: inst = 32'h24428800;
      23128: inst = 32'h8620000;
      23129: inst = 32'h2a0e0008;
      23130: inst = 32'h294f0003;
      23131: inst = 32'h11200000;
      23132: inst = 32'hd205a60;
      23133: inst = 32'h13e00000;
      23134: inst = 32'hfe0aa19;
      23135: inst = 32'h5be00000;
      23136: inst = 32'h244c8000;
      23137: inst = 32'h24428800;
      23138: inst = 32'h8620000;
      23139: inst = 32'h2a0e0000;
      23140: inst = 32'h294f0004;
      23141: inst = 32'h11200000;
      23142: inst = 32'hd205a6a;
      23143: inst = 32'h13e00000;
      23144: inst = 32'hfe0aa19;
      23145: inst = 32'h5be00000;
      23146: inst = 32'h244c8000;
      23147: inst = 32'h24428800;
      23148: inst = 32'h8620000;
      23149: inst = 32'h2a0e0008;
      23150: inst = 32'h294f0004;
      23151: inst = 32'h11200000;
      23152: inst = 32'hd205a74;
      23153: inst = 32'h13e00000;
      23154: inst = 32'hfe0aa19;
      23155: inst = 32'h5be00000;
      23156: inst = 32'h244c8000;
      23157: inst = 32'h24428800;
      23158: inst = 32'h8620000;
      23159: inst = 32'h2a0e0000;
      23160: inst = 32'h294f0005;
      23161: inst = 32'h11200000;
      23162: inst = 32'hd205a7e;
      23163: inst = 32'h13e00000;
      23164: inst = 32'hfe0aa19;
      23165: inst = 32'h5be00000;
      23166: inst = 32'h244c8000;
      23167: inst = 32'h24428800;
      23168: inst = 32'h8620000;
      23169: inst = 32'h2a0e0001;
      23170: inst = 32'h294f0005;
      23171: inst = 32'h11200000;
      23172: inst = 32'hd205a88;
      23173: inst = 32'h13e00000;
      23174: inst = 32'hfe0aa19;
      23175: inst = 32'h5be00000;
      23176: inst = 32'h244c8000;
      23177: inst = 32'h24428800;
      23178: inst = 32'h8620000;
      23179: inst = 32'h2a0e0000;
      23180: inst = 32'h294f0006;
      23181: inst = 32'h11200000;
      23182: inst = 32'hd205a92;
      23183: inst = 32'h13e00000;
      23184: inst = 32'hfe0aa19;
      23185: inst = 32'h5be00000;
      23186: inst = 32'h244c8000;
      23187: inst = 32'h24428800;
      23188: inst = 32'h8620000;
      23189: inst = 32'h2a0e0001;
      23190: inst = 32'h294f0006;
      23191: inst = 32'h11200000;
      23192: inst = 32'hd205a9c;
      23193: inst = 32'h13e00000;
      23194: inst = 32'hfe0aa19;
      23195: inst = 32'h5be00000;
      23196: inst = 32'h244c8000;
      23197: inst = 32'h24428800;
      23198: inst = 32'h8620000;
      23199: inst = 32'hc60d42c;
      23200: inst = 32'h2a0e0002;
      23201: inst = 32'h294f0002;
      23202: inst = 32'h11200000;
      23203: inst = 32'hd205aa7;
      23204: inst = 32'h13e00000;
      23205: inst = 32'hfe0aa19;
      23206: inst = 32'h5be00000;
      23207: inst = 32'h244c8000;
      23208: inst = 32'h24428800;
      23209: inst = 32'h8620000;
      23210: inst = 32'h2a0e0003;
      23211: inst = 32'h294f0002;
      23212: inst = 32'h11200000;
      23213: inst = 32'hd205ab1;
      23214: inst = 32'h13e00000;
      23215: inst = 32'hfe0aa19;
      23216: inst = 32'h5be00000;
      23217: inst = 32'h244c8000;
      23218: inst = 32'h24428800;
      23219: inst = 32'h8620000;
      23220: inst = 32'h2a0e0004;
      23221: inst = 32'h294f0002;
      23222: inst = 32'h11200000;
      23223: inst = 32'hd205abb;
      23224: inst = 32'h13e00000;
      23225: inst = 32'hfe0aa19;
      23226: inst = 32'h5be00000;
      23227: inst = 32'h244c8000;
      23228: inst = 32'h24428800;
      23229: inst = 32'h8620000;
      23230: inst = 32'h2a0e0005;
      23231: inst = 32'h294f0002;
      23232: inst = 32'h11200000;
      23233: inst = 32'hd205ac5;
      23234: inst = 32'h13e00000;
      23235: inst = 32'hfe0aa19;
      23236: inst = 32'h5be00000;
      23237: inst = 32'h244c8000;
      23238: inst = 32'h24428800;
      23239: inst = 32'h8620000;
      23240: inst = 32'h2a0e0006;
      23241: inst = 32'h294f0002;
      23242: inst = 32'h11200000;
      23243: inst = 32'hd205acf;
      23244: inst = 32'h13e00000;
      23245: inst = 32'hfe0aa19;
      23246: inst = 32'h5be00000;
      23247: inst = 32'h244c8000;
      23248: inst = 32'h24428800;
      23249: inst = 32'h8620000;
      23250: inst = 32'h2a0e0007;
      23251: inst = 32'h294f0002;
      23252: inst = 32'h11200000;
      23253: inst = 32'hd205ad9;
      23254: inst = 32'h13e00000;
      23255: inst = 32'hfe0aa19;
      23256: inst = 32'h5be00000;
      23257: inst = 32'h244c8000;
      23258: inst = 32'h24428800;
      23259: inst = 32'h8620000;
      23260: inst = 32'h2a0e0008;
      23261: inst = 32'h294f0002;
      23262: inst = 32'h11200000;
      23263: inst = 32'hd205ae3;
      23264: inst = 32'h13e00000;
      23265: inst = 32'hfe0aa19;
      23266: inst = 32'h5be00000;
      23267: inst = 32'h244c8000;
      23268: inst = 32'h24428800;
      23269: inst = 32'h8620000;
      23270: inst = 32'h2a0e0009;
      23271: inst = 32'h294f0002;
      23272: inst = 32'h11200000;
      23273: inst = 32'hd205aed;
      23274: inst = 32'h13e00000;
      23275: inst = 32'hfe0aa19;
      23276: inst = 32'h5be00000;
      23277: inst = 32'h244c8000;
      23278: inst = 32'h24428800;
      23279: inst = 32'h8620000;
      23280: inst = 32'h2a0e0002;
      23281: inst = 32'h294f0005;
      23282: inst = 32'h11200000;
      23283: inst = 32'hd205af7;
      23284: inst = 32'h13e00000;
      23285: inst = 32'hfe0aa19;
      23286: inst = 32'h5be00000;
      23287: inst = 32'h244c8000;
      23288: inst = 32'h24428800;
      23289: inst = 32'h8620000;
      23290: inst = 32'h2a0e0002;
      23291: inst = 32'h294f0006;
      23292: inst = 32'h11200000;
      23293: inst = 32'hd205b01;
      23294: inst = 32'h13e00000;
      23295: inst = 32'hfe0aa19;
      23296: inst = 32'h5be00000;
      23297: inst = 32'h244c8000;
      23298: inst = 32'h24428800;
      23299: inst = 32'h8620000;
      23300: inst = 32'h2a0e0003;
      23301: inst = 32'h294f000b;
      23302: inst = 32'h11200000;
      23303: inst = 32'hd205b0b;
      23304: inst = 32'h13e00000;
      23305: inst = 32'hfe0aa19;
      23306: inst = 32'h5be00000;
      23307: inst = 32'h244c8000;
      23308: inst = 32'h24428800;
      23309: inst = 32'h8620000;
      23310: inst = 32'h2a0e0006;
      23311: inst = 32'h294f000b;
      23312: inst = 32'h11200000;
      23313: inst = 32'hd205b15;
      23314: inst = 32'h13e00000;
      23315: inst = 32'hfe0aa19;
      23316: inst = 32'h5be00000;
      23317: inst = 32'h244c8000;
      23318: inst = 32'h24428800;
      23319: inst = 32'h8620000;
      23320: inst = 32'hc60f4ce;
      23321: inst = 32'h2a0e0001;
      23322: inst = 32'h294f0003;
      23323: inst = 32'h11200000;
      23324: inst = 32'hd205b20;
      23325: inst = 32'h13e00000;
      23326: inst = 32'hfe0aa19;
      23327: inst = 32'h5be00000;
      23328: inst = 32'h244c8000;
      23329: inst = 32'h24428800;
      23330: inst = 32'h8620000;
      23331: inst = 32'h2a0e0002;
      23332: inst = 32'h294f0003;
      23333: inst = 32'h11200000;
      23334: inst = 32'hd205b2a;
      23335: inst = 32'h13e00000;
      23336: inst = 32'hfe0aa19;
      23337: inst = 32'h5be00000;
      23338: inst = 32'h244c8000;
      23339: inst = 32'h24428800;
      23340: inst = 32'h8620000;
      23341: inst = 32'h2a0e0003;
      23342: inst = 32'h294f0003;
      23343: inst = 32'h11200000;
      23344: inst = 32'hd205b34;
      23345: inst = 32'h13e00000;
      23346: inst = 32'hfe0aa19;
      23347: inst = 32'h5be00000;
      23348: inst = 32'h244c8000;
      23349: inst = 32'h24428800;
      23350: inst = 32'h8620000;
      23351: inst = 32'h2a0e0004;
      23352: inst = 32'h294f0003;
      23353: inst = 32'h11200000;
      23354: inst = 32'hd205b3e;
      23355: inst = 32'h13e00000;
      23356: inst = 32'hfe0aa19;
      23357: inst = 32'h5be00000;
      23358: inst = 32'h244c8000;
      23359: inst = 32'h24428800;
      23360: inst = 32'h8620000;
      23361: inst = 32'h2a0e0005;
      23362: inst = 32'h294f0003;
      23363: inst = 32'h11200000;
      23364: inst = 32'hd205b48;
      23365: inst = 32'h13e00000;
      23366: inst = 32'hfe0aa19;
      23367: inst = 32'h5be00000;
      23368: inst = 32'h244c8000;
      23369: inst = 32'h24428800;
      23370: inst = 32'h8620000;
      23371: inst = 32'h2a0e0006;
      23372: inst = 32'h294f0003;
      23373: inst = 32'h11200000;
      23374: inst = 32'hd205b52;
      23375: inst = 32'h13e00000;
      23376: inst = 32'hfe0aa19;
      23377: inst = 32'h5be00000;
      23378: inst = 32'h244c8000;
      23379: inst = 32'h24428800;
      23380: inst = 32'h8620000;
      23381: inst = 32'h2a0e0007;
      23382: inst = 32'h294f0003;
      23383: inst = 32'h11200000;
      23384: inst = 32'hd205b5c;
      23385: inst = 32'h13e00000;
      23386: inst = 32'hfe0aa19;
      23387: inst = 32'h5be00000;
      23388: inst = 32'h244c8000;
      23389: inst = 32'h24428800;
      23390: inst = 32'h8620000;
      23391: inst = 32'h2a0e0009;
      23392: inst = 32'h294f0003;
      23393: inst = 32'h11200000;
      23394: inst = 32'hd205b66;
      23395: inst = 32'h13e00000;
      23396: inst = 32'hfe0aa19;
      23397: inst = 32'h5be00000;
      23398: inst = 32'h244c8000;
      23399: inst = 32'h24428800;
      23400: inst = 32'h8620000;
      23401: inst = 32'h2a0e0001;
      23402: inst = 32'h294f0004;
      23403: inst = 32'h11200000;
      23404: inst = 32'hd205b70;
      23405: inst = 32'h13e00000;
      23406: inst = 32'hfe0aa19;
      23407: inst = 32'h5be00000;
      23408: inst = 32'h244c8000;
      23409: inst = 32'h24428800;
      23410: inst = 32'h8620000;
      23411: inst = 32'h2a0e0002;
      23412: inst = 32'h294f0004;
      23413: inst = 32'h11200000;
      23414: inst = 32'hd205b7a;
      23415: inst = 32'h13e00000;
      23416: inst = 32'hfe0aa19;
      23417: inst = 32'h5be00000;
      23418: inst = 32'h244c8000;
      23419: inst = 32'h24428800;
      23420: inst = 32'h8620000;
      23421: inst = 32'h2a0e0003;
      23422: inst = 32'h294f0004;
      23423: inst = 32'h11200000;
      23424: inst = 32'hd205b84;
      23425: inst = 32'h13e00000;
      23426: inst = 32'hfe0aa19;
      23427: inst = 32'h5be00000;
      23428: inst = 32'h244c8000;
      23429: inst = 32'h24428800;
      23430: inst = 32'h8620000;
      23431: inst = 32'h2a0e0004;
      23432: inst = 32'h294f0004;
      23433: inst = 32'h11200000;
      23434: inst = 32'hd205b8e;
      23435: inst = 32'h13e00000;
      23436: inst = 32'hfe0aa19;
      23437: inst = 32'h5be00000;
      23438: inst = 32'h244c8000;
      23439: inst = 32'h24428800;
      23440: inst = 32'h8620000;
      23441: inst = 32'h2a0e0005;
      23442: inst = 32'h294f0004;
      23443: inst = 32'h11200000;
      23444: inst = 32'hd205b98;
      23445: inst = 32'h13e00000;
      23446: inst = 32'hfe0aa19;
      23447: inst = 32'h5be00000;
      23448: inst = 32'h244c8000;
      23449: inst = 32'h24428800;
      23450: inst = 32'h8620000;
      23451: inst = 32'h2a0e0006;
      23452: inst = 32'h294f0004;
      23453: inst = 32'h11200000;
      23454: inst = 32'hd205ba2;
      23455: inst = 32'h13e00000;
      23456: inst = 32'hfe0aa19;
      23457: inst = 32'h5be00000;
      23458: inst = 32'h244c8000;
      23459: inst = 32'h24428800;
      23460: inst = 32'h8620000;
      23461: inst = 32'h2a0e0007;
      23462: inst = 32'h294f0004;
      23463: inst = 32'h11200000;
      23464: inst = 32'hd205bac;
      23465: inst = 32'h13e00000;
      23466: inst = 32'hfe0aa19;
      23467: inst = 32'h5be00000;
      23468: inst = 32'h244c8000;
      23469: inst = 32'h24428800;
      23470: inst = 32'h8620000;
      23471: inst = 32'h2a0e0009;
      23472: inst = 32'h294f0004;
      23473: inst = 32'h11200000;
      23474: inst = 32'hd205bb6;
      23475: inst = 32'h13e00000;
      23476: inst = 32'hfe0aa19;
      23477: inst = 32'h5be00000;
      23478: inst = 32'h244c8000;
      23479: inst = 32'h24428800;
      23480: inst = 32'h8620000;
      23481: inst = 32'h2a0e0003;
      23482: inst = 32'h294f0005;
      23483: inst = 32'h11200000;
      23484: inst = 32'hd205bc0;
      23485: inst = 32'h13e00000;
      23486: inst = 32'hfe0aa19;
      23487: inst = 32'h5be00000;
      23488: inst = 32'h244c8000;
      23489: inst = 32'h24428800;
      23490: inst = 32'h8620000;
      23491: inst = 32'h2a0e0004;
      23492: inst = 32'h294f0005;
      23493: inst = 32'h11200000;
      23494: inst = 32'hd205bca;
      23495: inst = 32'h13e00000;
      23496: inst = 32'hfe0aa19;
      23497: inst = 32'h5be00000;
      23498: inst = 32'h244c8000;
      23499: inst = 32'h24428800;
      23500: inst = 32'h8620000;
      23501: inst = 32'h2a0e0005;
      23502: inst = 32'h294f0005;
      23503: inst = 32'h11200000;
      23504: inst = 32'hd205bd4;
      23505: inst = 32'h13e00000;
      23506: inst = 32'hfe0aa19;
      23507: inst = 32'h5be00000;
      23508: inst = 32'h244c8000;
      23509: inst = 32'h24428800;
      23510: inst = 32'h8620000;
      23511: inst = 32'h2a0e0006;
      23512: inst = 32'h294f0005;
      23513: inst = 32'h11200000;
      23514: inst = 32'hd205bde;
      23515: inst = 32'h13e00000;
      23516: inst = 32'hfe0aa19;
      23517: inst = 32'h5be00000;
      23518: inst = 32'h244c8000;
      23519: inst = 32'h24428800;
      23520: inst = 32'h8620000;
      23521: inst = 32'h2a0e0007;
      23522: inst = 32'h294f0005;
      23523: inst = 32'h11200000;
      23524: inst = 32'hd205be8;
      23525: inst = 32'h13e00000;
      23526: inst = 32'hfe0aa19;
      23527: inst = 32'h5be00000;
      23528: inst = 32'h244c8000;
      23529: inst = 32'h24428800;
      23530: inst = 32'h8620000;
      23531: inst = 32'h2a0e0008;
      23532: inst = 32'h294f0005;
      23533: inst = 32'h11200000;
      23534: inst = 32'hd205bf2;
      23535: inst = 32'h13e00000;
      23536: inst = 32'hfe0aa19;
      23537: inst = 32'h5be00000;
      23538: inst = 32'h244c8000;
      23539: inst = 32'h24428800;
      23540: inst = 32'h8620000;
      23541: inst = 32'h2a0e0009;
      23542: inst = 32'h294f0005;
      23543: inst = 32'h11200000;
      23544: inst = 32'hd205bfc;
      23545: inst = 32'h13e00000;
      23546: inst = 32'hfe0aa19;
      23547: inst = 32'h5be00000;
      23548: inst = 32'h244c8000;
      23549: inst = 32'h24428800;
      23550: inst = 32'h8620000;
      23551: inst = 32'h2a0e0003;
      23552: inst = 32'h294f0006;
      23553: inst = 32'h11200000;
      23554: inst = 32'hd205c06;
      23555: inst = 32'h13e00000;
      23556: inst = 32'hfe0aa19;
      23557: inst = 32'h5be00000;
      23558: inst = 32'h244c8000;
      23559: inst = 32'h24428800;
      23560: inst = 32'h8620000;
      23561: inst = 32'h2a0e0004;
      23562: inst = 32'h294f0006;
      23563: inst = 32'h11200000;
      23564: inst = 32'hd205c10;
      23565: inst = 32'h13e00000;
      23566: inst = 32'hfe0aa19;
      23567: inst = 32'h5be00000;
      23568: inst = 32'h244c8000;
      23569: inst = 32'h24428800;
      23570: inst = 32'h8620000;
      23571: inst = 32'h2a0e0005;
      23572: inst = 32'h294f0006;
      23573: inst = 32'h11200000;
      23574: inst = 32'hd205c1a;
      23575: inst = 32'h13e00000;
      23576: inst = 32'hfe0aa19;
      23577: inst = 32'h5be00000;
      23578: inst = 32'h244c8000;
      23579: inst = 32'h24428800;
      23580: inst = 32'h8620000;
      23581: inst = 32'h2a0e0006;
      23582: inst = 32'h294f0006;
      23583: inst = 32'h11200000;
      23584: inst = 32'hd205c24;
      23585: inst = 32'h13e00000;
      23586: inst = 32'hfe0aa19;
      23587: inst = 32'h5be00000;
      23588: inst = 32'h244c8000;
      23589: inst = 32'h24428800;
      23590: inst = 32'h8620000;
      23591: inst = 32'h2a0e0007;
      23592: inst = 32'h294f0006;
      23593: inst = 32'h11200000;
      23594: inst = 32'hd205c2e;
      23595: inst = 32'h13e00000;
      23596: inst = 32'hfe0aa19;
      23597: inst = 32'h5be00000;
      23598: inst = 32'h244c8000;
      23599: inst = 32'h24428800;
      23600: inst = 32'h8620000;
      23601: inst = 32'h2a0e0008;
      23602: inst = 32'h294f0006;
      23603: inst = 32'h11200000;
      23604: inst = 32'hd205c38;
      23605: inst = 32'h13e00000;
      23606: inst = 32'hfe0aa19;
      23607: inst = 32'h5be00000;
      23608: inst = 32'h244c8000;
      23609: inst = 32'h24428800;
      23610: inst = 32'h8620000;
      23611: inst = 32'h2a0e0009;
      23612: inst = 32'h294f0006;
      23613: inst = 32'h11200000;
      23614: inst = 32'hd205c42;
      23615: inst = 32'h13e00000;
      23616: inst = 32'hfe0aa19;
      23617: inst = 32'h5be00000;
      23618: inst = 32'h244c8000;
      23619: inst = 32'h24428800;
      23620: inst = 32'h8620000;
      23621: inst = 32'h2a0e0004;
      23622: inst = 32'h294f0008;
      23623: inst = 32'h11200000;
      23624: inst = 32'hd205c4c;
      23625: inst = 32'h13e00000;
      23626: inst = 32'hfe0aa19;
      23627: inst = 32'h5be00000;
      23628: inst = 32'h244c8000;
      23629: inst = 32'h24428800;
      23630: inst = 32'h8620000;
      23631: inst = 32'h2a0e0008;
      23632: inst = 32'h294f0008;
      23633: inst = 32'h11200000;
      23634: inst = 32'hd205c56;
      23635: inst = 32'h13e00000;
      23636: inst = 32'hfe0aa19;
      23637: inst = 32'h5be00000;
      23638: inst = 32'h244c8000;
      23639: inst = 32'h24428800;
      23640: inst = 32'h8620000;
      23641: inst = 32'h2a0e0004;
      23642: inst = 32'h294f0009;
      23643: inst = 32'h11200000;
      23644: inst = 32'hd205c60;
      23645: inst = 32'h13e00000;
      23646: inst = 32'hfe0aa19;
      23647: inst = 32'h5be00000;
      23648: inst = 32'h244c8000;
      23649: inst = 32'h24428800;
      23650: inst = 32'h8620000;
      23651: inst = 32'hc607841;
      23652: inst = 32'h2a0e0002;
      23653: inst = 32'h294f0007;
      23654: inst = 32'h11200000;
      23655: inst = 32'hd205c6b;
      23656: inst = 32'h13e00000;
      23657: inst = 32'hfe0aa19;
      23658: inst = 32'h5be00000;
      23659: inst = 32'h244c8000;
      23660: inst = 32'h24428800;
      23661: inst = 32'h8620000;
      23662: inst = 32'h2a0e0002;
      23663: inst = 32'h294f0008;
      23664: inst = 32'h11200000;
      23665: inst = 32'hd205c75;
      23666: inst = 32'h13e00000;
      23667: inst = 32'hfe0aa19;
      23668: inst = 32'h5be00000;
      23669: inst = 32'h244c8000;
      23670: inst = 32'h24428800;
      23671: inst = 32'h8620000;
      23672: inst = 32'hc60a000;
      23673: inst = 32'h2a0e0003;
      23674: inst = 32'h294f0007;
      23675: inst = 32'h11200000;
      23676: inst = 32'hd205c80;
      23677: inst = 32'h13e00000;
      23678: inst = 32'hfe0aa19;
      23679: inst = 32'h5be00000;
      23680: inst = 32'h244c8000;
      23681: inst = 32'h24428800;
      23682: inst = 32'h8620000;
      23683: inst = 32'h2a0e0004;
      23684: inst = 32'h294f0007;
      23685: inst = 32'h11200000;
      23686: inst = 32'hd205c8a;
      23687: inst = 32'h13e00000;
      23688: inst = 32'hfe0aa19;
      23689: inst = 32'h5be00000;
      23690: inst = 32'h244c8000;
      23691: inst = 32'h24428800;
      23692: inst = 32'h8620000;
      23693: inst = 32'h2a0e0005;
      23694: inst = 32'h294f0007;
      23695: inst = 32'h11200000;
      23696: inst = 32'hd205c94;
      23697: inst = 32'h13e00000;
      23698: inst = 32'hfe0aa19;
      23699: inst = 32'h5be00000;
      23700: inst = 32'h244c8000;
      23701: inst = 32'h24428800;
      23702: inst = 32'h8620000;
      23703: inst = 32'h2a0e0006;
      23704: inst = 32'h294f0007;
      23705: inst = 32'h11200000;
      23706: inst = 32'hd205c9e;
      23707: inst = 32'h13e00000;
      23708: inst = 32'hfe0aa19;
      23709: inst = 32'h5be00000;
      23710: inst = 32'h244c8000;
      23711: inst = 32'h24428800;
      23712: inst = 32'h8620000;
      23713: inst = 32'h2a0e0007;
      23714: inst = 32'h294f0007;
      23715: inst = 32'h11200000;
      23716: inst = 32'hd205ca8;
      23717: inst = 32'h13e00000;
      23718: inst = 32'hfe0aa19;
      23719: inst = 32'h5be00000;
      23720: inst = 32'h244c8000;
      23721: inst = 32'h24428800;
      23722: inst = 32'h8620000;
      23723: inst = 32'h2a0e0003;
      23724: inst = 32'h294f0008;
      23725: inst = 32'h11200000;
      23726: inst = 32'hd205cb2;
      23727: inst = 32'h13e00000;
      23728: inst = 32'hfe0aa19;
      23729: inst = 32'h5be00000;
      23730: inst = 32'h244c8000;
      23731: inst = 32'h24428800;
      23732: inst = 32'h8620000;
      23733: inst = 32'h2a0e0005;
      23734: inst = 32'h294f0008;
      23735: inst = 32'h11200000;
      23736: inst = 32'hd205cbc;
      23737: inst = 32'h13e00000;
      23738: inst = 32'hfe0aa19;
      23739: inst = 32'h5be00000;
      23740: inst = 32'h244c8000;
      23741: inst = 32'h24428800;
      23742: inst = 32'h8620000;
      23743: inst = 32'h2a0e0006;
      23744: inst = 32'h294f0008;
      23745: inst = 32'h11200000;
      23746: inst = 32'hd205cc6;
      23747: inst = 32'h13e00000;
      23748: inst = 32'hfe0aa19;
      23749: inst = 32'h5be00000;
      23750: inst = 32'h244c8000;
      23751: inst = 32'h24428800;
      23752: inst = 32'h8620000;
      23753: inst = 32'h2a0e0007;
      23754: inst = 32'h294f0008;
      23755: inst = 32'h11200000;
      23756: inst = 32'hd205cd0;
      23757: inst = 32'h13e00000;
      23758: inst = 32'hfe0aa19;
      23759: inst = 32'h5be00000;
      23760: inst = 32'h244c8000;
      23761: inst = 32'h24428800;
      23762: inst = 32'h8620000;
      23763: inst = 32'h2a0e0002;
      23764: inst = 32'h294f0009;
      23765: inst = 32'h11200000;
      23766: inst = 32'hd205cda;
      23767: inst = 32'h13e00000;
      23768: inst = 32'hfe0aa19;
      23769: inst = 32'h5be00000;
      23770: inst = 32'h244c8000;
      23771: inst = 32'h24428800;
      23772: inst = 32'h8620000;
      23773: inst = 32'h2a0e0003;
      23774: inst = 32'h294f0009;
      23775: inst = 32'h11200000;
      23776: inst = 32'hd205ce4;
      23777: inst = 32'h13e00000;
      23778: inst = 32'hfe0aa19;
      23779: inst = 32'h5be00000;
      23780: inst = 32'h244c8000;
      23781: inst = 32'h24428800;
      23782: inst = 32'h8620000;
      23783: inst = 32'h2a0e0005;
      23784: inst = 32'h294f0009;
      23785: inst = 32'h11200000;
      23786: inst = 32'hd205cee;
      23787: inst = 32'h13e00000;
      23788: inst = 32'hfe0aa19;
      23789: inst = 32'h5be00000;
      23790: inst = 32'h244c8000;
      23791: inst = 32'h24428800;
      23792: inst = 32'h8620000;
      23793: inst = 32'h2a0e0006;
      23794: inst = 32'h294f0009;
      23795: inst = 32'h11200000;
      23796: inst = 32'hd205cf8;
      23797: inst = 32'h13e00000;
      23798: inst = 32'hfe0aa19;
      23799: inst = 32'h5be00000;
      23800: inst = 32'h244c8000;
      23801: inst = 32'h24428800;
      23802: inst = 32'h8620000;
      23803: inst = 32'h2a0e0007;
      23804: inst = 32'h294f0009;
      23805: inst = 32'h11200000;
      23806: inst = 32'hd205d02;
      23807: inst = 32'h13e00000;
      23808: inst = 32'hfe0aa19;
      23809: inst = 32'h5be00000;
      23810: inst = 32'h244c8000;
      23811: inst = 32'h24428800;
      23812: inst = 32'h8620000;
      23813: inst = 32'hc6010ac;
      23814: inst = 32'h2a0e0002;
      23815: inst = 32'h294f000a;
      23816: inst = 32'h11200000;
      23817: inst = 32'hd205d0d;
      23818: inst = 32'h13e00000;
      23819: inst = 32'hfe0aa19;
      23820: inst = 32'h5be00000;
      23821: inst = 32'h244c8000;
      23822: inst = 32'h24428800;
      23823: inst = 32'h8620000;
      23824: inst = 32'h2a0e0003;
      23825: inst = 32'h294f000a;
      23826: inst = 32'h11200000;
      23827: inst = 32'hd205d17;
      23828: inst = 32'h13e00000;
      23829: inst = 32'hfe0aa19;
      23830: inst = 32'h5be00000;
      23831: inst = 32'h244c8000;
      23832: inst = 32'h24428800;
      23833: inst = 32'h8620000;
      23834: inst = 32'h2a0e0004;
      23835: inst = 32'h294f000a;
      23836: inst = 32'h11200000;
      23837: inst = 32'hd205d21;
      23838: inst = 32'h13e00000;
      23839: inst = 32'hfe0aa19;
      23840: inst = 32'h5be00000;
      23841: inst = 32'h244c8000;
      23842: inst = 32'h24428800;
      23843: inst = 32'h8620000;
      23844: inst = 32'h2a0e0005;
      23845: inst = 32'h294f000a;
      23846: inst = 32'h11200000;
      23847: inst = 32'hd205d2b;
      23848: inst = 32'h13e00000;
      23849: inst = 32'hfe0aa19;
      23850: inst = 32'h5be00000;
      23851: inst = 32'h244c8000;
      23852: inst = 32'h24428800;
      23853: inst = 32'h8620000;
      23854: inst = 32'h2a0e0006;
      23855: inst = 32'h294f000a;
      23856: inst = 32'h11200000;
      23857: inst = 32'hd205d35;
      23858: inst = 32'h13e00000;
      23859: inst = 32'hfe0aa19;
      23860: inst = 32'h5be00000;
      23861: inst = 32'h244c8000;
      23862: inst = 32'h24428800;
      23863: inst = 32'h8620000;
      23864: inst = 32'h2a0e0007;
      23865: inst = 32'h294f000a;
      23866: inst = 32'h11200000;
      23867: inst = 32'hd205d3f;
      23868: inst = 32'h13e00000;
      23869: inst = 32'hfe0aa19;
      23870: inst = 32'h5be00000;
      23871: inst = 32'h244c8000;
      23872: inst = 32'h24428800;
      23873: inst = 32'h8620000;
      23874: inst = 32'h13e00000;
      23875: inst = 32'hfe05d49;
      23876: inst = 32'h20200003;
      23877: inst = 32'h5be00000;
      23878: inst = 32'h13e00000;
      23879: inst = 32'hfe06126;
      23880: inst = 32'h5be00000;
      23881: inst = 32'h13e00000;
      23882: inst = 32'hfe06126;
      23883: inst = 32'h5be00000;
      23884: inst = 32'hc6018c3;
      23885: inst = 32'h2a0e000a;
      23886: inst = 32'h294f0000;
      23887: inst = 32'h11200000;
      23888: inst = 32'hd205d54;
      23889: inst = 32'h13e00000;
      23890: inst = 32'hfe0aa19;
      23891: inst = 32'h5be00000;
      23892: inst = 32'h244c8000;
      23893: inst = 32'h24428800;
      23894: inst = 32'h8620000;
      23895: inst = 32'h2a0e0009;
      23896: inst = 32'h294f0000;
      23897: inst = 32'h11200000;
      23898: inst = 32'hd205d5e;
      23899: inst = 32'h13e00000;
      23900: inst = 32'hfe0aa19;
      23901: inst = 32'h5be00000;
      23902: inst = 32'h244c8000;
      23903: inst = 32'h24428800;
      23904: inst = 32'h8620000;
      23905: inst = 32'h2a0e0008;
      23906: inst = 32'h294f0000;
      23907: inst = 32'h11200000;
      23908: inst = 32'hd205d68;
      23909: inst = 32'h13e00000;
      23910: inst = 32'hfe0aa19;
      23911: inst = 32'h5be00000;
      23912: inst = 32'h244c8000;
      23913: inst = 32'h24428800;
      23914: inst = 32'h8620000;
      23915: inst = 32'h2a0e0007;
      23916: inst = 32'h294f0000;
      23917: inst = 32'h11200000;
      23918: inst = 32'hd205d72;
      23919: inst = 32'h13e00000;
      23920: inst = 32'hfe0aa19;
      23921: inst = 32'h5be00000;
      23922: inst = 32'h244c8000;
      23923: inst = 32'h24428800;
      23924: inst = 32'h8620000;
      23925: inst = 32'h2a0e0006;
      23926: inst = 32'h294f0000;
      23927: inst = 32'h11200000;
      23928: inst = 32'hd205d7c;
      23929: inst = 32'h13e00000;
      23930: inst = 32'hfe0aa19;
      23931: inst = 32'h5be00000;
      23932: inst = 32'h244c8000;
      23933: inst = 32'h24428800;
      23934: inst = 32'h8620000;
      23935: inst = 32'h2a0e0005;
      23936: inst = 32'h294f0000;
      23937: inst = 32'h11200000;
      23938: inst = 32'hd205d86;
      23939: inst = 32'h13e00000;
      23940: inst = 32'hfe0aa19;
      23941: inst = 32'h5be00000;
      23942: inst = 32'h244c8000;
      23943: inst = 32'h24428800;
      23944: inst = 32'h8620000;
      23945: inst = 32'h2a0e0004;
      23946: inst = 32'h294f0000;
      23947: inst = 32'h11200000;
      23948: inst = 32'hd205d90;
      23949: inst = 32'h13e00000;
      23950: inst = 32'hfe0aa19;
      23951: inst = 32'h5be00000;
      23952: inst = 32'h244c8000;
      23953: inst = 32'h24428800;
      23954: inst = 32'h8620000;
      23955: inst = 32'h2a0e0003;
      23956: inst = 32'h294f0000;
      23957: inst = 32'h11200000;
      23958: inst = 32'hd205d9a;
      23959: inst = 32'h13e00000;
      23960: inst = 32'hfe0aa19;
      23961: inst = 32'h5be00000;
      23962: inst = 32'h244c8000;
      23963: inst = 32'h24428800;
      23964: inst = 32'h8620000;
      23965: inst = 32'h2a0e0002;
      23966: inst = 32'h294f0000;
      23967: inst = 32'h11200000;
      23968: inst = 32'hd205da4;
      23969: inst = 32'h13e00000;
      23970: inst = 32'hfe0aa19;
      23971: inst = 32'h5be00000;
      23972: inst = 32'h244c8000;
      23973: inst = 32'h24428800;
      23974: inst = 32'h8620000;
      23975: inst = 32'h2a0e0001;
      23976: inst = 32'h294f0000;
      23977: inst = 32'h11200000;
      23978: inst = 32'hd205dae;
      23979: inst = 32'h13e00000;
      23980: inst = 32'hfe0aa19;
      23981: inst = 32'h5be00000;
      23982: inst = 32'h244c8000;
      23983: inst = 32'h24428800;
      23984: inst = 32'h8620000;
      23985: inst = 32'h2a0e000a;
      23986: inst = 32'h294f0001;
      23987: inst = 32'h11200000;
      23988: inst = 32'hd205db8;
      23989: inst = 32'h13e00000;
      23990: inst = 32'hfe0aa19;
      23991: inst = 32'h5be00000;
      23992: inst = 32'h244c8000;
      23993: inst = 32'h24428800;
      23994: inst = 32'h8620000;
      23995: inst = 32'h2a0e0009;
      23996: inst = 32'h294f0001;
      23997: inst = 32'h11200000;
      23998: inst = 32'hd205dc2;
      23999: inst = 32'h13e00000;
      24000: inst = 32'hfe0aa19;
      24001: inst = 32'h5be00000;
      24002: inst = 32'h244c8000;
      24003: inst = 32'h24428800;
      24004: inst = 32'h8620000;
      24005: inst = 32'h2a0e0008;
      24006: inst = 32'h294f0001;
      24007: inst = 32'h11200000;
      24008: inst = 32'hd205dcc;
      24009: inst = 32'h13e00000;
      24010: inst = 32'hfe0aa19;
      24011: inst = 32'h5be00000;
      24012: inst = 32'h244c8000;
      24013: inst = 32'h24428800;
      24014: inst = 32'h8620000;
      24015: inst = 32'h2a0e0007;
      24016: inst = 32'h294f0001;
      24017: inst = 32'h11200000;
      24018: inst = 32'hd205dd6;
      24019: inst = 32'h13e00000;
      24020: inst = 32'hfe0aa19;
      24021: inst = 32'h5be00000;
      24022: inst = 32'h244c8000;
      24023: inst = 32'h24428800;
      24024: inst = 32'h8620000;
      24025: inst = 32'h2a0e0006;
      24026: inst = 32'h294f0001;
      24027: inst = 32'h11200000;
      24028: inst = 32'hd205de0;
      24029: inst = 32'h13e00000;
      24030: inst = 32'hfe0aa19;
      24031: inst = 32'h5be00000;
      24032: inst = 32'h244c8000;
      24033: inst = 32'h24428800;
      24034: inst = 32'h8620000;
      24035: inst = 32'h2a0e0005;
      24036: inst = 32'h294f0001;
      24037: inst = 32'h11200000;
      24038: inst = 32'hd205dea;
      24039: inst = 32'h13e00000;
      24040: inst = 32'hfe0aa19;
      24041: inst = 32'h5be00000;
      24042: inst = 32'h244c8000;
      24043: inst = 32'h24428800;
      24044: inst = 32'h8620000;
      24045: inst = 32'h2a0e0004;
      24046: inst = 32'h294f0001;
      24047: inst = 32'h11200000;
      24048: inst = 32'hd205df4;
      24049: inst = 32'h13e00000;
      24050: inst = 32'hfe0aa19;
      24051: inst = 32'h5be00000;
      24052: inst = 32'h244c8000;
      24053: inst = 32'h24428800;
      24054: inst = 32'h8620000;
      24055: inst = 32'h2a0e0003;
      24056: inst = 32'h294f0001;
      24057: inst = 32'h11200000;
      24058: inst = 32'hd205dfe;
      24059: inst = 32'h13e00000;
      24060: inst = 32'hfe0aa19;
      24061: inst = 32'h5be00000;
      24062: inst = 32'h244c8000;
      24063: inst = 32'h24428800;
      24064: inst = 32'h8620000;
      24065: inst = 32'h2a0e0002;
      24066: inst = 32'h294f0001;
      24067: inst = 32'h11200000;
      24068: inst = 32'hd205e08;
      24069: inst = 32'h13e00000;
      24070: inst = 32'hfe0aa19;
      24071: inst = 32'h5be00000;
      24072: inst = 32'h244c8000;
      24073: inst = 32'h24428800;
      24074: inst = 32'h8620000;
      24075: inst = 32'h2a0e0001;
      24076: inst = 32'h294f0001;
      24077: inst = 32'h11200000;
      24078: inst = 32'hd205e12;
      24079: inst = 32'h13e00000;
      24080: inst = 32'hfe0aa19;
      24081: inst = 32'h5be00000;
      24082: inst = 32'h244c8000;
      24083: inst = 32'h24428800;
      24084: inst = 32'h8620000;
      24085: inst = 32'h2a0e000a;
      24086: inst = 32'h294f0002;
      24087: inst = 32'h11200000;
      24088: inst = 32'hd205e1c;
      24089: inst = 32'h13e00000;
      24090: inst = 32'hfe0aa19;
      24091: inst = 32'h5be00000;
      24092: inst = 32'h244c8000;
      24093: inst = 32'h24428800;
      24094: inst = 32'h8620000;
      24095: inst = 32'h2a0e0009;
      24096: inst = 32'h294f0002;
      24097: inst = 32'h11200000;
      24098: inst = 32'hd205e26;
      24099: inst = 32'h13e00000;
      24100: inst = 32'hfe0aa19;
      24101: inst = 32'h5be00000;
      24102: inst = 32'h244c8000;
      24103: inst = 32'h24428800;
      24104: inst = 32'h8620000;
      24105: inst = 32'h2a0e000a;
      24106: inst = 32'h294f0003;
      24107: inst = 32'h11200000;
      24108: inst = 32'hd205e30;
      24109: inst = 32'h13e00000;
      24110: inst = 32'hfe0aa19;
      24111: inst = 32'h5be00000;
      24112: inst = 32'h244c8000;
      24113: inst = 32'h24428800;
      24114: inst = 32'h8620000;
      24115: inst = 32'h2a0e0002;
      24116: inst = 32'h294f0003;
      24117: inst = 32'h11200000;
      24118: inst = 32'hd205e3a;
      24119: inst = 32'h13e00000;
      24120: inst = 32'hfe0aa19;
      24121: inst = 32'h5be00000;
      24122: inst = 32'h244c8000;
      24123: inst = 32'h24428800;
      24124: inst = 32'h8620000;
      24125: inst = 32'h2a0e000a;
      24126: inst = 32'h294f0004;
      24127: inst = 32'h11200000;
      24128: inst = 32'hd205e44;
      24129: inst = 32'h13e00000;
      24130: inst = 32'hfe0aa19;
      24131: inst = 32'h5be00000;
      24132: inst = 32'h244c8000;
      24133: inst = 32'h24428800;
      24134: inst = 32'h8620000;
      24135: inst = 32'h2a0e0002;
      24136: inst = 32'h294f0004;
      24137: inst = 32'h11200000;
      24138: inst = 32'hd205e4e;
      24139: inst = 32'h13e00000;
      24140: inst = 32'hfe0aa19;
      24141: inst = 32'h5be00000;
      24142: inst = 32'h244c8000;
      24143: inst = 32'h24428800;
      24144: inst = 32'h8620000;
      24145: inst = 32'h2a0e000a;
      24146: inst = 32'h294f0005;
      24147: inst = 32'h11200000;
      24148: inst = 32'hd205e58;
      24149: inst = 32'h13e00000;
      24150: inst = 32'hfe0aa19;
      24151: inst = 32'h5be00000;
      24152: inst = 32'h244c8000;
      24153: inst = 32'h24428800;
      24154: inst = 32'h8620000;
      24155: inst = 32'h2a0e0009;
      24156: inst = 32'h294f0005;
      24157: inst = 32'h11200000;
      24158: inst = 32'hd205e62;
      24159: inst = 32'h13e00000;
      24160: inst = 32'hfe0aa19;
      24161: inst = 32'h5be00000;
      24162: inst = 32'h244c8000;
      24163: inst = 32'h24428800;
      24164: inst = 32'h8620000;
      24165: inst = 32'h2a0e000a;
      24166: inst = 32'h294f0006;
      24167: inst = 32'h11200000;
      24168: inst = 32'hd205e6c;
      24169: inst = 32'h13e00000;
      24170: inst = 32'hfe0aa19;
      24171: inst = 32'h5be00000;
      24172: inst = 32'h244c8000;
      24173: inst = 32'h24428800;
      24174: inst = 32'h8620000;
      24175: inst = 32'h2a0e0009;
      24176: inst = 32'h294f0006;
      24177: inst = 32'h11200000;
      24178: inst = 32'hd205e76;
      24179: inst = 32'h13e00000;
      24180: inst = 32'hfe0aa19;
      24181: inst = 32'h5be00000;
      24182: inst = 32'h244c8000;
      24183: inst = 32'h24428800;
      24184: inst = 32'h8620000;
      24185: inst = 32'hc60d42c;
      24186: inst = 32'h2a0e0008;
      24187: inst = 32'h294f0002;
      24188: inst = 32'h11200000;
      24189: inst = 32'hd205e81;
      24190: inst = 32'h13e00000;
      24191: inst = 32'hfe0aa19;
      24192: inst = 32'h5be00000;
      24193: inst = 32'h244c8000;
      24194: inst = 32'h24428800;
      24195: inst = 32'h8620000;
      24196: inst = 32'h2a0e0007;
      24197: inst = 32'h294f0002;
      24198: inst = 32'h11200000;
      24199: inst = 32'hd205e8b;
      24200: inst = 32'h13e00000;
      24201: inst = 32'hfe0aa19;
      24202: inst = 32'h5be00000;
      24203: inst = 32'h244c8000;
      24204: inst = 32'h24428800;
      24205: inst = 32'h8620000;
      24206: inst = 32'h2a0e0006;
      24207: inst = 32'h294f0002;
      24208: inst = 32'h11200000;
      24209: inst = 32'hd205e95;
      24210: inst = 32'h13e00000;
      24211: inst = 32'hfe0aa19;
      24212: inst = 32'h5be00000;
      24213: inst = 32'h244c8000;
      24214: inst = 32'h24428800;
      24215: inst = 32'h8620000;
      24216: inst = 32'h2a0e0005;
      24217: inst = 32'h294f0002;
      24218: inst = 32'h11200000;
      24219: inst = 32'hd205e9f;
      24220: inst = 32'h13e00000;
      24221: inst = 32'hfe0aa19;
      24222: inst = 32'h5be00000;
      24223: inst = 32'h244c8000;
      24224: inst = 32'h24428800;
      24225: inst = 32'h8620000;
      24226: inst = 32'h2a0e0004;
      24227: inst = 32'h294f0002;
      24228: inst = 32'h11200000;
      24229: inst = 32'hd205ea9;
      24230: inst = 32'h13e00000;
      24231: inst = 32'hfe0aa19;
      24232: inst = 32'h5be00000;
      24233: inst = 32'h244c8000;
      24234: inst = 32'h24428800;
      24235: inst = 32'h8620000;
      24236: inst = 32'h2a0e0003;
      24237: inst = 32'h294f0002;
      24238: inst = 32'h11200000;
      24239: inst = 32'hd205eb3;
      24240: inst = 32'h13e00000;
      24241: inst = 32'hfe0aa19;
      24242: inst = 32'h5be00000;
      24243: inst = 32'h244c8000;
      24244: inst = 32'h24428800;
      24245: inst = 32'h8620000;
      24246: inst = 32'h2a0e0002;
      24247: inst = 32'h294f0002;
      24248: inst = 32'h11200000;
      24249: inst = 32'hd205ebd;
      24250: inst = 32'h13e00000;
      24251: inst = 32'hfe0aa19;
      24252: inst = 32'h5be00000;
      24253: inst = 32'h244c8000;
      24254: inst = 32'h24428800;
      24255: inst = 32'h8620000;
      24256: inst = 32'h2a0e0001;
      24257: inst = 32'h294f0002;
      24258: inst = 32'h11200000;
      24259: inst = 32'hd205ec7;
      24260: inst = 32'h13e00000;
      24261: inst = 32'hfe0aa19;
      24262: inst = 32'h5be00000;
      24263: inst = 32'h244c8000;
      24264: inst = 32'h24428800;
      24265: inst = 32'h8620000;
      24266: inst = 32'h2a0e0008;
      24267: inst = 32'h294f0005;
      24268: inst = 32'h11200000;
      24269: inst = 32'hd205ed1;
      24270: inst = 32'h13e00000;
      24271: inst = 32'hfe0aa19;
      24272: inst = 32'h5be00000;
      24273: inst = 32'h244c8000;
      24274: inst = 32'h24428800;
      24275: inst = 32'h8620000;
      24276: inst = 32'h2a0e0008;
      24277: inst = 32'h294f0006;
      24278: inst = 32'h11200000;
      24279: inst = 32'hd205edb;
      24280: inst = 32'h13e00000;
      24281: inst = 32'hfe0aa19;
      24282: inst = 32'h5be00000;
      24283: inst = 32'h244c8000;
      24284: inst = 32'h24428800;
      24285: inst = 32'h8620000;
      24286: inst = 32'h2a0e0007;
      24287: inst = 32'h294f000b;
      24288: inst = 32'h11200000;
      24289: inst = 32'hd205ee5;
      24290: inst = 32'h13e00000;
      24291: inst = 32'hfe0aa19;
      24292: inst = 32'h5be00000;
      24293: inst = 32'h244c8000;
      24294: inst = 32'h24428800;
      24295: inst = 32'h8620000;
      24296: inst = 32'h2a0e0004;
      24297: inst = 32'h294f000b;
      24298: inst = 32'h11200000;
      24299: inst = 32'hd205eef;
      24300: inst = 32'h13e00000;
      24301: inst = 32'hfe0aa19;
      24302: inst = 32'h5be00000;
      24303: inst = 32'h244c8000;
      24304: inst = 32'h24428800;
      24305: inst = 32'h8620000;
      24306: inst = 32'hc60f4ce;
      24307: inst = 32'h2a0e0009;
      24308: inst = 32'h294f0003;
      24309: inst = 32'h11200000;
      24310: inst = 32'hd205efa;
      24311: inst = 32'h13e00000;
      24312: inst = 32'hfe0aa19;
      24313: inst = 32'h5be00000;
      24314: inst = 32'h244c8000;
      24315: inst = 32'h24428800;
      24316: inst = 32'h8620000;
      24317: inst = 32'h2a0e0008;
      24318: inst = 32'h294f0003;
      24319: inst = 32'h11200000;
      24320: inst = 32'hd205f04;
      24321: inst = 32'h13e00000;
      24322: inst = 32'hfe0aa19;
      24323: inst = 32'h5be00000;
      24324: inst = 32'h244c8000;
      24325: inst = 32'h24428800;
      24326: inst = 32'h8620000;
      24327: inst = 32'h2a0e0007;
      24328: inst = 32'h294f0003;
      24329: inst = 32'h11200000;
      24330: inst = 32'hd205f0e;
      24331: inst = 32'h13e00000;
      24332: inst = 32'hfe0aa19;
      24333: inst = 32'h5be00000;
      24334: inst = 32'h244c8000;
      24335: inst = 32'h24428800;
      24336: inst = 32'h8620000;
      24337: inst = 32'h2a0e0006;
      24338: inst = 32'h294f0003;
      24339: inst = 32'h11200000;
      24340: inst = 32'hd205f18;
      24341: inst = 32'h13e00000;
      24342: inst = 32'hfe0aa19;
      24343: inst = 32'h5be00000;
      24344: inst = 32'h244c8000;
      24345: inst = 32'h24428800;
      24346: inst = 32'h8620000;
      24347: inst = 32'h2a0e0005;
      24348: inst = 32'h294f0003;
      24349: inst = 32'h11200000;
      24350: inst = 32'hd205f22;
      24351: inst = 32'h13e00000;
      24352: inst = 32'hfe0aa19;
      24353: inst = 32'h5be00000;
      24354: inst = 32'h244c8000;
      24355: inst = 32'h24428800;
      24356: inst = 32'h8620000;
      24357: inst = 32'h2a0e0004;
      24358: inst = 32'h294f0003;
      24359: inst = 32'h11200000;
      24360: inst = 32'hd205f2c;
      24361: inst = 32'h13e00000;
      24362: inst = 32'hfe0aa19;
      24363: inst = 32'h5be00000;
      24364: inst = 32'h244c8000;
      24365: inst = 32'h24428800;
      24366: inst = 32'h8620000;
      24367: inst = 32'h2a0e0003;
      24368: inst = 32'h294f0003;
      24369: inst = 32'h11200000;
      24370: inst = 32'hd205f36;
      24371: inst = 32'h13e00000;
      24372: inst = 32'hfe0aa19;
      24373: inst = 32'h5be00000;
      24374: inst = 32'h244c8000;
      24375: inst = 32'h24428800;
      24376: inst = 32'h8620000;
      24377: inst = 32'h2a0e0001;
      24378: inst = 32'h294f0003;
      24379: inst = 32'h11200000;
      24380: inst = 32'hd205f40;
      24381: inst = 32'h13e00000;
      24382: inst = 32'hfe0aa19;
      24383: inst = 32'h5be00000;
      24384: inst = 32'h244c8000;
      24385: inst = 32'h24428800;
      24386: inst = 32'h8620000;
      24387: inst = 32'h2a0e0009;
      24388: inst = 32'h294f0004;
      24389: inst = 32'h11200000;
      24390: inst = 32'hd205f4a;
      24391: inst = 32'h13e00000;
      24392: inst = 32'hfe0aa19;
      24393: inst = 32'h5be00000;
      24394: inst = 32'h244c8000;
      24395: inst = 32'h24428800;
      24396: inst = 32'h8620000;
      24397: inst = 32'h2a0e0008;
      24398: inst = 32'h294f0004;
      24399: inst = 32'h11200000;
      24400: inst = 32'hd205f54;
      24401: inst = 32'h13e00000;
      24402: inst = 32'hfe0aa19;
      24403: inst = 32'h5be00000;
      24404: inst = 32'h244c8000;
      24405: inst = 32'h24428800;
      24406: inst = 32'h8620000;
      24407: inst = 32'h2a0e0007;
      24408: inst = 32'h294f0004;
      24409: inst = 32'h11200000;
      24410: inst = 32'hd205f5e;
      24411: inst = 32'h13e00000;
      24412: inst = 32'hfe0aa19;
      24413: inst = 32'h5be00000;
      24414: inst = 32'h244c8000;
      24415: inst = 32'h24428800;
      24416: inst = 32'h8620000;
      24417: inst = 32'h2a0e0006;
      24418: inst = 32'h294f0004;
      24419: inst = 32'h11200000;
      24420: inst = 32'hd205f68;
      24421: inst = 32'h13e00000;
      24422: inst = 32'hfe0aa19;
      24423: inst = 32'h5be00000;
      24424: inst = 32'h244c8000;
      24425: inst = 32'h24428800;
      24426: inst = 32'h8620000;
      24427: inst = 32'h2a0e0005;
      24428: inst = 32'h294f0004;
      24429: inst = 32'h11200000;
      24430: inst = 32'hd205f72;
      24431: inst = 32'h13e00000;
      24432: inst = 32'hfe0aa19;
      24433: inst = 32'h5be00000;
      24434: inst = 32'h244c8000;
      24435: inst = 32'h24428800;
      24436: inst = 32'h8620000;
      24437: inst = 32'h2a0e0004;
      24438: inst = 32'h294f0004;
      24439: inst = 32'h11200000;
      24440: inst = 32'hd205f7c;
      24441: inst = 32'h13e00000;
      24442: inst = 32'hfe0aa19;
      24443: inst = 32'h5be00000;
      24444: inst = 32'h244c8000;
      24445: inst = 32'h24428800;
      24446: inst = 32'h8620000;
      24447: inst = 32'h2a0e0003;
      24448: inst = 32'h294f0004;
      24449: inst = 32'h11200000;
      24450: inst = 32'hd205f86;
      24451: inst = 32'h13e00000;
      24452: inst = 32'hfe0aa19;
      24453: inst = 32'h5be00000;
      24454: inst = 32'h244c8000;
      24455: inst = 32'h24428800;
      24456: inst = 32'h8620000;
      24457: inst = 32'h2a0e0001;
      24458: inst = 32'h294f0004;
      24459: inst = 32'h11200000;
      24460: inst = 32'hd205f90;
      24461: inst = 32'h13e00000;
      24462: inst = 32'hfe0aa19;
      24463: inst = 32'h5be00000;
      24464: inst = 32'h244c8000;
      24465: inst = 32'h24428800;
      24466: inst = 32'h8620000;
      24467: inst = 32'h2a0e0007;
      24468: inst = 32'h294f0005;
      24469: inst = 32'h11200000;
      24470: inst = 32'hd205f9a;
      24471: inst = 32'h13e00000;
      24472: inst = 32'hfe0aa19;
      24473: inst = 32'h5be00000;
      24474: inst = 32'h244c8000;
      24475: inst = 32'h24428800;
      24476: inst = 32'h8620000;
      24477: inst = 32'h2a0e0006;
      24478: inst = 32'h294f0005;
      24479: inst = 32'h11200000;
      24480: inst = 32'hd205fa4;
      24481: inst = 32'h13e00000;
      24482: inst = 32'hfe0aa19;
      24483: inst = 32'h5be00000;
      24484: inst = 32'h244c8000;
      24485: inst = 32'h24428800;
      24486: inst = 32'h8620000;
      24487: inst = 32'h2a0e0005;
      24488: inst = 32'h294f0005;
      24489: inst = 32'h11200000;
      24490: inst = 32'hd205fae;
      24491: inst = 32'h13e00000;
      24492: inst = 32'hfe0aa19;
      24493: inst = 32'h5be00000;
      24494: inst = 32'h244c8000;
      24495: inst = 32'h24428800;
      24496: inst = 32'h8620000;
      24497: inst = 32'h2a0e0004;
      24498: inst = 32'h294f0005;
      24499: inst = 32'h11200000;
      24500: inst = 32'hd205fb8;
      24501: inst = 32'h13e00000;
      24502: inst = 32'hfe0aa19;
      24503: inst = 32'h5be00000;
      24504: inst = 32'h244c8000;
      24505: inst = 32'h24428800;
      24506: inst = 32'h8620000;
      24507: inst = 32'h2a0e0003;
      24508: inst = 32'h294f0005;
      24509: inst = 32'h11200000;
      24510: inst = 32'hd205fc2;
      24511: inst = 32'h13e00000;
      24512: inst = 32'hfe0aa19;
      24513: inst = 32'h5be00000;
      24514: inst = 32'h244c8000;
      24515: inst = 32'h24428800;
      24516: inst = 32'h8620000;
      24517: inst = 32'h2a0e0002;
      24518: inst = 32'h294f0005;
      24519: inst = 32'h11200000;
      24520: inst = 32'hd205fcc;
      24521: inst = 32'h13e00000;
      24522: inst = 32'hfe0aa19;
      24523: inst = 32'h5be00000;
      24524: inst = 32'h244c8000;
      24525: inst = 32'h24428800;
      24526: inst = 32'h8620000;
      24527: inst = 32'h2a0e0001;
      24528: inst = 32'h294f0005;
      24529: inst = 32'h11200000;
      24530: inst = 32'hd205fd6;
      24531: inst = 32'h13e00000;
      24532: inst = 32'hfe0aa19;
      24533: inst = 32'h5be00000;
      24534: inst = 32'h244c8000;
      24535: inst = 32'h24428800;
      24536: inst = 32'h8620000;
      24537: inst = 32'h2a0e0007;
      24538: inst = 32'h294f0006;
      24539: inst = 32'h11200000;
      24540: inst = 32'hd205fe0;
      24541: inst = 32'h13e00000;
      24542: inst = 32'hfe0aa19;
      24543: inst = 32'h5be00000;
      24544: inst = 32'h244c8000;
      24545: inst = 32'h24428800;
      24546: inst = 32'h8620000;
      24547: inst = 32'h2a0e0006;
      24548: inst = 32'h294f0006;
      24549: inst = 32'h11200000;
      24550: inst = 32'hd205fea;
      24551: inst = 32'h13e00000;
      24552: inst = 32'hfe0aa19;
      24553: inst = 32'h5be00000;
      24554: inst = 32'h244c8000;
      24555: inst = 32'h24428800;
      24556: inst = 32'h8620000;
      24557: inst = 32'h2a0e0005;
      24558: inst = 32'h294f0006;
      24559: inst = 32'h11200000;
      24560: inst = 32'hd205ff4;
      24561: inst = 32'h13e00000;
      24562: inst = 32'hfe0aa19;
      24563: inst = 32'h5be00000;
      24564: inst = 32'h244c8000;
      24565: inst = 32'h24428800;
      24566: inst = 32'h8620000;
      24567: inst = 32'h2a0e0004;
      24568: inst = 32'h294f0006;
      24569: inst = 32'h11200000;
      24570: inst = 32'hd205ffe;
      24571: inst = 32'h13e00000;
      24572: inst = 32'hfe0aa19;
      24573: inst = 32'h5be00000;
      24574: inst = 32'h244c8000;
      24575: inst = 32'h24428800;
      24576: inst = 32'h8620000;
      24577: inst = 32'h2a0e0003;
      24578: inst = 32'h294f0006;
      24579: inst = 32'h11200000;
      24580: inst = 32'hd206008;
      24581: inst = 32'h13e00000;
      24582: inst = 32'hfe0aa19;
      24583: inst = 32'h5be00000;
      24584: inst = 32'h244c8000;
      24585: inst = 32'h24428800;
      24586: inst = 32'h8620000;
      24587: inst = 32'h2a0e0002;
      24588: inst = 32'h294f0006;
      24589: inst = 32'h11200000;
      24590: inst = 32'hd206012;
      24591: inst = 32'h13e00000;
      24592: inst = 32'hfe0aa19;
      24593: inst = 32'h5be00000;
      24594: inst = 32'h244c8000;
      24595: inst = 32'h24428800;
      24596: inst = 32'h8620000;
      24597: inst = 32'h2a0e0001;
      24598: inst = 32'h294f0006;
      24599: inst = 32'h11200000;
      24600: inst = 32'hd20601c;
      24601: inst = 32'h13e00000;
      24602: inst = 32'hfe0aa19;
      24603: inst = 32'h5be00000;
      24604: inst = 32'h244c8000;
      24605: inst = 32'h24428800;
      24606: inst = 32'h8620000;
      24607: inst = 32'h2a0e0006;
      24608: inst = 32'h294f0008;
      24609: inst = 32'h11200000;
      24610: inst = 32'hd206026;
      24611: inst = 32'h13e00000;
      24612: inst = 32'hfe0aa19;
      24613: inst = 32'h5be00000;
      24614: inst = 32'h244c8000;
      24615: inst = 32'h24428800;
      24616: inst = 32'h8620000;
      24617: inst = 32'h2a0e0002;
      24618: inst = 32'h294f0008;
      24619: inst = 32'h11200000;
      24620: inst = 32'hd206030;
      24621: inst = 32'h13e00000;
      24622: inst = 32'hfe0aa19;
      24623: inst = 32'h5be00000;
      24624: inst = 32'h244c8000;
      24625: inst = 32'h24428800;
      24626: inst = 32'h8620000;
      24627: inst = 32'h2a0e0006;
      24628: inst = 32'h294f0009;
      24629: inst = 32'h11200000;
      24630: inst = 32'hd20603a;
      24631: inst = 32'h13e00000;
      24632: inst = 32'hfe0aa19;
      24633: inst = 32'h5be00000;
      24634: inst = 32'h244c8000;
      24635: inst = 32'h24428800;
      24636: inst = 32'h8620000;
      24637: inst = 32'hc607841;
      24638: inst = 32'h2a0e0008;
      24639: inst = 32'h294f0007;
      24640: inst = 32'h11200000;
      24641: inst = 32'hd206045;
      24642: inst = 32'h13e00000;
      24643: inst = 32'hfe0aa19;
      24644: inst = 32'h5be00000;
      24645: inst = 32'h244c8000;
      24646: inst = 32'h24428800;
      24647: inst = 32'h8620000;
      24648: inst = 32'h2a0e0008;
      24649: inst = 32'h294f0008;
      24650: inst = 32'h11200000;
      24651: inst = 32'hd20604f;
      24652: inst = 32'h13e00000;
      24653: inst = 32'hfe0aa19;
      24654: inst = 32'h5be00000;
      24655: inst = 32'h244c8000;
      24656: inst = 32'h24428800;
      24657: inst = 32'h8620000;
      24658: inst = 32'hc60a000;
      24659: inst = 32'h2a0e0007;
      24660: inst = 32'h294f0007;
      24661: inst = 32'h11200000;
      24662: inst = 32'hd20605a;
      24663: inst = 32'h13e00000;
      24664: inst = 32'hfe0aa19;
      24665: inst = 32'h5be00000;
      24666: inst = 32'h244c8000;
      24667: inst = 32'h24428800;
      24668: inst = 32'h8620000;
      24669: inst = 32'h2a0e0006;
      24670: inst = 32'h294f0007;
      24671: inst = 32'h11200000;
      24672: inst = 32'hd206064;
      24673: inst = 32'h13e00000;
      24674: inst = 32'hfe0aa19;
      24675: inst = 32'h5be00000;
      24676: inst = 32'h244c8000;
      24677: inst = 32'h24428800;
      24678: inst = 32'h8620000;
      24679: inst = 32'h2a0e0005;
      24680: inst = 32'h294f0007;
      24681: inst = 32'h11200000;
      24682: inst = 32'hd20606e;
      24683: inst = 32'h13e00000;
      24684: inst = 32'hfe0aa19;
      24685: inst = 32'h5be00000;
      24686: inst = 32'h244c8000;
      24687: inst = 32'h24428800;
      24688: inst = 32'h8620000;
      24689: inst = 32'h2a0e0004;
      24690: inst = 32'h294f0007;
      24691: inst = 32'h11200000;
      24692: inst = 32'hd206078;
      24693: inst = 32'h13e00000;
      24694: inst = 32'hfe0aa19;
      24695: inst = 32'h5be00000;
      24696: inst = 32'h244c8000;
      24697: inst = 32'h24428800;
      24698: inst = 32'h8620000;
      24699: inst = 32'h2a0e0003;
      24700: inst = 32'h294f0007;
      24701: inst = 32'h11200000;
      24702: inst = 32'hd206082;
      24703: inst = 32'h13e00000;
      24704: inst = 32'hfe0aa19;
      24705: inst = 32'h5be00000;
      24706: inst = 32'h244c8000;
      24707: inst = 32'h24428800;
      24708: inst = 32'h8620000;
      24709: inst = 32'h2a0e0007;
      24710: inst = 32'h294f0008;
      24711: inst = 32'h11200000;
      24712: inst = 32'hd20608c;
      24713: inst = 32'h13e00000;
      24714: inst = 32'hfe0aa19;
      24715: inst = 32'h5be00000;
      24716: inst = 32'h244c8000;
      24717: inst = 32'h24428800;
      24718: inst = 32'h8620000;
      24719: inst = 32'h2a0e0005;
      24720: inst = 32'h294f0008;
      24721: inst = 32'h11200000;
      24722: inst = 32'hd206096;
      24723: inst = 32'h13e00000;
      24724: inst = 32'hfe0aa19;
      24725: inst = 32'h5be00000;
      24726: inst = 32'h244c8000;
      24727: inst = 32'h24428800;
      24728: inst = 32'h8620000;
      24729: inst = 32'h2a0e0004;
      24730: inst = 32'h294f0008;
      24731: inst = 32'h11200000;
      24732: inst = 32'hd2060a0;
      24733: inst = 32'h13e00000;
      24734: inst = 32'hfe0aa19;
      24735: inst = 32'h5be00000;
      24736: inst = 32'h244c8000;
      24737: inst = 32'h24428800;
      24738: inst = 32'h8620000;
      24739: inst = 32'h2a0e0003;
      24740: inst = 32'h294f0008;
      24741: inst = 32'h11200000;
      24742: inst = 32'hd2060aa;
      24743: inst = 32'h13e00000;
      24744: inst = 32'hfe0aa19;
      24745: inst = 32'h5be00000;
      24746: inst = 32'h244c8000;
      24747: inst = 32'h24428800;
      24748: inst = 32'h8620000;
      24749: inst = 32'h2a0e0008;
      24750: inst = 32'h294f0009;
      24751: inst = 32'h11200000;
      24752: inst = 32'hd2060b4;
      24753: inst = 32'h13e00000;
      24754: inst = 32'hfe0aa19;
      24755: inst = 32'h5be00000;
      24756: inst = 32'h244c8000;
      24757: inst = 32'h24428800;
      24758: inst = 32'h8620000;
      24759: inst = 32'h2a0e0007;
      24760: inst = 32'h294f0009;
      24761: inst = 32'h11200000;
      24762: inst = 32'hd2060be;
      24763: inst = 32'h13e00000;
      24764: inst = 32'hfe0aa19;
      24765: inst = 32'h5be00000;
      24766: inst = 32'h244c8000;
      24767: inst = 32'h24428800;
      24768: inst = 32'h8620000;
      24769: inst = 32'h2a0e0005;
      24770: inst = 32'h294f0009;
      24771: inst = 32'h11200000;
      24772: inst = 32'hd2060c8;
      24773: inst = 32'h13e00000;
      24774: inst = 32'hfe0aa19;
      24775: inst = 32'h5be00000;
      24776: inst = 32'h244c8000;
      24777: inst = 32'h24428800;
      24778: inst = 32'h8620000;
      24779: inst = 32'h2a0e0004;
      24780: inst = 32'h294f0009;
      24781: inst = 32'h11200000;
      24782: inst = 32'hd2060d2;
      24783: inst = 32'h13e00000;
      24784: inst = 32'hfe0aa19;
      24785: inst = 32'h5be00000;
      24786: inst = 32'h244c8000;
      24787: inst = 32'h24428800;
      24788: inst = 32'h8620000;
      24789: inst = 32'h2a0e0003;
      24790: inst = 32'h294f0009;
      24791: inst = 32'h11200000;
      24792: inst = 32'hd2060dc;
      24793: inst = 32'h13e00000;
      24794: inst = 32'hfe0aa19;
      24795: inst = 32'h5be00000;
      24796: inst = 32'h244c8000;
      24797: inst = 32'h24428800;
      24798: inst = 32'h8620000;
      24799: inst = 32'hc6010ac;
      24800: inst = 32'h2a0e0008;
      24801: inst = 32'h294f000a;
      24802: inst = 32'h11200000;
      24803: inst = 32'hd2060e7;
      24804: inst = 32'h13e00000;
      24805: inst = 32'hfe0aa19;
      24806: inst = 32'h5be00000;
      24807: inst = 32'h244c8000;
      24808: inst = 32'h24428800;
      24809: inst = 32'h8620000;
      24810: inst = 32'h2a0e0007;
      24811: inst = 32'h294f000a;
      24812: inst = 32'h11200000;
      24813: inst = 32'hd2060f1;
      24814: inst = 32'h13e00000;
      24815: inst = 32'hfe0aa19;
      24816: inst = 32'h5be00000;
      24817: inst = 32'h244c8000;
      24818: inst = 32'h24428800;
      24819: inst = 32'h8620000;
      24820: inst = 32'h2a0e0006;
      24821: inst = 32'h294f000a;
      24822: inst = 32'h11200000;
      24823: inst = 32'hd2060fb;
      24824: inst = 32'h13e00000;
      24825: inst = 32'hfe0aa19;
      24826: inst = 32'h5be00000;
      24827: inst = 32'h244c8000;
      24828: inst = 32'h24428800;
      24829: inst = 32'h8620000;
      24830: inst = 32'h2a0e0005;
      24831: inst = 32'h294f000a;
      24832: inst = 32'h11200000;
      24833: inst = 32'hd206105;
      24834: inst = 32'h13e00000;
      24835: inst = 32'hfe0aa19;
      24836: inst = 32'h5be00000;
      24837: inst = 32'h244c8000;
      24838: inst = 32'h24428800;
      24839: inst = 32'h8620000;
      24840: inst = 32'h2a0e0004;
      24841: inst = 32'h294f000a;
      24842: inst = 32'h11200000;
      24843: inst = 32'hd20610f;
      24844: inst = 32'h13e00000;
      24845: inst = 32'hfe0aa19;
      24846: inst = 32'h5be00000;
      24847: inst = 32'h244c8000;
      24848: inst = 32'h24428800;
      24849: inst = 32'h8620000;
      24850: inst = 32'h2a0e0003;
      24851: inst = 32'h294f000a;
      24852: inst = 32'h11200000;
      24853: inst = 32'hd206119;
      24854: inst = 32'h13e00000;
      24855: inst = 32'hfe0aa19;
      24856: inst = 32'h5be00000;
      24857: inst = 32'h244c8000;
      24858: inst = 32'h24428800;
      24859: inst = 32'h8620000;
      24860: inst = 32'h13e00000;
      24861: inst = 32'hfe06123;
      24862: inst = 32'h20200001;
      24863: inst = 32'h5be00000;
      24864: inst = 32'h13e00000;
      24865: inst = 32'hfe06126;
      24866: inst = 32'h5be00000;
      24867: inst = 32'h13e00000;
      24868: inst = 32'hfe06126;
      24869: inst = 32'h5be00000;
      24870: inst = 32'h58000000;
      24871: inst = 32'h10408000;
      24872: inst = 32'hc400002;
      24873: inst = 32'h4420000;
      24874: inst = 32'h10600000;
      24875: inst = 32'hc600010;
      24876: inst = 32'h38421800;
      24877: inst = 32'h4042000f;
      24878: inst = 32'h1c40000f;
      24879: inst = 32'h58000000;
      24880: inst = 32'h58200000;
      24881: inst = 32'hc206b50;
      24882: inst = 32'h10408000;
      24883: inst = 32'hc403fe0;
      24884: inst = 32'h8220000;
      24885: inst = 32'h10408000;
      24886: inst = 32'hc403fe1;
      24887: inst = 32'h8220000;
      24888: inst = 32'h10408000;
      24889: inst = 32'hc403fe2;
      24890: inst = 32'h8220000;
      24891: inst = 32'h10408000;
      24892: inst = 32'hc403ff5;
      24893: inst = 32'h8220000;
      24894: inst = 32'h10408000;
      24895: inst = 32'hc403ff8;
      24896: inst = 32'h8220000;
      24897: inst = 32'h10408000;
      24898: inst = 32'hc403ff9;
      24899: inst = 32'h8220000;
      24900: inst = 32'h10408000;
      24901: inst = 32'hc403ffd;
      24902: inst = 32'h8220000;
      24903: inst = 32'h10408000;
      24904: inst = 32'hc403ffe;
      24905: inst = 32'h8220000;
      24906: inst = 32'h10408000;
      24907: inst = 32'hc403fff;
      24908: inst = 32'h8220000;
      24909: inst = 32'h10408000;
      24910: inst = 32'hc404000;
      24911: inst = 32'h8220000;
      24912: inst = 32'h10408000;
      24913: inst = 32'hc404001;
      24914: inst = 32'h8220000;
      24915: inst = 32'h10408000;
      24916: inst = 32'hc404002;
      24917: inst = 32'h8220000;
      24918: inst = 32'h10408000;
      24919: inst = 32'hc404003;
      24920: inst = 32'h8220000;
      24921: inst = 32'h10408000;
      24922: inst = 32'hc404004;
      24923: inst = 32'h8220000;
      24924: inst = 32'h10408000;
      24925: inst = 32'hc404005;
      24926: inst = 32'h8220000;
      24927: inst = 32'h10408000;
      24928: inst = 32'hc404006;
      24929: inst = 32'h8220000;
      24930: inst = 32'h10408000;
      24931: inst = 32'hc404007;
      24932: inst = 32'h8220000;
      24933: inst = 32'h10408000;
      24934: inst = 32'hc404008;
      24935: inst = 32'h8220000;
      24936: inst = 32'h10408000;
      24937: inst = 32'hc404009;
      24938: inst = 32'h8220000;
      24939: inst = 32'h10408000;
      24940: inst = 32'hc40400a;
      24941: inst = 32'h8220000;
      24942: inst = 32'h10408000;
      24943: inst = 32'hc40400b;
      24944: inst = 32'h8220000;
      24945: inst = 32'h10408000;
      24946: inst = 32'hc40400c;
      24947: inst = 32'h8220000;
      24948: inst = 32'h10408000;
      24949: inst = 32'hc40400d;
      24950: inst = 32'h8220000;
      24951: inst = 32'h10408000;
      24952: inst = 32'hc40400e;
      24953: inst = 32'h8220000;
      24954: inst = 32'h10408000;
      24955: inst = 32'hc40400f;
      24956: inst = 32'h8220000;
      24957: inst = 32'h10408000;
      24958: inst = 32'hc404010;
      24959: inst = 32'h8220000;
      24960: inst = 32'h10408000;
      24961: inst = 32'hc404011;
      24962: inst = 32'h8220000;
      24963: inst = 32'h10408000;
      24964: inst = 32'hc404012;
      24965: inst = 32'h8220000;
      24966: inst = 32'h10408000;
      24967: inst = 32'hc404013;
      24968: inst = 32'h8220000;
      24969: inst = 32'h10408000;
      24970: inst = 32'hc404014;
      24971: inst = 32'h8220000;
      24972: inst = 32'h10408000;
      24973: inst = 32'hc404015;
      24974: inst = 32'h8220000;
      24975: inst = 32'h10408000;
      24976: inst = 32'hc404016;
      24977: inst = 32'h8220000;
      24978: inst = 32'h10408000;
      24979: inst = 32'hc404017;
      24980: inst = 32'h8220000;
      24981: inst = 32'h10408000;
      24982: inst = 32'hc404018;
      24983: inst = 32'h8220000;
      24984: inst = 32'h10408000;
      24985: inst = 32'hc404019;
      24986: inst = 32'h8220000;
      24987: inst = 32'h10408000;
      24988: inst = 32'hc40401a;
      24989: inst = 32'h8220000;
      24990: inst = 32'h10408000;
      24991: inst = 32'hc40401b;
      24992: inst = 32'h8220000;
      24993: inst = 32'h10408000;
      24994: inst = 32'hc40401c;
      24995: inst = 32'h8220000;
      24996: inst = 32'h10408000;
      24997: inst = 32'hc40401d;
      24998: inst = 32'h8220000;
      24999: inst = 32'h10408000;
      25000: inst = 32'hc40401e;
      25001: inst = 32'h8220000;
      25002: inst = 32'h10408000;
      25003: inst = 32'hc40401f;
      25004: inst = 32'h8220000;
      25005: inst = 32'h10408000;
      25006: inst = 32'hc404020;
      25007: inst = 32'h8220000;
      25008: inst = 32'h10408000;
      25009: inst = 32'hc404021;
      25010: inst = 32'h8220000;
      25011: inst = 32'h10408000;
      25012: inst = 32'hc404022;
      25013: inst = 32'h8220000;
      25014: inst = 32'h10408000;
      25015: inst = 32'hc404023;
      25016: inst = 32'h8220000;
      25017: inst = 32'h10408000;
      25018: inst = 32'hc404024;
      25019: inst = 32'h8220000;
      25020: inst = 32'h10408000;
      25021: inst = 32'hc404025;
      25022: inst = 32'h8220000;
      25023: inst = 32'h10408000;
      25024: inst = 32'hc404026;
      25025: inst = 32'h8220000;
      25026: inst = 32'h10408000;
      25027: inst = 32'hc404027;
      25028: inst = 32'h8220000;
      25029: inst = 32'h10408000;
      25030: inst = 32'hc404028;
      25031: inst = 32'h8220000;
      25032: inst = 32'h10408000;
      25033: inst = 32'hc404029;
      25034: inst = 32'h8220000;
      25035: inst = 32'h10408000;
      25036: inst = 32'hc40402a;
      25037: inst = 32'h8220000;
      25038: inst = 32'h10408000;
      25039: inst = 32'hc40402b;
      25040: inst = 32'h8220000;
      25041: inst = 32'h10408000;
      25042: inst = 32'hc40402c;
      25043: inst = 32'h8220000;
      25044: inst = 32'h10408000;
      25045: inst = 32'hc40402d;
      25046: inst = 32'h8220000;
      25047: inst = 32'h10408000;
      25048: inst = 32'hc40402e;
      25049: inst = 32'h8220000;
      25050: inst = 32'h10408000;
      25051: inst = 32'hc40402f;
      25052: inst = 32'h8220000;
      25053: inst = 32'h10408000;
      25054: inst = 32'hc404030;
      25055: inst = 32'h8220000;
      25056: inst = 32'h10408000;
      25057: inst = 32'hc404031;
      25058: inst = 32'h8220000;
      25059: inst = 32'h10408000;
      25060: inst = 32'hc404032;
      25061: inst = 32'h8220000;
      25062: inst = 32'h10408000;
      25063: inst = 32'hc404033;
      25064: inst = 32'h8220000;
      25065: inst = 32'h10408000;
      25066: inst = 32'hc404034;
      25067: inst = 32'h8220000;
      25068: inst = 32'h10408000;
      25069: inst = 32'hc404035;
      25070: inst = 32'h8220000;
      25071: inst = 32'h10408000;
      25072: inst = 32'hc404036;
      25073: inst = 32'h8220000;
      25074: inst = 32'h10408000;
      25075: inst = 32'hc404037;
      25076: inst = 32'h8220000;
      25077: inst = 32'h10408000;
      25078: inst = 32'hc404038;
      25079: inst = 32'h8220000;
      25080: inst = 32'h10408000;
      25081: inst = 32'hc404039;
      25082: inst = 32'h8220000;
      25083: inst = 32'h10408000;
      25084: inst = 32'hc40403a;
      25085: inst = 32'h8220000;
      25086: inst = 32'h10408000;
      25087: inst = 32'hc40403b;
      25088: inst = 32'h8220000;
      25089: inst = 32'h10408000;
      25090: inst = 32'hc40403c;
      25091: inst = 32'h8220000;
      25092: inst = 32'h10408000;
      25093: inst = 32'hc40403d;
      25094: inst = 32'h8220000;
      25095: inst = 32'h10408000;
      25096: inst = 32'hc40403e;
      25097: inst = 32'h8220000;
      25098: inst = 32'h10408000;
      25099: inst = 32'hc40403f;
      25100: inst = 32'h8220000;
      25101: inst = 32'h10408000;
      25102: inst = 32'hc404040;
      25103: inst = 32'h8220000;
      25104: inst = 32'h10408000;
      25105: inst = 32'hc404041;
      25106: inst = 32'h8220000;
      25107: inst = 32'h10408000;
      25108: inst = 32'hc404042;
      25109: inst = 32'h8220000;
      25110: inst = 32'h10408000;
      25111: inst = 32'hc404054;
      25112: inst = 32'h8220000;
      25113: inst = 32'h10408000;
      25114: inst = 32'hc404057;
      25115: inst = 32'h8220000;
      25116: inst = 32'h10408000;
      25117: inst = 32'hc404058;
      25118: inst = 32'h8220000;
      25119: inst = 32'h10408000;
      25120: inst = 32'hc40405c;
      25121: inst = 32'h8220000;
      25122: inst = 32'h10408000;
      25123: inst = 32'hc40405d;
      25124: inst = 32'h8220000;
      25125: inst = 32'h10408000;
      25126: inst = 32'hc40405e;
      25127: inst = 32'h8220000;
      25128: inst = 32'h10408000;
      25129: inst = 32'hc40405f;
      25130: inst = 32'h8220000;
      25131: inst = 32'h10408000;
      25132: inst = 32'hc404060;
      25133: inst = 32'h8220000;
      25134: inst = 32'h10408000;
      25135: inst = 32'hc404061;
      25136: inst = 32'h8220000;
      25137: inst = 32'h10408000;
      25138: inst = 32'hc404062;
      25139: inst = 32'h8220000;
      25140: inst = 32'h10408000;
      25141: inst = 32'hc404063;
      25142: inst = 32'h8220000;
      25143: inst = 32'h10408000;
      25144: inst = 32'hc404064;
      25145: inst = 32'h8220000;
      25146: inst = 32'h10408000;
      25147: inst = 32'hc404065;
      25148: inst = 32'h8220000;
      25149: inst = 32'h10408000;
      25150: inst = 32'hc404066;
      25151: inst = 32'h8220000;
      25152: inst = 32'h10408000;
      25153: inst = 32'hc404067;
      25154: inst = 32'h8220000;
      25155: inst = 32'h10408000;
      25156: inst = 32'hc404068;
      25157: inst = 32'h8220000;
      25158: inst = 32'h10408000;
      25159: inst = 32'hc404069;
      25160: inst = 32'h8220000;
      25161: inst = 32'h10408000;
      25162: inst = 32'hc40406a;
      25163: inst = 32'h8220000;
      25164: inst = 32'h10408000;
      25165: inst = 32'hc40406b;
      25166: inst = 32'h8220000;
      25167: inst = 32'h10408000;
      25168: inst = 32'hc40406c;
      25169: inst = 32'h8220000;
      25170: inst = 32'h10408000;
      25171: inst = 32'hc40406d;
      25172: inst = 32'h8220000;
      25173: inst = 32'h10408000;
      25174: inst = 32'hc40406e;
      25175: inst = 32'h8220000;
      25176: inst = 32'h10408000;
      25177: inst = 32'hc40406f;
      25178: inst = 32'h8220000;
      25179: inst = 32'h10408000;
      25180: inst = 32'hc404070;
      25181: inst = 32'h8220000;
      25182: inst = 32'h10408000;
      25183: inst = 32'hc404071;
      25184: inst = 32'h8220000;
      25185: inst = 32'h10408000;
      25186: inst = 32'hc404072;
      25187: inst = 32'h8220000;
      25188: inst = 32'h10408000;
      25189: inst = 32'hc404073;
      25190: inst = 32'h8220000;
      25191: inst = 32'h10408000;
      25192: inst = 32'hc404074;
      25193: inst = 32'h8220000;
      25194: inst = 32'h10408000;
      25195: inst = 32'hc404075;
      25196: inst = 32'h8220000;
      25197: inst = 32'h10408000;
      25198: inst = 32'hc404076;
      25199: inst = 32'h8220000;
      25200: inst = 32'h10408000;
      25201: inst = 32'hc404077;
      25202: inst = 32'h8220000;
      25203: inst = 32'h10408000;
      25204: inst = 32'hc404078;
      25205: inst = 32'h8220000;
      25206: inst = 32'h10408000;
      25207: inst = 32'hc404079;
      25208: inst = 32'h8220000;
      25209: inst = 32'h10408000;
      25210: inst = 32'hc40407a;
      25211: inst = 32'h8220000;
      25212: inst = 32'h10408000;
      25213: inst = 32'hc40407b;
      25214: inst = 32'h8220000;
      25215: inst = 32'h10408000;
      25216: inst = 32'hc40407c;
      25217: inst = 32'h8220000;
      25218: inst = 32'h10408000;
      25219: inst = 32'hc40407d;
      25220: inst = 32'h8220000;
      25221: inst = 32'h10408000;
      25222: inst = 32'hc40407e;
      25223: inst = 32'h8220000;
      25224: inst = 32'h10408000;
      25225: inst = 32'hc40407f;
      25226: inst = 32'h8220000;
      25227: inst = 32'h10408000;
      25228: inst = 32'hc404080;
      25229: inst = 32'h8220000;
      25230: inst = 32'h10408000;
      25231: inst = 32'hc404081;
      25232: inst = 32'h8220000;
      25233: inst = 32'h10408000;
      25234: inst = 32'hc404082;
      25235: inst = 32'h8220000;
      25236: inst = 32'h10408000;
      25237: inst = 32'hc404083;
      25238: inst = 32'h8220000;
      25239: inst = 32'h10408000;
      25240: inst = 32'hc404084;
      25241: inst = 32'h8220000;
      25242: inst = 32'h10408000;
      25243: inst = 32'hc404085;
      25244: inst = 32'h8220000;
      25245: inst = 32'h10408000;
      25246: inst = 32'hc404086;
      25247: inst = 32'h8220000;
      25248: inst = 32'h10408000;
      25249: inst = 32'hc404087;
      25250: inst = 32'h8220000;
      25251: inst = 32'h10408000;
      25252: inst = 32'hc404088;
      25253: inst = 32'h8220000;
      25254: inst = 32'h10408000;
      25255: inst = 32'hc404089;
      25256: inst = 32'h8220000;
      25257: inst = 32'h10408000;
      25258: inst = 32'hc40408a;
      25259: inst = 32'h8220000;
      25260: inst = 32'h10408000;
      25261: inst = 32'hc40408b;
      25262: inst = 32'h8220000;
      25263: inst = 32'h10408000;
      25264: inst = 32'hc40408c;
      25265: inst = 32'h8220000;
      25266: inst = 32'h10408000;
      25267: inst = 32'hc40408d;
      25268: inst = 32'h8220000;
      25269: inst = 32'h10408000;
      25270: inst = 32'hc40408e;
      25271: inst = 32'h8220000;
      25272: inst = 32'h10408000;
      25273: inst = 32'hc40408f;
      25274: inst = 32'h8220000;
      25275: inst = 32'h10408000;
      25276: inst = 32'hc404090;
      25277: inst = 32'h8220000;
      25278: inst = 32'h10408000;
      25279: inst = 32'hc404091;
      25280: inst = 32'h8220000;
      25281: inst = 32'h10408000;
      25282: inst = 32'hc404092;
      25283: inst = 32'h8220000;
      25284: inst = 32'h10408000;
      25285: inst = 32'hc404093;
      25286: inst = 32'h8220000;
      25287: inst = 32'h10408000;
      25288: inst = 32'hc404094;
      25289: inst = 32'h8220000;
      25290: inst = 32'h10408000;
      25291: inst = 32'hc404095;
      25292: inst = 32'h8220000;
      25293: inst = 32'h10408000;
      25294: inst = 32'hc404096;
      25295: inst = 32'h8220000;
      25296: inst = 32'h10408000;
      25297: inst = 32'hc404097;
      25298: inst = 32'h8220000;
      25299: inst = 32'h10408000;
      25300: inst = 32'hc404098;
      25301: inst = 32'h8220000;
      25302: inst = 32'h10408000;
      25303: inst = 32'hc404099;
      25304: inst = 32'h8220000;
      25305: inst = 32'h10408000;
      25306: inst = 32'hc40409a;
      25307: inst = 32'h8220000;
      25308: inst = 32'h10408000;
      25309: inst = 32'hc40409b;
      25310: inst = 32'h8220000;
      25311: inst = 32'h10408000;
      25312: inst = 32'hc40409c;
      25313: inst = 32'h8220000;
      25314: inst = 32'h10408000;
      25315: inst = 32'hc40409d;
      25316: inst = 32'h8220000;
      25317: inst = 32'h10408000;
      25318: inst = 32'hc40409e;
      25319: inst = 32'h8220000;
      25320: inst = 32'h10408000;
      25321: inst = 32'hc40409f;
      25322: inst = 32'h8220000;
      25323: inst = 32'h10408000;
      25324: inst = 32'hc4040a0;
      25325: inst = 32'h8220000;
      25326: inst = 32'h10408000;
      25327: inst = 32'hc4040a1;
      25328: inst = 32'h8220000;
      25329: inst = 32'h10408000;
      25330: inst = 32'hc4040a2;
      25331: inst = 32'h8220000;
      25332: inst = 32'h10408000;
      25333: inst = 32'hc4040af;
      25334: inst = 32'h8220000;
      25335: inst = 32'h10408000;
      25336: inst = 32'hc4040b2;
      25337: inst = 32'h8220000;
      25338: inst = 32'h10408000;
      25339: inst = 32'hc4040b7;
      25340: inst = 32'h8220000;
      25341: inst = 32'h10408000;
      25342: inst = 32'hc4040b8;
      25343: inst = 32'h8220000;
      25344: inst = 32'h10408000;
      25345: inst = 32'hc4040bb;
      25346: inst = 32'h8220000;
      25347: inst = 32'h10408000;
      25348: inst = 32'hc4040bc;
      25349: inst = 32'h8220000;
      25350: inst = 32'h10408000;
      25351: inst = 32'hc4040bd;
      25352: inst = 32'h8220000;
      25353: inst = 32'h10408000;
      25354: inst = 32'hc4040be;
      25355: inst = 32'h8220000;
      25356: inst = 32'h10408000;
      25357: inst = 32'hc4040bf;
      25358: inst = 32'h8220000;
      25359: inst = 32'h10408000;
      25360: inst = 32'hc4040c0;
      25361: inst = 32'h8220000;
      25362: inst = 32'h10408000;
      25363: inst = 32'hc4040c1;
      25364: inst = 32'h8220000;
      25365: inst = 32'h10408000;
      25366: inst = 32'hc4040c2;
      25367: inst = 32'h8220000;
      25368: inst = 32'h10408000;
      25369: inst = 32'hc4040c3;
      25370: inst = 32'h8220000;
      25371: inst = 32'h10408000;
      25372: inst = 32'hc4040c4;
      25373: inst = 32'h8220000;
      25374: inst = 32'h10408000;
      25375: inst = 32'hc4040c5;
      25376: inst = 32'h8220000;
      25377: inst = 32'h10408000;
      25378: inst = 32'hc4040c6;
      25379: inst = 32'h8220000;
      25380: inst = 32'h10408000;
      25381: inst = 32'hc4040c7;
      25382: inst = 32'h8220000;
      25383: inst = 32'h10408000;
      25384: inst = 32'hc4040c8;
      25385: inst = 32'h8220000;
      25386: inst = 32'h10408000;
      25387: inst = 32'hc4040c9;
      25388: inst = 32'h8220000;
      25389: inst = 32'h10408000;
      25390: inst = 32'hc4040ca;
      25391: inst = 32'h8220000;
      25392: inst = 32'h10408000;
      25393: inst = 32'hc4040cb;
      25394: inst = 32'h8220000;
      25395: inst = 32'h10408000;
      25396: inst = 32'hc4040cc;
      25397: inst = 32'h8220000;
      25398: inst = 32'h10408000;
      25399: inst = 32'hc4040cd;
      25400: inst = 32'h8220000;
      25401: inst = 32'h10408000;
      25402: inst = 32'hc4040ce;
      25403: inst = 32'h8220000;
      25404: inst = 32'h10408000;
      25405: inst = 32'hc4040cf;
      25406: inst = 32'h8220000;
      25407: inst = 32'h10408000;
      25408: inst = 32'hc4040d0;
      25409: inst = 32'h8220000;
      25410: inst = 32'h10408000;
      25411: inst = 32'hc4040d1;
      25412: inst = 32'h8220000;
      25413: inst = 32'h10408000;
      25414: inst = 32'hc4040d2;
      25415: inst = 32'h8220000;
      25416: inst = 32'h10408000;
      25417: inst = 32'hc4040d3;
      25418: inst = 32'h8220000;
      25419: inst = 32'h10408000;
      25420: inst = 32'hc4040d4;
      25421: inst = 32'h8220000;
      25422: inst = 32'h10408000;
      25423: inst = 32'hc4040d5;
      25424: inst = 32'h8220000;
      25425: inst = 32'h10408000;
      25426: inst = 32'hc4040d6;
      25427: inst = 32'h8220000;
      25428: inst = 32'h10408000;
      25429: inst = 32'hc4040d7;
      25430: inst = 32'h8220000;
      25431: inst = 32'h10408000;
      25432: inst = 32'hc4040d8;
      25433: inst = 32'h8220000;
      25434: inst = 32'h10408000;
      25435: inst = 32'hc4040d9;
      25436: inst = 32'h8220000;
      25437: inst = 32'h10408000;
      25438: inst = 32'hc4040da;
      25439: inst = 32'h8220000;
      25440: inst = 32'h10408000;
      25441: inst = 32'hc4040db;
      25442: inst = 32'h8220000;
      25443: inst = 32'h10408000;
      25444: inst = 32'hc4040dc;
      25445: inst = 32'h8220000;
      25446: inst = 32'h10408000;
      25447: inst = 32'hc4040dd;
      25448: inst = 32'h8220000;
      25449: inst = 32'h10408000;
      25450: inst = 32'hc4040de;
      25451: inst = 32'h8220000;
      25452: inst = 32'h10408000;
      25453: inst = 32'hc4040df;
      25454: inst = 32'h8220000;
      25455: inst = 32'h10408000;
      25456: inst = 32'hc4040e0;
      25457: inst = 32'h8220000;
      25458: inst = 32'h10408000;
      25459: inst = 32'hc4040e1;
      25460: inst = 32'h8220000;
      25461: inst = 32'h10408000;
      25462: inst = 32'hc4040e2;
      25463: inst = 32'h8220000;
      25464: inst = 32'h10408000;
      25465: inst = 32'hc4040e3;
      25466: inst = 32'h8220000;
      25467: inst = 32'h10408000;
      25468: inst = 32'hc4040e4;
      25469: inst = 32'h8220000;
      25470: inst = 32'h10408000;
      25471: inst = 32'hc4040e5;
      25472: inst = 32'h8220000;
      25473: inst = 32'h10408000;
      25474: inst = 32'hc4040e6;
      25475: inst = 32'h8220000;
      25476: inst = 32'h10408000;
      25477: inst = 32'hc4040e7;
      25478: inst = 32'h8220000;
      25479: inst = 32'h10408000;
      25480: inst = 32'hc4040e8;
      25481: inst = 32'h8220000;
      25482: inst = 32'h10408000;
      25483: inst = 32'hc4040e9;
      25484: inst = 32'h8220000;
      25485: inst = 32'h10408000;
      25486: inst = 32'hc4040ea;
      25487: inst = 32'h8220000;
      25488: inst = 32'h10408000;
      25489: inst = 32'hc4040eb;
      25490: inst = 32'h8220000;
      25491: inst = 32'h10408000;
      25492: inst = 32'hc4040ec;
      25493: inst = 32'h8220000;
      25494: inst = 32'h10408000;
      25495: inst = 32'hc4040ed;
      25496: inst = 32'h8220000;
      25497: inst = 32'h10408000;
      25498: inst = 32'hc4040ee;
      25499: inst = 32'h8220000;
      25500: inst = 32'h10408000;
      25501: inst = 32'hc4040ef;
      25502: inst = 32'h8220000;
      25503: inst = 32'h10408000;
      25504: inst = 32'hc4040f0;
      25505: inst = 32'h8220000;
      25506: inst = 32'h10408000;
      25507: inst = 32'hc4040f1;
      25508: inst = 32'h8220000;
      25509: inst = 32'h10408000;
      25510: inst = 32'hc4040f2;
      25511: inst = 32'h8220000;
      25512: inst = 32'h10408000;
      25513: inst = 32'hc4040f3;
      25514: inst = 32'h8220000;
      25515: inst = 32'h10408000;
      25516: inst = 32'hc4040f4;
      25517: inst = 32'h8220000;
      25518: inst = 32'h10408000;
      25519: inst = 32'hc4040f5;
      25520: inst = 32'h8220000;
      25521: inst = 32'h10408000;
      25522: inst = 32'hc4040f6;
      25523: inst = 32'h8220000;
      25524: inst = 32'h10408000;
      25525: inst = 32'hc4040f7;
      25526: inst = 32'h8220000;
      25527: inst = 32'h10408000;
      25528: inst = 32'hc4040f8;
      25529: inst = 32'h8220000;
      25530: inst = 32'h10408000;
      25531: inst = 32'hc4040f9;
      25532: inst = 32'h8220000;
      25533: inst = 32'h10408000;
      25534: inst = 32'hc4040fa;
      25535: inst = 32'h8220000;
      25536: inst = 32'h10408000;
      25537: inst = 32'hc4040fb;
      25538: inst = 32'h8220000;
      25539: inst = 32'h10408000;
      25540: inst = 32'hc4040fc;
      25541: inst = 32'h8220000;
      25542: inst = 32'h10408000;
      25543: inst = 32'hc4040fd;
      25544: inst = 32'h8220000;
      25545: inst = 32'h10408000;
      25546: inst = 32'hc4040fe;
      25547: inst = 32'h8220000;
      25548: inst = 32'h10408000;
      25549: inst = 32'hc4040ff;
      25550: inst = 32'h8220000;
      25551: inst = 32'h10408000;
      25552: inst = 32'hc404100;
      25553: inst = 32'h8220000;
      25554: inst = 32'h10408000;
      25555: inst = 32'hc404101;
      25556: inst = 32'h8220000;
      25557: inst = 32'h10408000;
      25558: inst = 32'hc404102;
      25559: inst = 32'h8220000;
      25560: inst = 32'h10408000;
      25561: inst = 32'hc40414c;
      25562: inst = 32'h8220000;
      25563: inst = 32'h10408000;
      25564: inst = 32'hc40414d;
      25565: inst = 32'h8220000;
      25566: inst = 32'h10408000;
      25567: inst = 32'hc40414e;
      25568: inst = 32'h8220000;
      25569: inst = 32'h10408000;
      25570: inst = 32'hc40415d;
      25571: inst = 32'h8220000;
      25572: inst = 32'h10408000;
      25573: inst = 32'hc40415e;
      25574: inst = 32'h8220000;
      25575: inst = 32'h10408000;
      25576: inst = 32'hc40415f;
      25577: inst = 32'h8220000;
      25578: inst = 32'h10408000;
      25579: inst = 32'hc404160;
      25580: inst = 32'h8220000;
      25581: inst = 32'h10408000;
      25582: inst = 32'hc404161;
      25583: inst = 32'h8220000;
      25584: inst = 32'h10408000;
      25585: inst = 32'hc404162;
      25586: inst = 32'h8220000;
      25587: inst = 32'h10408000;
      25588: inst = 32'hc4041ac;
      25589: inst = 32'h8220000;
      25590: inst = 32'h10408000;
      25591: inst = 32'hc4041ad;
      25592: inst = 32'h8220000;
      25593: inst = 32'h10408000;
      25594: inst = 32'hc4041ae;
      25595: inst = 32'h8220000;
      25596: inst = 32'h10408000;
      25597: inst = 32'hc4041bd;
      25598: inst = 32'h8220000;
      25599: inst = 32'h10408000;
      25600: inst = 32'hc4041be;
      25601: inst = 32'h8220000;
      25602: inst = 32'h10408000;
      25603: inst = 32'hc4041bf;
      25604: inst = 32'h8220000;
      25605: inst = 32'h10408000;
      25606: inst = 32'hc4041c0;
      25607: inst = 32'h8220000;
      25608: inst = 32'h10408000;
      25609: inst = 32'hc4041c1;
      25610: inst = 32'h8220000;
      25611: inst = 32'h10408000;
      25612: inst = 32'hc4041c2;
      25613: inst = 32'h8220000;
      25614: inst = 32'h10408000;
      25615: inst = 32'hc40420c;
      25616: inst = 32'h8220000;
      25617: inst = 32'h10408000;
      25618: inst = 32'hc40420d;
      25619: inst = 32'h8220000;
      25620: inst = 32'h10408000;
      25621: inst = 32'hc40420e;
      25622: inst = 32'h8220000;
      25623: inst = 32'h10408000;
      25624: inst = 32'hc40421d;
      25625: inst = 32'h8220000;
      25626: inst = 32'h10408000;
      25627: inst = 32'hc40421e;
      25628: inst = 32'h8220000;
      25629: inst = 32'h10408000;
      25630: inst = 32'hc40421f;
      25631: inst = 32'h8220000;
      25632: inst = 32'h10408000;
      25633: inst = 32'hc404220;
      25634: inst = 32'h8220000;
      25635: inst = 32'h10408000;
      25636: inst = 32'hc404221;
      25637: inst = 32'h8220000;
      25638: inst = 32'h10408000;
      25639: inst = 32'hc404222;
      25640: inst = 32'h8220000;
      25641: inst = 32'h10408000;
      25642: inst = 32'hc40426c;
      25643: inst = 32'h8220000;
      25644: inst = 32'h10408000;
      25645: inst = 32'hc40426d;
      25646: inst = 32'h8220000;
      25647: inst = 32'h10408000;
      25648: inst = 32'hc40426e;
      25649: inst = 32'h8220000;
      25650: inst = 32'h10408000;
      25651: inst = 32'hc40427d;
      25652: inst = 32'h8220000;
      25653: inst = 32'h10408000;
      25654: inst = 32'hc40427e;
      25655: inst = 32'h8220000;
      25656: inst = 32'h10408000;
      25657: inst = 32'hc40427f;
      25658: inst = 32'h8220000;
      25659: inst = 32'h10408000;
      25660: inst = 32'hc404280;
      25661: inst = 32'h8220000;
      25662: inst = 32'h10408000;
      25663: inst = 32'hc404281;
      25664: inst = 32'h8220000;
      25665: inst = 32'h10408000;
      25666: inst = 32'hc404282;
      25667: inst = 32'h8220000;
      25668: inst = 32'h10408000;
      25669: inst = 32'hc4042cc;
      25670: inst = 32'h8220000;
      25671: inst = 32'h10408000;
      25672: inst = 32'hc4042cd;
      25673: inst = 32'h8220000;
      25674: inst = 32'h10408000;
      25675: inst = 32'hc4042ce;
      25676: inst = 32'h8220000;
      25677: inst = 32'h10408000;
      25678: inst = 32'hc4042dd;
      25679: inst = 32'h8220000;
      25680: inst = 32'h10408000;
      25681: inst = 32'hc4042de;
      25682: inst = 32'h8220000;
      25683: inst = 32'h10408000;
      25684: inst = 32'hc4042df;
      25685: inst = 32'h8220000;
      25686: inst = 32'h10408000;
      25687: inst = 32'hc4042e0;
      25688: inst = 32'h8220000;
      25689: inst = 32'h10408000;
      25690: inst = 32'hc4042e1;
      25691: inst = 32'h8220000;
      25692: inst = 32'h10408000;
      25693: inst = 32'hc4042e2;
      25694: inst = 32'h8220000;
      25695: inst = 32'h10408000;
      25696: inst = 32'hc40432c;
      25697: inst = 32'h8220000;
      25698: inst = 32'h10408000;
      25699: inst = 32'hc40432d;
      25700: inst = 32'h8220000;
      25701: inst = 32'h10408000;
      25702: inst = 32'hc40432e;
      25703: inst = 32'h8220000;
      25704: inst = 32'h10408000;
      25705: inst = 32'hc40433d;
      25706: inst = 32'h8220000;
      25707: inst = 32'h10408000;
      25708: inst = 32'hc40433e;
      25709: inst = 32'h8220000;
      25710: inst = 32'h10408000;
      25711: inst = 32'hc40433f;
      25712: inst = 32'h8220000;
      25713: inst = 32'h10408000;
      25714: inst = 32'hc404340;
      25715: inst = 32'h8220000;
      25716: inst = 32'h10408000;
      25717: inst = 32'hc404341;
      25718: inst = 32'h8220000;
      25719: inst = 32'h10408000;
      25720: inst = 32'hc404342;
      25721: inst = 32'h8220000;
      25722: inst = 32'h10408000;
      25723: inst = 32'hc40438c;
      25724: inst = 32'h8220000;
      25725: inst = 32'h10408000;
      25726: inst = 32'hc40438d;
      25727: inst = 32'h8220000;
      25728: inst = 32'h10408000;
      25729: inst = 32'hc40438e;
      25730: inst = 32'h8220000;
      25731: inst = 32'h10408000;
      25732: inst = 32'hc40439d;
      25733: inst = 32'h8220000;
      25734: inst = 32'h10408000;
      25735: inst = 32'hc40439e;
      25736: inst = 32'h8220000;
      25737: inst = 32'h10408000;
      25738: inst = 32'hc40439f;
      25739: inst = 32'h8220000;
      25740: inst = 32'h10408000;
      25741: inst = 32'hc4043a0;
      25742: inst = 32'h8220000;
      25743: inst = 32'h10408000;
      25744: inst = 32'hc4043a1;
      25745: inst = 32'h8220000;
      25746: inst = 32'h10408000;
      25747: inst = 32'hc4043a2;
      25748: inst = 32'h8220000;
      25749: inst = 32'h10408000;
      25750: inst = 32'hc4043ec;
      25751: inst = 32'h8220000;
      25752: inst = 32'h10408000;
      25753: inst = 32'hc4043ed;
      25754: inst = 32'h8220000;
      25755: inst = 32'h10408000;
      25756: inst = 32'hc4043ee;
      25757: inst = 32'h8220000;
      25758: inst = 32'h10408000;
      25759: inst = 32'hc4043fd;
      25760: inst = 32'h8220000;
      25761: inst = 32'h10408000;
      25762: inst = 32'hc4043fe;
      25763: inst = 32'h8220000;
      25764: inst = 32'h10408000;
      25765: inst = 32'hc4043ff;
      25766: inst = 32'h8220000;
      25767: inst = 32'h10408000;
      25768: inst = 32'hc404400;
      25769: inst = 32'h8220000;
      25770: inst = 32'h10408000;
      25771: inst = 32'hc404401;
      25772: inst = 32'h8220000;
      25773: inst = 32'h10408000;
      25774: inst = 32'hc404402;
      25775: inst = 32'h8220000;
      25776: inst = 32'h10408000;
      25777: inst = 32'hc40444c;
      25778: inst = 32'h8220000;
      25779: inst = 32'h10408000;
      25780: inst = 32'hc40444d;
      25781: inst = 32'h8220000;
      25782: inst = 32'h10408000;
      25783: inst = 32'hc40444e;
      25784: inst = 32'h8220000;
      25785: inst = 32'h10408000;
      25786: inst = 32'hc40445d;
      25787: inst = 32'h8220000;
      25788: inst = 32'h10408000;
      25789: inst = 32'hc40445e;
      25790: inst = 32'h8220000;
      25791: inst = 32'h10408000;
      25792: inst = 32'hc40445f;
      25793: inst = 32'h8220000;
      25794: inst = 32'h10408000;
      25795: inst = 32'hc404460;
      25796: inst = 32'h8220000;
      25797: inst = 32'h10408000;
      25798: inst = 32'hc404461;
      25799: inst = 32'h8220000;
      25800: inst = 32'h10408000;
      25801: inst = 32'hc404462;
      25802: inst = 32'h8220000;
      25803: inst = 32'h10408000;
      25804: inst = 32'hc4044ac;
      25805: inst = 32'h8220000;
      25806: inst = 32'h10408000;
      25807: inst = 32'hc4044ad;
      25808: inst = 32'h8220000;
      25809: inst = 32'h10408000;
      25810: inst = 32'hc4044ae;
      25811: inst = 32'h8220000;
      25812: inst = 32'h10408000;
      25813: inst = 32'hc4044bd;
      25814: inst = 32'h8220000;
      25815: inst = 32'h10408000;
      25816: inst = 32'hc4044be;
      25817: inst = 32'h8220000;
      25818: inst = 32'h10408000;
      25819: inst = 32'hc4044bf;
      25820: inst = 32'h8220000;
      25821: inst = 32'h10408000;
      25822: inst = 32'hc4044c0;
      25823: inst = 32'h8220000;
      25824: inst = 32'h10408000;
      25825: inst = 32'hc4044c1;
      25826: inst = 32'h8220000;
      25827: inst = 32'h10408000;
      25828: inst = 32'hc4044c2;
      25829: inst = 32'h8220000;
      25830: inst = 32'h10408000;
      25831: inst = 32'hc40450c;
      25832: inst = 32'h8220000;
      25833: inst = 32'h10408000;
      25834: inst = 32'hc40450d;
      25835: inst = 32'h8220000;
      25836: inst = 32'h10408000;
      25837: inst = 32'hc40450e;
      25838: inst = 32'h8220000;
      25839: inst = 32'h10408000;
      25840: inst = 32'hc40451d;
      25841: inst = 32'h8220000;
      25842: inst = 32'h10408000;
      25843: inst = 32'hc40451e;
      25844: inst = 32'h8220000;
      25845: inst = 32'h10408000;
      25846: inst = 32'hc40451f;
      25847: inst = 32'h8220000;
      25848: inst = 32'h10408000;
      25849: inst = 32'hc404520;
      25850: inst = 32'h8220000;
      25851: inst = 32'h10408000;
      25852: inst = 32'hc404521;
      25853: inst = 32'h8220000;
      25854: inst = 32'h10408000;
      25855: inst = 32'hc404522;
      25856: inst = 32'h8220000;
      25857: inst = 32'h10408000;
      25858: inst = 32'hc40456c;
      25859: inst = 32'h8220000;
      25860: inst = 32'h10408000;
      25861: inst = 32'hc40456d;
      25862: inst = 32'h8220000;
      25863: inst = 32'h10408000;
      25864: inst = 32'hc40456e;
      25865: inst = 32'h8220000;
      25866: inst = 32'h10408000;
      25867: inst = 32'hc40457d;
      25868: inst = 32'h8220000;
      25869: inst = 32'h10408000;
      25870: inst = 32'hc40457e;
      25871: inst = 32'h8220000;
      25872: inst = 32'h10408000;
      25873: inst = 32'hc40457f;
      25874: inst = 32'h8220000;
      25875: inst = 32'h10408000;
      25876: inst = 32'hc404580;
      25877: inst = 32'h8220000;
      25878: inst = 32'h10408000;
      25879: inst = 32'hc404581;
      25880: inst = 32'h8220000;
      25881: inst = 32'h10408000;
      25882: inst = 32'hc404582;
      25883: inst = 32'h8220000;
      25884: inst = 32'h10408000;
      25885: inst = 32'hc4045cc;
      25886: inst = 32'h8220000;
      25887: inst = 32'h10408000;
      25888: inst = 32'hc4045cd;
      25889: inst = 32'h8220000;
      25890: inst = 32'h10408000;
      25891: inst = 32'hc4045ce;
      25892: inst = 32'h8220000;
      25893: inst = 32'h10408000;
      25894: inst = 32'hc4045dd;
      25895: inst = 32'h8220000;
      25896: inst = 32'h10408000;
      25897: inst = 32'hc4045de;
      25898: inst = 32'h8220000;
      25899: inst = 32'h10408000;
      25900: inst = 32'hc4045df;
      25901: inst = 32'h8220000;
      25902: inst = 32'h10408000;
      25903: inst = 32'hc4045e0;
      25904: inst = 32'h8220000;
      25905: inst = 32'h10408000;
      25906: inst = 32'hc4045e1;
      25907: inst = 32'h8220000;
      25908: inst = 32'h10408000;
      25909: inst = 32'hc4045e2;
      25910: inst = 32'h8220000;
      25911: inst = 32'h10408000;
      25912: inst = 32'hc40462c;
      25913: inst = 32'h8220000;
      25914: inst = 32'h10408000;
      25915: inst = 32'hc40462d;
      25916: inst = 32'h8220000;
      25917: inst = 32'h10408000;
      25918: inst = 32'hc40462e;
      25919: inst = 32'h8220000;
      25920: inst = 32'h10408000;
      25921: inst = 32'hc40463d;
      25922: inst = 32'h8220000;
      25923: inst = 32'h10408000;
      25924: inst = 32'hc40463e;
      25925: inst = 32'h8220000;
      25926: inst = 32'h10408000;
      25927: inst = 32'hc40463f;
      25928: inst = 32'h8220000;
      25929: inst = 32'h10408000;
      25930: inst = 32'hc404640;
      25931: inst = 32'h8220000;
      25932: inst = 32'h10408000;
      25933: inst = 32'hc404641;
      25934: inst = 32'h8220000;
      25935: inst = 32'h10408000;
      25936: inst = 32'hc404642;
      25937: inst = 32'h8220000;
      25938: inst = 32'h10408000;
      25939: inst = 32'hc40464e;
      25940: inst = 32'h8220000;
      25941: inst = 32'h10408000;
      25942: inst = 32'hc40464f;
      25943: inst = 32'h8220000;
      25944: inst = 32'h10408000;
      25945: inst = 32'hc404650;
      25946: inst = 32'h8220000;
      25947: inst = 32'h10408000;
      25948: inst = 32'hc404651;
      25949: inst = 32'h8220000;
      25950: inst = 32'h10408000;
      25951: inst = 32'hc404652;
      25952: inst = 32'h8220000;
      25953: inst = 32'h10408000;
      25954: inst = 32'hc404653;
      25955: inst = 32'h8220000;
      25956: inst = 32'h10408000;
      25957: inst = 32'hc404654;
      25958: inst = 32'h8220000;
      25959: inst = 32'h10408000;
      25960: inst = 32'hc404655;
      25961: inst = 32'h8220000;
      25962: inst = 32'h10408000;
      25963: inst = 32'hc404656;
      25964: inst = 32'h8220000;
      25965: inst = 32'h10408000;
      25966: inst = 32'hc404657;
      25967: inst = 32'h8220000;
      25968: inst = 32'h10408000;
      25969: inst = 32'hc404658;
      25970: inst = 32'h8220000;
      25971: inst = 32'h10408000;
      25972: inst = 32'hc404659;
      25973: inst = 32'h8220000;
      25974: inst = 32'h10408000;
      25975: inst = 32'hc40465a;
      25976: inst = 32'h8220000;
      25977: inst = 32'h10408000;
      25978: inst = 32'hc40465b;
      25979: inst = 32'h8220000;
      25980: inst = 32'h10408000;
      25981: inst = 32'hc40465c;
      25982: inst = 32'h8220000;
      25983: inst = 32'h10408000;
      25984: inst = 32'hc40465d;
      25985: inst = 32'h8220000;
      25986: inst = 32'h10408000;
      25987: inst = 32'hc40465e;
      25988: inst = 32'h8220000;
      25989: inst = 32'h10408000;
      25990: inst = 32'hc40465f;
      25991: inst = 32'h8220000;
      25992: inst = 32'h10408000;
      25993: inst = 32'hc404660;
      25994: inst = 32'h8220000;
      25995: inst = 32'h10408000;
      25996: inst = 32'hc404661;
      25997: inst = 32'h8220000;
      25998: inst = 32'h10408000;
      25999: inst = 32'hc404662;
      26000: inst = 32'h8220000;
      26001: inst = 32'h10408000;
      26002: inst = 32'hc404663;
      26003: inst = 32'h8220000;
      26004: inst = 32'h10408000;
      26005: inst = 32'hc404664;
      26006: inst = 32'h8220000;
      26007: inst = 32'h10408000;
      26008: inst = 32'hc404665;
      26009: inst = 32'h8220000;
      26010: inst = 32'h10408000;
      26011: inst = 32'hc404666;
      26012: inst = 32'h8220000;
      26013: inst = 32'h10408000;
      26014: inst = 32'hc404667;
      26015: inst = 32'h8220000;
      26016: inst = 32'h10408000;
      26017: inst = 32'hc404668;
      26018: inst = 32'h8220000;
      26019: inst = 32'h10408000;
      26020: inst = 32'hc404669;
      26021: inst = 32'h8220000;
      26022: inst = 32'h10408000;
      26023: inst = 32'hc40466e;
      26024: inst = 32'h8220000;
      26025: inst = 32'h10408000;
      26026: inst = 32'hc40466f;
      26027: inst = 32'h8220000;
      26028: inst = 32'h10408000;
      26029: inst = 32'hc404673;
      26030: inst = 32'h8220000;
      26031: inst = 32'h10408000;
      26032: inst = 32'hc404676;
      26033: inst = 32'h8220000;
      26034: inst = 32'h10408000;
      26035: inst = 32'hc40468c;
      26036: inst = 32'h8220000;
      26037: inst = 32'h10408000;
      26038: inst = 32'hc40468d;
      26039: inst = 32'h8220000;
      26040: inst = 32'h10408000;
      26041: inst = 32'hc40468e;
      26042: inst = 32'h8220000;
      26043: inst = 32'h10408000;
      26044: inst = 32'hc40469d;
      26045: inst = 32'h8220000;
      26046: inst = 32'h10408000;
      26047: inst = 32'hc40469e;
      26048: inst = 32'h8220000;
      26049: inst = 32'h10408000;
      26050: inst = 32'hc40469f;
      26051: inst = 32'h8220000;
      26052: inst = 32'h10408000;
      26053: inst = 32'hc4046a0;
      26054: inst = 32'h8220000;
      26055: inst = 32'h10408000;
      26056: inst = 32'hc4046a1;
      26057: inst = 32'h8220000;
      26058: inst = 32'h10408000;
      26059: inst = 32'hc4046a2;
      26060: inst = 32'h8220000;
      26061: inst = 32'h10408000;
      26062: inst = 32'hc4046ae;
      26063: inst = 32'h8220000;
      26064: inst = 32'h10408000;
      26065: inst = 32'hc4046af;
      26066: inst = 32'h8220000;
      26067: inst = 32'h10408000;
      26068: inst = 32'hc4046b0;
      26069: inst = 32'h8220000;
      26070: inst = 32'h10408000;
      26071: inst = 32'hc4046b1;
      26072: inst = 32'h8220000;
      26073: inst = 32'h10408000;
      26074: inst = 32'hc4046b2;
      26075: inst = 32'h8220000;
      26076: inst = 32'h10408000;
      26077: inst = 32'hc4046b3;
      26078: inst = 32'h8220000;
      26079: inst = 32'h10408000;
      26080: inst = 32'hc4046b4;
      26081: inst = 32'h8220000;
      26082: inst = 32'h10408000;
      26083: inst = 32'hc4046b5;
      26084: inst = 32'h8220000;
      26085: inst = 32'h10408000;
      26086: inst = 32'hc4046b6;
      26087: inst = 32'h8220000;
      26088: inst = 32'h10408000;
      26089: inst = 32'hc4046b7;
      26090: inst = 32'h8220000;
      26091: inst = 32'h10408000;
      26092: inst = 32'hc4046b8;
      26093: inst = 32'h8220000;
      26094: inst = 32'h10408000;
      26095: inst = 32'hc4046b9;
      26096: inst = 32'h8220000;
      26097: inst = 32'h10408000;
      26098: inst = 32'hc4046ba;
      26099: inst = 32'h8220000;
      26100: inst = 32'h10408000;
      26101: inst = 32'hc4046bb;
      26102: inst = 32'h8220000;
      26103: inst = 32'h10408000;
      26104: inst = 32'hc4046bc;
      26105: inst = 32'h8220000;
      26106: inst = 32'h10408000;
      26107: inst = 32'hc4046bd;
      26108: inst = 32'h8220000;
      26109: inst = 32'h10408000;
      26110: inst = 32'hc4046be;
      26111: inst = 32'h8220000;
      26112: inst = 32'h10408000;
      26113: inst = 32'hc4046bf;
      26114: inst = 32'h8220000;
      26115: inst = 32'h10408000;
      26116: inst = 32'hc4046c0;
      26117: inst = 32'h8220000;
      26118: inst = 32'h10408000;
      26119: inst = 32'hc4046c1;
      26120: inst = 32'h8220000;
      26121: inst = 32'h10408000;
      26122: inst = 32'hc4046c2;
      26123: inst = 32'h8220000;
      26124: inst = 32'h10408000;
      26125: inst = 32'hc4046c3;
      26126: inst = 32'h8220000;
      26127: inst = 32'h10408000;
      26128: inst = 32'hc4046c4;
      26129: inst = 32'h8220000;
      26130: inst = 32'h10408000;
      26131: inst = 32'hc4046c5;
      26132: inst = 32'h8220000;
      26133: inst = 32'h10408000;
      26134: inst = 32'hc4046c6;
      26135: inst = 32'h8220000;
      26136: inst = 32'h10408000;
      26137: inst = 32'hc4046c7;
      26138: inst = 32'h8220000;
      26139: inst = 32'h10408000;
      26140: inst = 32'hc4046c8;
      26141: inst = 32'h8220000;
      26142: inst = 32'h10408000;
      26143: inst = 32'hc4046c9;
      26144: inst = 32'h8220000;
      26145: inst = 32'h10408000;
      26146: inst = 32'hc4046ce;
      26147: inst = 32'h8220000;
      26148: inst = 32'h10408000;
      26149: inst = 32'hc4046cf;
      26150: inst = 32'h8220000;
      26151: inst = 32'h10408000;
      26152: inst = 32'hc4046d0;
      26153: inst = 32'h8220000;
      26154: inst = 32'h10408000;
      26155: inst = 32'hc4046d1;
      26156: inst = 32'h8220000;
      26157: inst = 32'h10408000;
      26158: inst = 32'hc4046d6;
      26159: inst = 32'h8220000;
      26160: inst = 32'h10408000;
      26161: inst = 32'hc4046ec;
      26162: inst = 32'h8220000;
      26163: inst = 32'h10408000;
      26164: inst = 32'hc4046ed;
      26165: inst = 32'h8220000;
      26166: inst = 32'h10408000;
      26167: inst = 32'hc4046ee;
      26168: inst = 32'h8220000;
      26169: inst = 32'h10408000;
      26170: inst = 32'hc4046fd;
      26171: inst = 32'h8220000;
      26172: inst = 32'h10408000;
      26173: inst = 32'hc4046fe;
      26174: inst = 32'h8220000;
      26175: inst = 32'h10408000;
      26176: inst = 32'hc4046ff;
      26177: inst = 32'h8220000;
      26178: inst = 32'h10408000;
      26179: inst = 32'hc404700;
      26180: inst = 32'h8220000;
      26181: inst = 32'h10408000;
      26182: inst = 32'hc404701;
      26183: inst = 32'h8220000;
      26184: inst = 32'h10408000;
      26185: inst = 32'hc404702;
      26186: inst = 32'h8220000;
      26187: inst = 32'h10408000;
      26188: inst = 32'hc40470e;
      26189: inst = 32'h8220000;
      26190: inst = 32'h10408000;
      26191: inst = 32'hc40470f;
      26192: inst = 32'h8220000;
      26193: inst = 32'h10408000;
      26194: inst = 32'hc404710;
      26195: inst = 32'h8220000;
      26196: inst = 32'h10408000;
      26197: inst = 32'hc404711;
      26198: inst = 32'h8220000;
      26199: inst = 32'h10408000;
      26200: inst = 32'hc404712;
      26201: inst = 32'h8220000;
      26202: inst = 32'h10408000;
      26203: inst = 32'hc404713;
      26204: inst = 32'h8220000;
      26205: inst = 32'h10408000;
      26206: inst = 32'hc404714;
      26207: inst = 32'h8220000;
      26208: inst = 32'h10408000;
      26209: inst = 32'hc404715;
      26210: inst = 32'h8220000;
      26211: inst = 32'h10408000;
      26212: inst = 32'hc404716;
      26213: inst = 32'h8220000;
      26214: inst = 32'h10408000;
      26215: inst = 32'hc404717;
      26216: inst = 32'h8220000;
      26217: inst = 32'h10408000;
      26218: inst = 32'hc404718;
      26219: inst = 32'h8220000;
      26220: inst = 32'h10408000;
      26221: inst = 32'hc404719;
      26222: inst = 32'h8220000;
      26223: inst = 32'h10408000;
      26224: inst = 32'hc40471a;
      26225: inst = 32'h8220000;
      26226: inst = 32'h10408000;
      26227: inst = 32'hc40471b;
      26228: inst = 32'h8220000;
      26229: inst = 32'h10408000;
      26230: inst = 32'hc40471c;
      26231: inst = 32'h8220000;
      26232: inst = 32'h10408000;
      26233: inst = 32'hc40471d;
      26234: inst = 32'h8220000;
      26235: inst = 32'h10408000;
      26236: inst = 32'hc40471e;
      26237: inst = 32'h8220000;
      26238: inst = 32'h10408000;
      26239: inst = 32'hc40471f;
      26240: inst = 32'h8220000;
      26241: inst = 32'h10408000;
      26242: inst = 32'hc404720;
      26243: inst = 32'h8220000;
      26244: inst = 32'h10408000;
      26245: inst = 32'hc404721;
      26246: inst = 32'h8220000;
      26247: inst = 32'h10408000;
      26248: inst = 32'hc404722;
      26249: inst = 32'h8220000;
      26250: inst = 32'h10408000;
      26251: inst = 32'hc404723;
      26252: inst = 32'h8220000;
      26253: inst = 32'h10408000;
      26254: inst = 32'hc404724;
      26255: inst = 32'h8220000;
      26256: inst = 32'h10408000;
      26257: inst = 32'hc404725;
      26258: inst = 32'h8220000;
      26259: inst = 32'h10408000;
      26260: inst = 32'hc404726;
      26261: inst = 32'h8220000;
      26262: inst = 32'h10408000;
      26263: inst = 32'hc404727;
      26264: inst = 32'h8220000;
      26265: inst = 32'h10408000;
      26266: inst = 32'hc404728;
      26267: inst = 32'h8220000;
      26268: inst = 32'h10408000;
      26269: inst = 32'hc404729;
      26270: inst = 32'h8220000;
      26271: inst = 32'h10408000;
      26272: inst = 32'hc40472a;
      26273: inst = 32'h8220000;
      26274: inst = 32'h10408000;
      26275: inst = 32'hc40472f;
      26276: inst = 32'h8220000;
      26277: inst = 32'h10408000;
      26278: inst = 32'hc404736;
      26279: inst = 32'h8220000;
      26280: inst = 32'h10408000;
      26281: inst = 32'hc404737;
      26282: inst = 32'h8220000;
      26283: inst = 32'h10408000;
      26284: inst = 32'hc404738;
      26285: inst = 32'h8220000;
      26286: inst = 32'h10408000;
      26287: inst = 32'hc40474c;
      26288: inst = 32'h8220000;
      26289: inst = 32'h10408000;
      26290: inst = 32'hc40474d;
      26291: inst = 32'h8220000;
      26292: inst = 32'h10408000;
      26293: inst = 32'hc40474e;
      26294: inst = 32'h8220000;
      26295: inst = 32'h10408000;
      26296: inst = 32'hc40475d;
      26297: inst = 32'h8220000;
      26298: inst = 32'h10408000;
      26299: inst = 32'hc40475e;
      26300: inst = 32'h8220000;
      26301: inst = 32'h10408000;
      26302: inst = 32'hc40475f;
      26303: inst = 32'h8220000;
      26304: inst = 32'h10408000;
      26305: inst = 32'hc404760;
      26306: inst = 32'h8220000;
      26307: inst = 32'h10408000;
      26308: inst = 32'hc404761;
      26309: inst = 32'h8220000;
      26310: inst = 32'h10408000;
      26311: inst = 32'hc404762;
      26312: inst = 32'h8220000;
      26313: inst = 32'h10408000;
      26314: inst = 32'hc40476e;
      26315: inst = 32'h8220000;
      26316: inst = 32'h10408000;
      26317: inst = 32'hc40476f;
      26318: inst = 32'h8220000;
      26319: inst = 32'h10408000;
      26320: inst = 32'hc404770;
      26321: inst = 32'h8220000;
      26322: inst = 32'h10408000;
      26323: inst = 32'hc4047ac;
      26324: inst = 32'h8220000;
      26325: inst = 32'h10408000;
      26326: inst = 32'hc4047ad;
      26327: inst = 32'h8220000;
      26328: inst = 32'h10408000;
      26329: inst = 32'hc4047ae;
      26330: inst = 32'h8220000;
      26331: inst = 32'h10408000;
      26332: inst = 32'hc4047bd;
      26333: inst = 32'h8220000;
      26334: inst = 32'h10408000;
      26335: inst = 32'hc4047be;
      26336: inst = 32'h8220000;
      26337: inst = 32'h10408000;
      26338: inst = 32'hc4047bf;
      26339: inst = 32'h8220000;
      26340: inst = 32'h10408000;
      26341: inst = 32'hc4047c0;
      26342: inst = 32'h8220000;
      26343: inst = 32'h10408000;
      26344: inst = 32'hc4047c1;
      26345: inst = 32'h8220000;
      26346: inst = 32'h10408000;
      26347: inst = 32'hc4047c2;
      26348: inst = 32'h8220000;
      26349: inst = 32'h10408000;
      26350: inst = 32'hc4047ce;
      26351: inst = 32'h8220000;
      26352: inst = 32'h10408000;
      26353: inst = 32'hc4047cf;
      26354: inst = 32'h8220000;
      26355: inst = 32'h10408000;
      26356: inst = 32'hc4047d0;
      26357: inst = 32'h8220000;
      26358: inst = 32'h10408000;
      26359: inst = 32'hc40480c;
      26360: inst = 32'h8220000;
      26361: inst = 32'h10408000;
      26362: inst = 32'hc40480d;
      26363: inst = 32'h8220000;
      26364: inst = 32'h10408000;
      26365: inst = 32'hc40480e;
      26366: inst = 32'h8220000;
      26367: inst = 32'h10408000;
      26368: inst = 32'hc40481d;
      26369: inst = 32'h8220000;
      26370: inst = 32'h10408000;
      26371: inst = 32'hc40481e;
      26372: inst = 32'h8220000;
      26373: inst = 32'h10408000;
      26374: inst = 32'hc40481f;
      26375: inst = 32'h8220000;
      26376: inst = 32'h10408000;
      26377: inst = 32'hc404820;
      26378: inst = 32'h8220000;
      26379: inst = 32'h10408000;
      26380: inst = 32'hc404821;
      26381: inst = 32'h8220000;
      26382: inst = 32'h10408000;
      26383: inst = 32'hc404822;
      26384: inst = 32'h8220000;
      26385: inst = 32'h10408000;
      26386: inst = 32'hc40482e;
      26387: inst = 32'h8220000;
      26388: inst = 32'h10408000;
      26389: inst = 32'hc40482f;
      26390: inst = 32'h8220000;
      26391: inst = 32'h10408000;
      26392: inst = 32'hc404830;
      26393: inst = 32'h8220000;
      26394: inst = 32'h10408000;
      26395: inst = 32'hc40486c;
      26396: inst = 32'h8220000;
      26397: inst = 32'h10408000;
      26398: inst = 32'hc40486d;
      26399: inst = 32'h8220000;
      26400: inst = 32'h10408000;
      26401: inst = 32'hc40486e;
      26402: inst = 32'h8220000;
      26403: inst = 32'h10408000;
      26404: inst = 32'hc40487d;
      26405: inst = 32'h8220000;
      26406: inst = 32'h10408000;
      26407: inst = 32'hc40487e;
      26408: inst = 32'h8220000;
      26409: inst = 32'h10408000;
      26410: inst = 32'hc40487f;
      26411: inst = 32'h8220000;
      26412: inst = 32'h10408000;
      26413: inst = 32'hc404880;
      26414: inst = 32'h8220000;
      26415: inst = 32'h10408000;
      26416: inst = 32'hc404881;
      26417: inst = 32'h8220000;
      26418: inst = 32'h10408000;
      26419: inst = 32'hc404882;
      26420: inst = 32'h8220000;
      26421: inst = 32'h10408000;
      26422: inst = 32'hc40488e;
      26423: inst = 32'h8220000;
      26424: inst = 32'h10408000;
      26425: inst = 32'hc40488f;
      26426: inst = 32'h8220000;
      26427: inst = 32'h10408000;
      26428: inst = 32'hc404890;
      26429: inst = 32'h8220000;
      26430: inst = 32'h10408000;
      26431: inst = 32'hc4048cc;
      26432: inst = 32'h8220000;
      26433: inst = 32'h10408000;
      26434: inst = 32'hc4048cd;
      26435: inst = 32'h8220000;
      26436: inst = 32'h10408000;
      26437: inst = 32'hc4048ce;
      26438: inst = 32'h8220000;
      26439: inst = 32'h10408000;
      26440: inst = 32'hc4048dd;
      26441: inst = 32'h8220000;
      26442: inst = 32'h10408000;
      26443: inst = 32'hc4048de;
      26444: inst = 32'h8220000;
      26445: inst = 32'h10408000;
      26446: inst = 32'hc4048df;
      26447: inst = 32'h8220000;
      26448: inst = 32'h10408000;
      26449: inst = 32'hc4048e0;
      26450: inst = 32'h8220000;
      26451: inst = 32'h10408000;
      26452: inst = 32'hc4048e1;
      26453: inst = 32'h8220000;
      26454: inst = 32'h10408000;
      26455: inst = 32'hc4048e2;
      26456: inst = 32'h8220000;
      26457: inst = 32'h10408000;
      26458: inst = 32'hc4048ee;
      26459: inst = 32'h8220000;
      26460: inst = 32'h10408000;
      26461: inst = 32'hc4048ef;
      26462: inst = 32'h8220000;
      26463: inst = 32'h10408000;
      26464: inst = 32'hc4048f0;
      26465: inst = 32'h8220000;
      26466: inst = 32'h10408000;
      26467: inst = 32'hc40492c;
      26468: inst = 32'h8220000;
      26469: inst = 32'h10408000;
      26470: inst = 32'hc40492d;
      26471: inst = 32'h8220000;
      26472: inst = 32'h10408000;
      26473: inst = 32'hc40492e;
      26474: inst = 32'h8220000;
      26475: inst = 32'h10408000;
      26476: inst = 32'hc40493d;
      26477: inst = 32'h8220000;
      26478: inst = 32'h10408000;
      26479: inst = 32'hc40493e;
      26480: inst = 32'h8220000;
      26481: inst = 32'h10408000;
      26482: inst = 32'hc40493f;
      26483: inst = 32'h8220000;
      26484: inst = 32'h10408000;
      26485: inst = 32'hc404940;
      26486: inst = 32'h8220000;
      26487: inst = 32'h10408000;
      26488: inst = 32'hc404941;
      26489: inst = 32'h8220000;
      26490: inst = 32'h10408000;
      26491: inst = 32'hc404942;
      26492: inst = 32'h8220000;
      26493: inst = 32'h10408000;
      26494: inst = 32'hc40494e;
      26495: inst = 32'h8220000;
      26496: inst = 32'h10408000;
      26497: inst = 32'hc40494f;
      26498: inst = 32'h8220000;
      26499: inst = 32'h10408000;
      26500: inst = 32'hc404950;
      26501: inst = 32'h8220000;
      26502: inst = 32'h10408000;
      26503: inst = 32'hc404986;
      26504: inst = 32'h8220000;
      26505: inst = 32'h10408000;
      26506: inst = 32'hc404987;
      26507: inst = 32'h8220000;
      26508: inst = 32'h10408000;
      26509: inst = 32'hc404988;
      26510: inst = 32'h8220000;
      26511: inst = 32'h10408000;
      26512: inst = 32'hc404989;
      26513: inst = 32'h8220000;
      26514: inst = 32'h10408000;
      26515: inst = 32'hc40498a;
      26516: inst = 32'h8220000;
      26517: inst = 32'h10408000;
      26518: inst = 32'hc40498b;
      26519: inst = 32'h8220000;
      26520: inst = 32'h10408000;
      26521: inst = 32'hc40498c;
      26522: inst = 32'h8220000;
      26523: inst = 32'h10408000;
      26524: inst = 32'hc40498d;
      26525: inst = 32'h8220000;
      26526: inst = 32'h10408000;
      26527: inst = 32'hc40498e;
      26528: inst = 32'h8220000;
      26529: inst = 32'h10408000;
      26530: inst = 32'hc40499d;
      26531: inst = 32'h8220000;
      26532: inst = 32'h10408000;
      26533: inst = 32'hc40499e;
      26534: inst = 32'h8220000;
      26535: inst = 32'h10408000;
      26536: inst = 32'hc40499f;
      26537: inst = 32'h8220000;
      26538: inst = 32'h10408000;
      26539: inst = 32'hc4049a0;
      26540: inst = 32'h8220000;
      26541: inst = 32'h10408000;
      26542: inst = 32'hc4049a1;
      26543: inst = 32'h8220000;
      26544: inst = 32'h10408000;
      26545: inst = 32'hc4049a2;
      26546: inst = 32'h8220000;
      26547: inst = 32'h10408000;
      26548: inst = 32'hc4049ae;
      26549: inst = 32'h8220000;
      26550: inst = 32'h10408000;
      26551: inst = 32'hc4049af;
      26552: inst = 32'h8220000;
      26553: inst = 32'h10408000;
      26554: inst = 32'hc4049b0;
      26555: inst = 32'h8220000;
      26556: inst = 32'h10408000;
      26557: inst = 32'hc4049e6;
      26558: inst = 32'h8220000;
      26559: inst = 32'h10408000;
      26560: inst = 32'hc4049e7;
      26561: inst = 32'h8220000;
      26562: inst = 32'h10408000;
      26563: inst = 32'hc4049e8;
      26564: inst = 32'h8220000;
      26565: inst = 32'h10408000;
      26566: inst = 32'hc4049e9;
      26567: inst = 32'h8220000;
      26568: inst = 32'h10408000;
      26569: inst = 32'hc4049ea;
      26570: inst = 32'h8220000;
      26571: inst = 32'h10408000;
      26572: inst = 32'hc4049eb;
      26573: inst = 32'h8220000;
      26574: inst = 32'h10408000;
      26575: inst = 32'hc4049ec;
      26576: inst = 32'h8220000;
      26577: inst = 32'h10408000;
      26578: inst = 32'hc4049ed;
      26579: inst = 32'h8220000;
      26580: inst = 32'h10408000;
      26581: inst = 32'hc4049ee;
      26582: inst = 32'h8220000;
      26583: inst = 32'h10408000;
      26584: inst = 32'hc4049fd;
      26585: inst = 32'h8220000;
      26586: inst = 32'h10408000;
      26587: inst = 32'hc4049fe;
      26588: inst = 32'h8220000;
      26589: inst = 32'h10408000;
      26590: inst = 32'hc4049ff;
      26591: inst = 32'h8220000;
      26592: inst = 32'h10408000;
      26593: inst = 32'hc404a00;
      26594: inst = 32'h8220000;
      26595: inst = 32'h10408000;
      26596: inst = 32'hc404a01;
      26597: inst = 32'h8220000;
      26598: inst = 32'h10408000;
      26599: inst = 32'hc404a02;
      26600: inst = 32'h8220000;
      26601: inst = 32'h10408000;
      26602: inst = 32'hc404a0e;
      26603: inst = 32'h8220000;
      26604: inst = 32'h10408000;
      26605: inst = 32'hc404a0f;
      26606: inst = 32'h8220000;
      26607: inst = 32'h10408000;
      26608: inst = 32'hc404a10;
      26609: inst = 32'h8220000;
      26610: inst = 32'h10408000;
      26611: inst = 32'hc404a46;
      26612: inst = 32'h8220000;
      26613: inst = 32'h10408000;
      26614: inst = 32'hc404a47;
      26615: inst = 32'h8220000;
      26616: inst = 32'h10408000;
      26617: inst = 32'hc404a48;
      26618: inst = 32'h8220000;
      26619: inst = 32'h10408000;
      26620: inst = 32'hc404a49;
      26621: inst = 32'h8220000;
      26622: inst = 32'h10408000;
      26623: inst = 32'hc404a4a;
      26624: inst = 32'h8220000;
      26625: inst = 32'h10408000;
      26626: inst = 32'hc404a4b;
      26627: inst = 32'h8220000;
      26628: inst = 32'h10408000;
      26629: inst = 32'hc404a4c;
      26630: inst = 32'h8220000;
      26631: inst = 32'h10408000;
      26632: inst = 32'hc404a4d;
      26633: inst = 32'h8220000;
      26634: inst = 32'h10408000;
      26635: inst = 32'hc404a4e;
      26636: inst = 32'h8220000;
      26637: inst = 32'h10408000;
      26638: inst = 32'hc404a5d;
      26639: inst = 32'h8220000;
      26640: inst = 32'h10408000;
      26641: inst = 32'hc404a5e;
      26642: inst = 32'h8220000;
      26643: inst = 32'h10408000;
      26644: inst = 32'hc404a5f;
      26645: inst = 32'h8220000;
      26646: inst = 32'h10408000;
      26647: inst = 32'hc404a60;
      26648: inst = 32'h8220000;
      26649: inst = 32'h10408000;
      26650: inst = 32'hc404a61;
      26651: inst = 32'h8220000;
      26652: inst = 32'h10408000;
      26653: inst = 32'hc404a62;
      26654: inst = 32'h8220000;
      26655: inst = 32'h10408000;
      26656: inst = 32'hc404a6e;
      26657: inst = 32'h8220000;
      26658: inst = 32'h10408000;
      26659: inst = 32'hc404a6f;
      26660: inst = 32'h8220000;
      26661: inst = 32'h10408000;
      26662: inst = 32'hc404a70;
      26663: inst = 32'h8220000;
      26664: inst = 32'h10408000;
      26665: inst = 32'hc404abd;
      26666: inst = 32'h8220000;
      26667: inst = 32'h10408000;
      26668: inst = 32'hc404abe;
      26669: inst = 32'h8220000;
      26670: inst = 32'h10408000;
      26671: inst = 32'hc404abf;
      26672: inst = 32'h8220000;
      26673: inst = 32'h10408000;
      26674: inst = 32'hc404ac0;
      26675: inst = 32'h8220000;
      26676: inst = 32'h10408000;
      26677: inst = 32'hc404ac1;
      26678: inst = 32'h8220000;
      26679: inst = 32'h10408000;
      26680: inst = 32'hc404ac2;
      26681: inst = 32'h8220000;
      26682: inst = 32'h10408000;
      26683: inst = 32'hc404ace;
      26684: inst = 32'h8220000;
      26685: inst = 32'h10408000;
      26686: inst = 32'hc404acf;
      26687: inst = 32'h8220000;
      26688: inst = 32'h10408000;
      26689: inst = 32'hc404ad0;
      26690: inst = 32'h8220000;
      26691: inst = 32'h10408000;
      26692: inst = 32'hc404b1d;
      26693: inst = 32'h8220000;
      26694: inst = 32'h10408000;
      26695: inst = 32'hc404b1e;
      26696: inst = 32'h8220000;
      26697: inst = 32'h10408000;
      26698: inst = 32'hc404b1f;
      26699: inst = 32'h8220000;
      26700: inst = 32'h10408000;
      26701: inst = 32'hc404b20;
      26702: inst = 32'h8220000;
      26703: inst = 32'h10408000;
      26704: inst = 32'hc404b21;
      26705: inst = 32'h8220000;
      26706: inst = 32'h10408000;
      26707: inst = 32'hc404b22;
      26708: inst = 32'h8220000;
      26709: inst = 32'h10408000;
      26710: inst = 32'hc404b23;
      26711: inst = 32'h8220000;
      26712: inst = 32'h10408000;
      26713: inst = 32'hc404b24;
      26714: inst = 32'h8220000;
      26715: inst = 32'h10408000;
      26716: inst = 32'hc404b25;
      26717: inst = 32'h8220000;
      26718: inst = 32'h10408000;
      26719: inst = 32'hc404b26;
      26720: inst = 32'h8220000;
      26721: inst = 32'h10408000;
      26722: inst = 32'hc404b27;
      26723: inst = 32'h8220000;
      26724: inst = 32'h10408000;
      26725: inst = 32'hc404b28;
      26726: inst = 32'h8220000;
      26727: inst = 32'h10408000;
      26728: inst = 32'hc404b29;
      26729: inst = 32'h8220000;
      26730: inst = 32'h10408000;
      26731: inst = 32'hc404b2a;
      26732: inst = 32'h8220000;
      26733: inst = 32'h10408000;
      26734: inst = 32'hc404b2b;
      26735: inst = 32'h8220000;
      26736: inst = 32'h10408000;
      26737: inst = 32'hc404b2c;
      26738: inst = 32'h8220000;
      26739: inst = 32'h10408000;
      26740: inst = 32'hc404b2d;
      26741: inst = 32'h8220000;
      26742: inst = 32'h10408000;
      26743: inst = 32'hc404b2e;
      26744: inst = 32'h8220000;
      26745: inst = 32'h10408000;
      26746: inst = 32'hc404b2f;
      26747: inst = 32'h8220000;
      26748: inst = 32'h10408000;
      26749: inst = 32'hc404b30;
      26750: inst = 32'h8220000;
      26751: inst = 32'h10408000;
      26752: inst = 32'hc404b7d;
      26753: inst = 32'h8220000;
      26754: inst = 32'h10408000;
      26755: inst = 32'hc404b7e;
      26756: inst = 32'h8220000;
      26757: inst = 32'h10408000;
      26758: inst = 32'hc404b7f;
      26759: inst = 32'h8220000;
      26760: inst = 32'h10408000;
      26761: inst = 32'hc404b80;
      26762: inst = 32'h8220000;
      26763: inst = 32'h10408000;
      26764: inst = 32'hc404b81;
      26765: inst = 32'h8220000;
      26766: inst = 32'h10408000;
      26767: inst = 32'hc404b82;
      26768: inst = 32'h8220000;
      26769: inst = 32'h10408000;
      26770: inst = 32'hc404b83;
      26771: inst = 32'h8220000;
      26772: inst = 32'h10408000;
      26773: inst = 32'hc404b84;
      26774: inst = 32'h8220000;
      26775: inst = 32'h10408000;
      26776: inst = 32'hc404b85;
      26777: inst = 32'h8220000;
      26778: inst = 32'h10408000;
      26779: inst = 32'hc404b86;
      26780: inst = 32'h8220000;
      26781: inst = 32'h10408000;
      26782: inst = 32'hc404b87;
      26783: inst = 32'h8220000;
      26784: inst = 32'h10408000;
      26785: inst = 32'hc404b88;
      26786: inst = 32'h8220000;
      26787: inst = 32'h10408000;
      26788: inst = 32'hc404b89;
      26789: inst = 32'h8220000;
      26790: inst = 32'h10408000;
      26791: inst = 32'hc404b8a;
      26792: inst = 32'h8220000;
      26793: inst = 32'h10408000;
      26794: inst = 32'hc404b8b;
      26795: inst = 32'h8220000;
      26796: inst = 32'h10408000;
      26797: inst = 32'hc404b8c;
      26798: inst = 32'h8220000;
      26799: inst = 32'h10408000;
      26800: inst = 32'hc404b8d;
      26801: inst = 32'h8220000;
      26802: inst = 32'h10408000;
      26803: inst = 32'hc404b8e;
      26804: inst = 32'h8220000;
      26805: inst = 32'h10408000;
      26806: inst = 32'hc404b8f;
      26807: inst = 32'h8220000;
      26808: inst = 32'h10408000;
      26809: inst = 32'hc404b90;
      26810: inst = 32'h8220000;
      26811: inst = 32'h10408000;
      26812: inst = 32'hc404bdd;
      26813: inst = 32'h8220000;
      26814: inst = 32'h10408000;
      26815: inst = 32'hc404bde;
      26816: inst = 32'h8220000;
      26817: inst = 32'h10408000;
      26818: inst = 32'hc404bdf;
      26819: inst = 32'h8220000;
      26820: inst = 32'h10408000;
      26821: inst = 32'hc404be0;
      26822: inst = 32'h8220000;
      26823: inst = 32'h10408000;
      26824: inst = 32'hc404be1;
      26825: inst = 32'h8220000;
      26826: inst = 32'h10408000;
      26827: inst = 32'hc404be2;
      26828: inst = 32'h8220000;
      26829: inst = 32'h10408000;
      26830: inst = 32'hc404be3;
      26831: inst = 32'h8220000;
      26832: inst = 32'h10408000;
      26833: inst = 32'hc404be4;
      26834: inst = 32'h8220000;
      26835: inst = 32'h10408000;
      26836: inst = 32'hc404be5;
      26837: inst = 32'h8220000;
      26838: inst = 32'h10408000;
      26839: inst = 32'hc404be6;
      26840: inst = 32'h8220000;
      26841: inst = 32'h10408000;
      26842: inst = 32'hc404be7;
      26843: inst = 32'h8220000;
      26844: inst = 32'h10408000;
      26845: inst = 32'hc404be8;
      26846: inst = 32'h8220000;
      26847: inst = 32'h10408000;
      26848: inst = 32'hc404be9;
      26849: inst = 32'h8220000;
      26850: inst = 32'h10408000;
      26851: inst = 32'hc404bea;
      26852: inst = 32'h8220000;
      26853: inst = 32'h10408000;
      26854: inst = 32'hc404beb;
      26855: inst = 32'h8220000;
      26856: inst = 32'h10408000;
      26857: inst = 32'hc404bec;
      26858: inst = 32'h8220000;
      26859: inst = 32'h10408000;
      26860: inst = 32'hc404bed;
      26861: inst = 32'h8220000;
      26862: inst = 32'h10408000;
      26863: inst = 32'hc404bee;
      26864: inst = 32'h8220000;
      26865: inst = 32'h10408000;
      26866: inst = 32'hc404bef;
      26867: inst = 32'h8220000;
      26868: inst = 32'h10408000;
      26869: inst = 32'hc404bf0;
      26870: inst = 32'h8220000;
      26871: inst = 32'h10408000;
      26872: inst = 32'hc404c3d;
      26873: inst = 32'h8220000;
      26874: inst = 32'h10408000;
      26875: inst = 32'hc404c3e;
      26876: inst = 32'h8220000;
      26877: inst = 32'h10408000;
      26878: inst = 32'hc404c3f;
      26879: inst = 32'h8220000;
      26880: inst = 32'h10408000;
      26881: inst = 32'hc404c40;
      26882: inst = 32'h8220000;
      26883: inst = 32'h10408000;
      26884: inst = 32'hc404c41;
      26885: inst = 32'h8220000;
      26886: inst = 32'h10408000;
      26887: inst = 32'hc404c42;
      26888: inst = 32'h8220000;
      26889: inst = 32'h10408000;
      26890: inst = 32'hc404c9d;
      26891: inst = 32'h8220000;
      26892: inst = 32'h10408000;
      26893: inst = 32'hc404c9e;
      26894: inst = 32'h8220000;
      26895: inst = 32'h10408000;
      26896: inst = 32'hc404c9f;
      26897: inst = 32'h8220000;
      26898: inst = 32'h10408000;
      26899: inst = 32'hc404ca0;
      26900: inst = 32'h8220000;
      26901: inst = 32'h10408000;
      26902: inst = 32'hc404ca1;
      26903: inst = 32'h8220000;
      26904: inst = 32'h10408000;
      26905: inst = 32'hc404ca2;
      26906: inst = 32'h8220000;
      26907: inst = 32'h10408000;
      26908: inst = 32'hc404cfd;
      26909: inst = 32'h8220000;
      26910: inst = 32'h10408000;
      26911: inst = 32'hc404cfe;
      26912: inst = 32'h8220000;
      26913: inst = 32'h10408000;
      26914: inst = 32'hc404cff;
      26915: inst = 32'h8220000;
      26916: inst = 32'h10408000;
      26917: inst = 32'hc404d00;
      26918: inst = 32'h8220000;
      26919: inst = 32'h10408000;
      26920: inst = 32'hc404d01;
      26921: inst = 32'h8220000;
      26922: inst = 32'h10408000;
      26923: inst = 32'hc404d02;
      26924: inst = 32'h8220000;
      26925: inst = 32'h10408000;
      26926: inst = 32'hc404d25;
      26927: inst = 32'h8220000;
      26928: inst = 32'h10408000;
      26929: inst = 32'hc404d26;
      26930: inst = 32'h8220000;
      26931: inst = 32'h10408000;
      26932: inst = 32'hc404d27;
      26933: inst = 32'h8220000;
      26934: inst = 32'h10408000;
      26935: inst = 32'hc404d28;
      26936: inst = 32'h8220000;
      26937: inst = 32'h10408000;
      26938: inst = 32'hc404d29;
      26939: inst = 32'h8220000;
      26940: inst = 32'h10408000;
      26941: inst = 32'hc404d2a;
      26942: inst = 32'h8220000;
      26943: inst = 32'h10408000;
      26944: inst = 32'hc404d2b;
      26945: inst = 32'h8220000;
      26946: inst = 32'h10408000;
      26947: inst = 32'hc404d2c;
      26948: inst = 32'h8220000;
      26949: inst = 32'h10408000;
      26950: inst = 32'hc404d2d;
      26951: inst = 32'h8220000;
      26952: inst = 32'h10408000;
      26953: inst = 32'hc404d2e;
      26954: inst = 32'h8220000;
      26955: inst = 32'h10408000;
      26956: inst = 32'hc404d2f;
      26957: inst = 32'h8220000;
      26958: inst = 32'h10408000;
      26959: inst = 32'hc404d30;
      26960: inst = 32'h8220000;
      26961: inst = 32'h10408000;
      26962: inst = 32'hc404d31;
      26963: inst = 32'h8220000;
      26964: inst = 32'h10408000;
      26965: inst = 32'hc404d32;
      26966: inst = 32'h8220000;
      26967: inst = 32'h10408000;
      26968: inst = 32'hc404d33;
      26969: inst = 32'h8220000;
      26970: inst = 32'h10408000;
      26971: inst = 32'hc404d34;
      26972: inst = 32'h8220000;
      26973: inst = 32'h10408000;
      26974: inst = 32'hc404d35;
      26975: inst = 32'h8220000;
      26976: inst = 32'h10408000;
      26977: inst = 32'hc404d36;
      26978: inst = 32'h8220000;
      26979: inst = 32'h10408000;
      26980: inst = 32'hc404d37;
      26981: inst = 32'h8220000;
      26982: inst = 32'h10408000;
      26983: inst = 32'hc404d38;
      26984: inst = 32'h8220000;
      26985: inst = 32'h10408000;
      26986: inst = 32'hc404d39;
      26987: inst = 32'h8220000;
      26988: inst = 32'h10408000;
      26989: inst = 32'hc404d3a;
      26990: inst = 32'h8220000;
      26991: inst = 32'h10408000;
      26992: inst = 32'hc404d5d;
      26993: inst = 32'h8220000;
      26994: inst = 32'h10408000;
      26995: inst = 32'hc404d5e;
      26996: inst = 32'h8220000;
      26997: inst = 32'h10408000;
      26998: inst = 32'hc404d5f;
      26999: inst = 32'h8220000;
      27000: inst = 32'h10408000;
      27001: inst = 32'hc404d60;
      27002: inst = 32'h8220000;
      27003: inst = 32'h10408000;
      27004: inst = 32'hc404d61;
      27005: inst = 32'h8220000;
      27006: inst = 32'h10408000;
      27007: inst = 32'hc404d62;
      27008: inst = 32'h8220000;
      27009: inst = 32'h10408000;
      27010: inst = 32'hc404d85;
      27011: inst = 32'h8220000;
      27012: inst = 32'h10408000;
      27013: inst = 32'hc404d86;
      27014: inst = 32'h8220000;
      27015: inst = 32'h10408000;
      27016: inst = 32'hc404d87;
      27017: inst = 32'h8220000;
      27018: inst = 32'h10408000;
      27019: inst = 32'hc404d88;
      27020: inst = 32'h8220000;
      27021: inst = 32'h10408000;
      27022: inst = 32'hc404d89;
      27023: inst = 32'h8220000;
      27024: inst = 32'h10408000;
      27025: inst = 32'hc404d8a;
      27026: inst = 32'h8220000;
      27027: inst = 32'h10408000;
      27028: inst = 32'hc404d8b;
      27029: inst = 32'h8220000;
      27030: inst = 32'h10408000;
      27031: inst = 32'hc404d8c;
      27032: inst = 32'h8220000;
      27033: inst = 32'h10408000;
      27034: inst = 32'hc404d8d;
      27035: inst = 32'h8220000;
      27036: inst = 32'h10408000;
      27037: inst = 32'hc404d8e;
      27038: inst = 32'h8220000;
      27039: inst = 32'h10408000;
      27040: inst = 32'hc404d8f;
      27041: inst = 32'h8220000;
      27042: inst = 32'h10408000;
      27043: inst = 32'hc404d90;
      27044: inst = 32'h8220000;
      27045: inst = 32'h10408000;
      27046: inst = 32'hc404d91;
      27047: inst = 32'h8220000;
      27048: inst = 32'h10408000;
      27049: inst = 32'hc404d92;
      27050: inst = 32'h8220000;
      27051: inst = 32'h10408000;
      27052: inst = 32'hc404d93;
      27053: inst = 32'h8220000;
      27054: inst = 32'h10408000;
      27055: inst = 32'hc404d94;
      27056: inst = 32'h8220000;
      27057: inst = 32'h10408000;
      27058: inst = 32'hc404d95;
      27059: inst = 32'h8220000;
      27060: inst = 32'h10408000;
      27061: inst = 32'hc404d96;
      27062: inst = 32'h8220000;
      27063: inst = 32'h10408000;
      27064: inst = 32'hc404d97;
      27065: inst = 32'h8220000;
      27066: inst = 32'h10408000;
      27067: inst = 32'hc404d98;
      27068: inst = 32'h8220000;
      27069: inst = 32'h10408000;
      27070: inst = 32'hc404d99;
      27071: inst = 32'h8220000;
      27072: inst = 32'h10408000;
      27073: inst = 32'hc404d9a;
      27074: inst = 32'h8220000;
      27075: inst = 32'h10408000;
      27076: inst = 32'hc404dbd;
      27077: inst = 32'h8220000;
      27078: inst = 32'h10408000;
      27079: inst = 32'hc404dbe;
      27080: inst = 32'h8220000;
      27081: inst = 32'h10408000;
      27082: inst = 32'hc404dbf;
      27083: inst = 32'h8220000;
      27084: inst = 32'h10408000;
      27085: inst = 32'hc404dc0;
      27086: inst = 32'h8220000;
      27087: inst = 32'h10408000;
      27088: inst = 32'hc404dc1;
      27089: inst = 32'h8220000;
      27090: inst = 32'h10408000;
      27091: inst = 32'hc404dc2;
      27092: inst = 32'h8220000;
      27093: inst = 32'h10408000;
      27094: inst = 32'hc404de5;
      27095: inst = 32'h8220000;
      27096: inst = 32'h10408000;
      27097: inst = 32'hc404de6;
      27098: inst = 32'h8220000;
      27099: inst = 32'h10408000;
      27100: inst = 32'hc404de7;
      27101: inst = 32'h8220000;
      27102: inst = 32'h10408000;
      27103: inst = 32'hc404de8;
      27104: inst = 32'h8220000;
      27105: inst = 32'h10408000;
      27106: inst = 32'hc404de9;
      27107: inst = 32'h8220000;
      27108: inst = 32'h10408000;
      27109: inst = 32'hc404dea;
      27110: inst = 32'h8220000;
      27111: inst = 32'h10408000;
      27112: inst = 32'hc404deb;
      27113: inst = 32'h8220000;
      27114: inst = 32'h10408000;
      27115: inst = 32'hc404dec;
      27116: inst = 32'h8220000;
      27117: inst = 32'h10408000;
      27118: inst = 32'hc404ded;
      27119: inst = 32'h8220000;
      27120: inst = 32'h10408000;
      27121: inst = 32'hc404dee;
      27122: inst = 32'h8220000;
      27123: inst = 32'h10408000;
      27124: inst = 32'hc404def;
      27125: inst = 32'h8220000;
      27126: inst = 32'h10408000;
      27127: inst = 32'hc404df0;
      27128: inst = 32'h8220000;
      27129: inst = 32'h10408000;
      27130: inst = 32'hc404df1;
      27131: inst = 32'h8220000;
      27132: inst = 32'h10408000;
      27133: inst = 32'hc404df2;
      27134: inst = 32'h8220000;
      27135: inst = 32'h10408000;
      27136: inst = 32'hc404df3;
      27137: inst = 32'h8220000;
      27138: inst = 32'h10408000;
      27139: inst = 32'hc404df4;
      27140: inst = 32'h8220000;
      27141: inst = 32'h10408000;
      27142: inst = 32'hc404df5;
      27143: inst = 32'h8220000;
      27144: inst = 32'h10408000;
      27145: inst = 32'hc404df6;
      27146: inst = 32'h8220000;
      27147: inst = 32'h10408000;
      27148: inst = 32'hc404df7;
      27149: inst = 32'h8220000;
      27150: inst = 32'h10408000;
      27151: inst = 32'hc404df8;
      27152: inst = 32'h8220000;
      27153: inst = 32'h10408000;
      27154: inst = 32'hc404df9;
      27155: inst = 32'h8220000;
      27156: inst = 32'h10408000;
      27157: inst = 32'hc404dfa;
      27158: inst = 32'h8220000;
      27159: inst = 32'h10408000;
      27160: inst = 32'hc404e1d;
      27161: inst = 32'h8220000;
      27162: inst = 32'h10408000;
      27163: inst = 32'hc404e1e;
      27164: inst = 32'h8220000;
      27165: inst = 32'h10408000;
      27166: inst = 32'hc404e1f;
      27167: inst = 32'h8220000;
      27168: inst = 32'h10408000;
      27169: inst = 32'hc404e20;
      27170: inst = 32'h8220000;
      27171: inst = 32'h10408000;
      27172: inst = 32'hc404e21;
      27173: inst = 32'h8220000;
      27174: inst = 32'h10408000;
      27175: inst = 32'hc404e22;
      27176: inst = 32'h8220000;
      27177: inst = 32'h10408000;
      27178: inst = 32'hc404e58;
      27179: inst = 32'h8220000;
      27180: inst = 32'h10408000;
      27181: inst = 32'hc404e59;
      27182: inst = 32'h8220000;
      27183: inst = 32'h10408000;
      27184: inst = 32'hc404e5a;
      27185: inst = 32'h8220000;
      27186: inst = 32'h10408000;
      27187: inst = 32'hc404e7d;
      27188: inst = 32'h8220000;
      27189: inst = 32'h10408000;
      27190: inst = 32'hc404e7e;
      27191: inst = 32'h8220000;
      27192: inst = 32'h10408000;
      27193: inst = 32'hc404e7f;
      27194: inst = 32'h8220000;
      27195: inst = 32'h10408000;
      27196: inst = 32'hc404e80;
      27197: inst = 32'h8220000;
      27198: inst = 32'h10408000;
      27199: inst = 32'hc404e81;
      27200: inst = 32'h8220000;
      27201: inst = 32'h10408000;
      27202: inst = 32'hc404e82;
      27203: inst = 32'h8220000;
      27204: inst = 32'h10408000;
      27205: inst = 32'hc404eb8;
      27206: inst = 32'h8220000;
      27207: inst = 32'h10408000;
      27208: inst = 32'hc404eb9;
      27209: inst = 32'h8220000;
      27210: inst = 32'h10408000;
      27211: inst = 32'hc404eba;
      27212: inst = 32'h8220000;
      27213: inst = 32'h10408000;
      27214: inst = 32'hc404edd;
      27215: inst = 32'h8220000;
      27216: inst = 32'h10408000;
      27217: inst = 32'hc404ede;
      27218: inst = 32'h8220000;
      27219: inst = 32'h10408000;
      27220: inst = 32'hc404edf;
      27221: inst = 32'h8220000;
      27222: inst = 32'h10408000;
      27223: inst = 32'hc404ee0;
      27224: inst = 32'h8220000;
      27225: inst = 32'h10408000;
      27226: inst = 32'hc404ee1;
      27227: inst = 32'h8220000;
      27228: inst = 32'h10408000;
      27229: inst = 32'hc404ee2;
      27230: inst = 32'h8220000;
      27231: inst = 32'h10408000;
      27232: inst = 32'hc404f18;
      27233: inst = 32'h8220000;
      27234: inst = 32'h10408000;
      27235: inst = 32'hc404f19;
      27236: inst = 32'h8220000;
      27237: inst = 32'h10408000;
      27238: inst = 32'hc404f1a;
      27239: inst = 32'h8220000;
      27240: inst = 32'h10408000;
      27241: inst = 32'hc404f3d;
      27242: inst = 32'h8220000;
      27243: inst = 32'h10408000;
      27244: inst = 32'hc404f3e;
      27245: inst = 32'h8220000;
      27246: inst = 32'h10408000;
      27247: inst = 32'hc404f3f;
      27248: inst = 32'h8220000;
      27249: inst = 32'h10408000;
      27250: inst = 32'hc404f40;
      27251: inst = 32'h8220000;
      27252: inst = 32'h10408000;
      27253: inst = 32'hc404f41;
      27254: inst = 32'h8220000;
      27255: inst = 32'h10408000;
      27256: inst = 32'hc404f42;
      27257: inst = 32'h8220000;
      27258: inst = 32'h10408000;
      27259: inst = 32'hc404f78;
      27260: inst = 32'h8220000;
      27261: inst = 32'h10408000;
      27262: inst = 32'hc404f79;
      27263: inst = 32'h8220000;
      27264: inst = 32'h10408000;
      27265: inst = 32'hc404f7a;
      27266: inst = 32'h8220000;
      27267: inst = 32'h10408000;
      27268: inst = 32'hc404f9d;
      27269: inst = 32'h8220000;
      27270: inst = 32'h10408000;
      27271: inst = 32'hc404f9e;
      27272: inst = 32'h8220000;
      27273: inst = 32'h10408000;
      27274: inst = 32'hc404f9f;
      27275: inst = 32'h8220000;
      27276: inst = 32'h10408000;
      27277: inst = 32'hc404fa0;
      27278: inst = 32'h8220000;
      27279: inst = 32'h10408000;
      27280: inst = 32'hc404fa1;
      27281: inst = 32'h8220000;
      27282: inst = 32'h10408000;
      27283: inst = 32'hc404fa2;
      27284: inst = 32'h8220000;
      27285: inst = 32'h10408000;
      27286: inst = 32'hc404fd8;
      27287: inst = 32'h8220000;
      27288: inst = 32'h10408000;
      27289: inst = 32'hc404fd9;
      27290: inst = 32'h8220000;
      27291: inst = 32'h10408000;
      27292: inst = 32'hc404fda;
      27293: inst = 32'h8220000;
      27294: inst = 32'h10408000;
      27295: inst = 32'hc404ffd;
      27296: inst = 32'h8220000;
      27297: inst = 32'h10408000;
      27298: inst = 32'hc404ffe;
      27299: inst = 32'h8220000;
      27300: inst = 32'h10408000;
      27301: inst = 32'hc404fff;
      27302: inst = 32'h8220000;
      27303: inst = 32'h10408000;
      27304: inst = 32'hc405000;
      27305: inst = 32'h8220000;
      27306: inst = 32'h10408000;
      27307: inst = 32'hc405001;
      27308: inst = 32'h8220000;
      27309: inst = 32'h10408000;
      27310: inst = 32'hc405002;
      27311: inst = 32'h8220000;
      27312: inst = 32'h10408000;
      27313: inst = 32'hc405038;
      27314: inst = 32'h8220000;
      27315: inst = 32'h10408000;
      27316: inst = 32'hc405039;
      27317: inst = 32'h8220000;
      27318: inst = 32'h10408000;
      27319: inst = 32'hc40503a;
      27320: inst = 32'h8220000;
      27321: inst = 32'h10408000;
      27322: inst = 32'hc40505d;
      27323: inst = 32'h8220000;
      27324: inst = 32'h10408000;
      27325: inst = 32'hc40505e;
      27326: inst = 32'h8220000;
      27327: inst = 32'h10408000;
      27328: inst = 32'hc40505f;
      27329: inst = 32'h8220000;
      27330: inst = 32'h10408000;
      27331: inst = 32'hc405060;
      27332: inst = 32'h8220000;
      27333: inst = 32'h10408000;
      27334: inst = 32'hc405061;
      27335: inst = 32'h8220000;
      27336: inst = 32'h10408000;
      27337: inst = 32'hc405062;
      27338: inst = 32'h8220000;
      27339: inst = 32'h10408000;
      27340: inst = 32'hc405098;
      27341: inst = 32'h8220000;
      27342: inst = 32'h10408000;
      27343: inst = 32'hc405099;
      27344: inst = 32'h8220000;
      27345: inst = 32'h10408000;
      27346: inst = 32'hc40509a;
      27347: inst = 32'h8220000;
      27348: inst = 32'h10408000;
      27349: inst = 32'hc40509b;
      27350: inst = 32'h8220000;
      27351: inst = 32'h10408000;
      27352: inst = 32'hc40509c;
      27353: inst = 32'h8220000;
      27354: inst = 32'h10408000;
      27355: inst = 32'hc40509d;
      27356: inst = 32'h8220000;
      27357: inst = 32'h10408000;
      27358: inst = 32'hc40509e;
      27359: inst = 32'h8220000;
      27360: inst = 32'h10408000;
      27361: inst = 32'hc40509f;
      27362: inst = 32'h8220000;
      27363: inst = 32'h10408000;
      27364: inst = 32'hc4050a0;
      27365: inst = 32'h8220000;
      27366: inst = 32'h10408000;
      27367: inst = 32'hc4050a1;
      27368: inst = 32'h8220000;
      27369: inst = 32'h10408000;
      27370: inst = 32'hc4050a2;
      27371: inst = 32'h8220000;
      27372: inst = 32'h10408000;
      27373: inst = 32'hc4050a3;
      27374: inst = 32'h8220000;
      27375: inst = 32'h10408000;
      27376: inst = 32'hc4050a4;
      27377: inst = 32'h8220000;
      27378: inst = 32'h10408000;
      27379: inst = 32'hc4050a5;
      27380: inst = 32'h8220000;
      27381: inst = 32'h10408000;
      27382: inst = 32'hc4050a6;
      27383: inst = 32'h8220000;
      27384: inst = 32'h10408000;
      27385: inst = 32'hc4050a7;
      27386: inst = 32'h8220000;
      27387: inst = 32'h10408000;
      27388: inst = 32'hc4050a8;
      27389: inst = 32'h8220000;
      27390: inst = 32'h10408000;
      27391: inst = 32'hc4050a9;
      27392: inst = 32'h8220000;
      27393: inst = 32'h10408000;
      27394: inst = 32'hc4050aa;
      27395: inst = 32'h8220000;
      27396: inst = 32'h10408000;
      27397: inst = 32'hc4050ab;
      27398: inst = 32'h8220000;
      27399: inst = 32'h10408000;
      27400: inst = 32'hc4050ac;
      27401: inst = 32'h8220000;
      27402: inst = 32'h10408000;
      27403: inst = 32'hc4050ad;
      27404: inst = 32'h8220000;
      27405: inst = 32'h10408000;
      27406: inst = 32'hc4050ae;
      27407: inst = 32'h8220000;
      27408: inst = 32'h10408000;
      27409: inst = 32'hc4050af;
      27410: inst = 32'h8220000;
      27411: inst = 32'h10408000;
      27412: inst = 32'hc4050b0;
      27413: inst = 32'h8220000;
      27414: inst = 32'h10408000;
      27415: inst = 32'hc4050b1;
      27416: inst = 32'h8220000;
      27417: inst = 32'h10408000;
      27418: inst = 32'hc4050b2;
      27419: inst = 32'h8220000;
      27420: inst = 32'h10408000;
      27421: inst = 32'hc4050b3;
      27422: inst = 32'h8220000;
      27423: inst = 32'h10408000;
      27424: inst = 32'hc4050b4;
      27425: inst = 32'h8220000;
      27426: inst = 32'h10408000;
      27427: inst = 32'hc4050b5;
      27428: inst = 32'h8220000;
      27429: inst = 32'h10408000;
      27430: inst = 32'hc4050b6;
      27431: inst = 32'h8220000;
      27432: inst = 32'h10408000;
      27433: inst = 32'hc4050b7;
      27434: inst = 32'h8220000;
      27435: inst = 32'h10408000;
      27436: inst = 32'hc4050b8;
      27437: inst = 32'h8220000;
      27438: inst = 32'h10408000;
      27439: inst = 32'hc4050b9;
      27440: inst = 32'h8220000;
      27441: inst = 32'h10408000;
      27442: inst = 32'hc4050ba;
      27443: inst = 32'h8220000;
      27444: inst = 32'h10408000;
      27445: inst = 32'hc4050bb;
      27446: inst = 32'h8220000;
      27447: inst = 32'h10408000;
      27448: inst = 32'hc4050bc;
      27449: inst = 32'h8220000;
      27450: inst = 32'h10408000;
      27451: inst = 32'hc4050bd;
      27452: inst = 32'h8220000;
      27453: inst = 32'h10408000;
      27454: inst = 32'hc4050be;
      27455: inst = 32'h8220000;
      27456: inst = 32'h10408000;
      27457: inst = 32'hc4050bf;
      27458: inst = 32'h8220000;
      27459: inst = 32'h10408000;
      27460: inst = 32'hc4050c0;
      27461: inst = 32'h8220000;
      27462: inst = 32'h10408000;
      27463: inst = 32'hc4050c1;
      27464: inst = 32'h8220000;
      27465: inst = 32'h10408000;
      27466: inst = 32'hc4050c2;
      27467: inst = 32'h8220000;
      27468: inst = 32'h10408000;
      27469: inst = 32'hc4050f8;
      27470: inst = 32'h8220000;
      27471: inst = 32'h10408000;
      27472: inst = 32'hc4050f9;
      27473: inst = 32'h8220000;
      27474: inst = 32'h10408000;
      27475: inst = 32'hc4050fa;
      27476: inst = 32'h8220000;
      27477: inst = 32'h10408000;
      27478: inst = 32'hc4050fb;
      27479: inst = 32'h8220000;
      27480: inst = 32'h10408000;
      27481: inst = 32'hc4050fc;
      27482: inst = 32'h8220000;
      27483: inst = 32'h10408000;
      27484: inst = 32'hc4050fd;
      27485: inst = 32'h8220000;
      27486: inst = 32'h10408000;
      27487: inst = 32'hc4050fe;
      27488: inst = 32'h8220000;
      27489: inst = 32'h10408000;
      27490: inst = 32'hc4050ff;
      27491: inst = 32'h8220000;
      27492: inst = 32'h10408000;
      27493: inst = 32'hc405100;
      27494: inst = 32'h8220000;
      27495: inst = 32'h10408000;
      27496: inst = 32'hc405101;
      27497: inst = 32'h8220000;
      27498: inst = 32'h10408000;
      27499: inst = 32'hc405102;
      27500: inst = 32'h8220000;
      27501: inst = 32'h10408000;
      27502: inst = 32'hc405103;
      27503: inst = 32'h8220000;
      27504: inst = 32'h10408000;
      27505: inst = 32'hc405104;
      27506: inst = 32'h8220000;
      27507: inst = 32'h10408000;
      27508: inst = 32'hc405105;
      27509: inst = 32'h8220000;
      27510: inst = 32'h10408000;
      27511: inst = 32'hc405106;
      27512: inst = 32'h8220000;
      27513: inst = 32'h10408000;
      27514: inst = 32'hc405107;
      27515: inst = 32'h8220000;
      27516: inst = 32'h10408000;
      27517: inst = 32'hc405108;
      27518: inst = 32'h8220000;
      27519: inst = 32'h10408000;
      27520: inst = 32'hc405109;
      27521: inst = 32'h8220000;
      27522: inst = 32'h10408000;
      27523: inst = 32'hc40510a;
      27524: inst = 32'h8220000;
      27525: inst = 32'h10408000;
      27526: inst = 32'hc40510b;
      27527: inst = 32'h8220000;
      27528: inst = 32'h10408000;
      27529: inst = 32'hc40510c;
      27530: inst = 32'h8220000;
      27531: inst = 32'h10408000;
      27532: inst = 32'hc40510d;
      27533: inst = 32'h8220000;
      27534: inst = 32'h10408000;
      27535: inst = 32'hc40510e;
      27536: inst = 32'h8220000;
      27537: inst = 32'h10408000;
      27538: inst = 32'hc40510f;
      27539: inst = 32'h8220000;
      27540: inst = 32'h10408000;
      27541: inst = 32'hc405110;
      27542: inst = 32'h8220000;
      27543: inst = 32'h10408000;
      27544: inst = 32'hc405111;
      27545: inst = 32'h8220000;
      27546: inst = 32'h10408000;
      27547: inst = 32'hc405112;
      27548: inst = 32'h8220000;
      27549: inst = 32'h10408000;
      27550: inst = 32'hc405113;
      27551: inst = 32'h8220000;
      27552: inst = 32'h10408000;
      27553: inst = 32'hc405114;
      27554: inst = 32'h8220000;
      27555: inst = 32'h10408000;
      27556: inst = 32'hc405115;
      27557: inst = 32'h8220000;
      27558: inst = 32'h10408000;
      27559: inst = 32'hc405116;
      27560: inst = 32'h8220000;
      27561: inst = 32'h10408000;
      27562: inst = 32'hc405117;
      27563: inst = 32'h8220000;
      27564: inst = 32'h10408000;
      27565: inst = 32'hc405118;
      27566: inst = 32'h8220000;
      27567: inst = 32'h10408000;
      27568: inst = 32'hc405119;
      27569: inst = 32'h8220000;
      27570: inst = 32'h10408000;
      27571: inst = 32'hc40511a;
      27572: inst = 32'h8220000;
      27573: inst = 32'h10408000;
      27574: inst = 32'hc40511b;
      27575: inst = 32'h8220000;
      27576: inst = 32'h10408000;
      27577: inst = 32'hc40511c;
      27578: inst = 32'h8220000;
      27579: inst = 32'h10408000;
      27580: inst = 32'hc40511d;
      27581: inst = 32'h8220000;
      27582: inst = 32'h10408000;
      27583: inst = 32'hc40511e;
      27584: inst = 32'h8220000;
      27585: inst = 32'h10408000;
      27586: inst = 32'hc40511f;
      27587: inst = 32'h8220000;
      27588: inst = 32'h10408000;
      27589: inst = 32'hc405120;
      27590: inst = 32'h8220000;
      27591: inst = 32'h10408000;
      27592: inst = 32'hc405121;
      27593: inst = 32'h8220000;
      27594: inst = 32'h10408000;
      27595: inst = 32'hc405122;
      27596: inst = 32'h8220000;
      27597: inst = 32'h10408000;
      27598: inst = 32'hc405136;
      27599: inst = 32'h8220000;
      27600: inst = 32'h10408000;
      27601: inst = 32'hc405137;
      27602: inst = 32'h8220000;
      27603: inst = 32'h10408000;
      27604: inst = 32'hc405138;
      27605: inst = 32'h8220000;
      27606: inst = 32'h10408000;
      27607: inst = 32'hc405158;
      27608: inst = 32'h8220000;
      27609: inst = 32'h10408000;
      27610: inst = 32'hc405159;
      27611: inst = 32'h8220000;
      27612: inst = 32'h10408000;
      27613: inst = 32'hc40515a;
      27614: inst = 32'h8220000;
      27615: inst = 32'h10408000;
      27616: inst = 32'hc40515b;
      27617: inst = 32'h8220000;
      27618: inst = 32'h10408000;
      27619: inst = 32'hc40515c;
      27620: inst = 32'h8220000;
      27621: inst = 32'h10408000;
      27622: inst = 32'hc40515d;
      27623: inst = 32'h8220000;
      27624: inst = 32'h10408000;
      27625: inst = 32'hc40515e;
      27626: inst = 32'h8220000;
      27627: inst = 32'h10408000;
      27628: inst = 32'hc40515f;
      27629: inst = 32'h8220000;
      27630: inst = 32'h10408000;
      27631: inst = 32'hc405160;
      27632: inst = 32'h8220000;
      27633: inst = 32'h10408000;
      27634: inst = 32'hc405161;
      27635: inst = 32'h8220000;
      27636: inst = 32'h10408000;
      27637: inst = 32'hc405162;
      27638: inst = 32'h8220000;
      27639: inst = 32'h10408000;
      27640: inst = 32'hc405163;
      27641: inst = 32'h8220000;
      27642: inst = 32'h10408000;
      27643: inst = 32'hc405164;
      27644: inst = 32'h8220000;
      27645: inst = 32'h10408000;
      27646: inst = 32'hc405165;
      27647: inst = 32'h8220000;
      27648: inst = 32'h10408000;
      27649: inst = 32'hc405166;
      27650: inst = 32'h8220000;
      27651: inst = 32'h10408000;
      27652: inst = 32'hc405167;
      27653: inst = 32'h8220000;
      27654: inst = 32'h10408000;
      27655: inst = 32'hc405168;
      27656: inst = 32'h8220000;
      27657: inst = 32'h10408000;
      27658: inst = 32'hc405169;
      27659: inst = 32'h8220000;
      27660: inst = 32'h10408000;
      27661: inst = 32'hc40516a;
      27662: inst = 32'h8220000;
      27663: inst = 32'h10408000;
      27664: inst = 32'hc40516b;
      27665: inst = 32'h8220000;
      27666: inst = 32'h10408000;
      27667: inst = 32'hc40516c;
      27668: inst = 32'h8220000;
      27669: inst = 32'h10408000;
      27670: inst = 32'hc40516d;
      27671: inst = 32'h8220000;
      27672: inst = 32'h10408000;
      27673: inst = 32'hc40516e;
      27674: inst = 32'h8220000;
      27675: inst = 32'h10408000;
      27676: inst = 32'hc40516f;
      27677: inst = 32'h8220000;
      27678: inst = 32'h10408000;
      27679: inst = 32'hc405170;
      27680: inst = 32'h8220000;
      27681: inst = 32'h10408000;
      27682: inst = 32'hc405171;
      27683: inst = 32'h8220000;
      27684: inst = 32'h10408000;
      27685: inst = 32'hc405172;
      27686: inst = 32'h8220000;
      27687: inst = 32'h10408000;
      27688: inst = 32'hc405173;
      27689: inst = 32'h8220000;
      27690: inst = 32'h10408000;
      27691: inst = 32'hc405174;
      27692: inst = 32'h8220000;
      27693: inst = 32'h10408000;
      27694: inst = 32'hc405175;
      27695: inst = 32'h8220000;
      27696: inst = 32'h10408000;
      27697: inst = 32'hc405176;
      27698: inst = 32'h8220000;
      27699: inst = 32'h10408000;
      27700: inst = 32'hc405177;
      27701: inst = 32'h8220000;
      27702: inst = 32'h10408000;
      27703: inst = 32'hc405178;
      27704: inst = 32'h8220000;
      27705: inst = 32'h10408000;
      27706: inst = 32'hc405179;
      27707: inst = 32'h8220000;
      27708: inst = 32'h10408000;
      27709: inst = 32'hc40517a;
      27710: inst = 32'h8220000;
      27711: inst = 32'h10408000;
      27712: inst = 32'hc40517b;
      27713: inst = 32'h8220000;
      27714: inst = 32'h10408000;
      27715: inst = 32'hc40517c;
      27716: inst = 32'h8220000;
      27717: inst = 32'h10408000;
      27718: inst = 32'hc40517d;
      27719: inst = 32'h8220000;
      27720: inst = 32'h10408000;
      27721: inst = 32'hc40517e;
      27722: inst = 32'h8220000;
      27723: inst = 32'h10408000;
      27724: inst = 32'hc40517f;
      27725: inst = 32'h8220000;
      27726: inst = 32'h10408000;
      27727: inst = 32'hc405180;
      27728: inst = 32'h8220000;
      27729: inst = 32'h10408000;
      27730: inst = 32'hc405181;
      27731: inst = 32'h8220000;
      27732: inst = 32'h10408000;
      27733: inst = 32'hc405182;
      27734: inst = 32'h8220000;
      27735: inst = 32'h10408000;
      27736: inst = 32'hc405196;
      27737: inst = 32'h8220000;
      27738: inst = 32'h10408000;
      27739: inst = 32'hc405197;
      27740: inst = 32'h8220000;
      27741: inst = 32'h10408000;
      27742: inst = 32'hc405198;
      27743: inst = 32'h8220000;
      27744: inst = 32'h10408000;
      27745: inst = 32'hc4051dd;
      27746: inst = 32'h8220000;
      27747: inst = 32'h10408000;
      27748: inst = 32'hc4051de;
      27749: inst = 32'h8220000;
      27750: inst = 32'h10408000;
      27751: inst = 32'hc4051df;
      27752: inst = 32'h8220000;
      27753: inst = 32'h10408000;
      27754: inst = 32'hc4051e0;
      27755: inst = 32'h8220000;
      27756: inst = 32'h10408000;
      27757: inst = 32'hc4051e1;
      27758: inst = 32'h8220000;
      27759: inst = 32'h10408000;
      27760: inst = 32'hc4051e2;
      27761: inst = 32'h8220000;
      27762: inst = 32'h10408000;
      27763: inst = 32'hc4051f6;
      27764: inst = 32'h8220000;
      27765: inst = 32'h10408000;
      27766: inst = 32'hc4051f7;
      27767: inst = 32'h8220000;
      27768: inst = 32'h10408000;
      27769: inst = 32'hc4051f8;
      27770: inst = 32'h8220000;
      27771: inst = 32'h10408000;
      27772: inst = 32'hc40523d;
      27773: inst = 32'h8220000;
      27774: inst = 32'h10408000;
      27775: inst = 32'hc40523e;
      27776: inst = 32'h8220000;
      27777: inst = 32'h10408000;
      27778: inst = 32'hc40523f;
      27779: inst = 32'h8220000;
      27780: inst = 32'h10408000;
      27781: inst = 32'hc405240;
      27782: inst = 32'h8220000;
      27783: inst = 32'h10408000;
      27784: inst = 32'hc405241;
      27785: inst = 32'h8220000;
      27786: inst = 32'h10408000;
      27787: inst = 32'hc405242;
      27788: inst = 32'h8220000;
      27789: inst = 32'h10408000;
      27790: inst = 32'hc405256;
      27791: inst = 32'h8220000;
      27792: inst = 32'h10408000;
      27793: inst = 32'hc405257;
      27794: inst = 32'h8220000;
      27795: inst = 32'h10408000;
      27796: inst = 32'hc405258;
      27797: inst = 32'h8220000;
      27798: inst = 32'h10408000;
      27799: inst = 32'hc40529d;
      27800: inst = 32'h8220000;
      27801: inst = 32'h10408000;
      27802: inst = 32'hc40529e;
      27803: inst = 32'h8220000;
      27804: inst = 32'h10408000;
      27805: inst = 32'hc40529f;
      27806: inst = 32'h8220000;
      27807: inst = 32'h10408000;
      27808: inst = 32'hc4052a0;
      27809: inst = 32'h8220000;
      27810: inst = 32'h10408000;
      27811: inst = 32'hc4052a1;
      27812: inst = 32'h8220000;
      27813: inst = 32'h10408000;
      27814: inst = 32'hc4052a2;
      27815: inst = 32'h8220000;
      27816: inst = 32'h10408000;
      27817: inst = 32'hc4052b6;
      27818: inst = 32'h8220000;
      27819: inst = 32'h10408000;
      27820: inst = 32'hc4052b7;
      27821: inst = 32'h8220000;
      27822: inst = 32'h10408000;
      27823: inst = 32'hc4052b8;
      27824: inst = 32'h8220000;
      27825: inst = 32'h10408000;
      27826: inst = 32'hc4052fd;
      27827: inst = 32'h8220000;
      27828: inst = 32'h10408000;
      27829: inst = 32'hc4052fe;
      27830: inst = 32'h8220000;
      27831: inst = 32'h10408000;
      27832: inst = 32'hc4052ff;
      27833: inst = 32'h8220000;
      27834: inst = 32'h10408000;
      27835: inst = 32'hc405300;
      27836: inst = 32'h8220000;
      27837: inst = 32'h10408000;
      27838: inst = 32'hc405301;
      27839: inst = 32'h8220000;
      27840: inst = 32'h10408000;
      27841: inst = 32'hc405302;
      27842: inst = 32'h8220000;
      27843: inst = 32'h10408000;
      27844: inst = 32'hc405316;
      27845: inst = 32'h8220000;
      27846: inst = 32'h10408000;
      27847: inst = 32'hc405317;
      27848: inst = 32'h8220000;
      27849: inst = 32'h10408000;
      27850: inst = 32'hc405318;
      27851: inst = 32'h8220000;
      27852: inst = 32'h10408000;
      27853: inst = 32'hc40535d;
      27854: inst = 32'h8220000;
      27855: inst = 32'h10408000;
      27856: inst = 32'hc40535e;
      27857: inst = 32'h8220000;
      27858: inst = 32'h10408000;
      27859: inst = 32'hc40535f;
      27860: inst = 32'h8220000;
      27861: inst = 32'h10408000;
      27862: inst = 32'hc405360;
      27863: inst = 32'h8220000;
      27864: inst = 32'h10408000;
      27865: inst = 32'hc405361;
      27866: inst = 32'h8220000;
      27867: inst = 32'h10408000;
      27868: inst = 32'hc405362;
      27869: inst = 32'h8220000;
      27870: inst = 32'h10408000;
      27871: inst = 32'hc405376;
      27872: inst = 32'h8220000;
      27873: inst = 32'h10408000;
      27874: inst = 32'hc405377;
      27875: inst = 32'h8220000;
      27876: inst = 32'h10408000;
      27877: inst = 32'hc405378;
      27878: inst = 32'h8220000;
      27879: inst = 32'h10408000;
      27880: inst = 32'hc4053bd;
      27881: inst = 32'h8220000;
      27882: inst = 32'h10408000;
      27883: inst = 32'hc4053be;
      27884: inst = 32'h8220000;
      27885: inst = 32'h10408000;
      27886: inst = 32'hc4053bf;
      27887: inst = 32'h8220000;
      27888: inst = 32'h10408000;
      27889: inst = 32'hc4053c0;
      27890: inst = 32'h8220000;
      27891: inst = 32'h10408000;
      27892: inst = 32'hc4053c1;
      27893: inst = 32'h8220000;
      27894: inst = 32'h10408000;
      27895: inst = 32'hc4053c2;
      27896: inst = 32'h8220000;
      27897: inst = 32'h10408000;
      27898: inst = 32'hc4053d6;
      27899: inst = 32'h8220000;
      27900: inst = 32'h10408000;
      27901: inst = 32'hc4053d7;
      27902: inst = 32'h8220000;
      27903: inst = 32'h10408000;
      27904: inst = 32'hc4053d8;
      27905: inst = 32'h8220000;
      27906: inst = 32'h10408000;
      27907: inst = 32'hc40541d;
      27908: inst = 32'h8220000;
      27909: inst = 32'h10408000;
      27910: inst = 32'hc40541e;
      27911: inst = 32'h8220000;
      27912: inst = 32'h10408000;
      27913: inst = 32'hc40541f;
      27914: inst = 32'h8220000;
      27915: inst = 32'h10408000;
      27916: inst = 32'hc405420;
      27917: inst = 32'h8220000;
      27918: inst = 32'h10408000;
      27919: inst = 32'hc405421;
      27920: inst = 32'h8220000;
      27921: inst = 32'h10408000;
      27922: inst = 32'hc405422;
      27923: inst = 32'h8220000;
      27924: inst = 32'h10408000;
      27925: inst = 32'hc405436;
      27926: inst = 32'h8220000;
      27927: inst = 32'h10408000;
      27928: inst = 32'hc405437;
      27929: inst = 32'h8220000;
      27930: inst = 32'h10408000;
      27931: inst = 32'hc405438;
      27932: inst = 32'h8220000;
      27933: inst = 32'h10408000;
      27934: inst = 32'hc405439;
      27935: inst = 32'h8220000;
      27936: inst = 32'h10408000;
      27937: inst = 32'hc40543a;
      27938: inst = 32'h8220000;
      27939: inst = 32'h10408000;
      27940: inst = 32'hc40543b;
      27941: inst = 32'h8220000;
      27942: inst = 32'h10408000;
      27943: inst = 32'hc40543c;
      27944: inst = 32'h8220000;
      27945: inst = 32'h10408000;
      27946: inst = 32'hc40543d;
      27947: inst = 32'h8220000;
      27948: inst = 32'h10408000;
      27949: inst = 32'hc40543e;
      27950: inst = 32'h8220000;
      27951: inst = 32'h10408000;
      27952: inst = 32'hc40543f;
      27953: inst = 32'h8220000;
      27954: inst = 32'h10408000;
      27955: inst = 32'hc405440;
      27956: inst = 32'h8220000;
      27957: inst = 32'h10408000;
      27958: inst = 32'hc405441;
      27959: inst = 32'h8220000;
      27960: inst = 32'h10408000;
      27961: inst = 32'hc405442;
      27962: inst = 32'h8220000;
      27963: inst = 32'h10408000;
      27964: inst = 32'hc405443;
      27965: inst = 32'h8220000;
      27966: inst = 32'h10408000;
      27967: inst = 32'hc405444;
      27968: inst = 32'h8220000;
      27969: inst = 32'h10408000;
      27970: inst = 32'hc405445;
      27971: inst = 32'h8220000;
      27972: inst = 32'h10408000;
      27973: inst = 32'hc405446;
      27974: inst = 32'h8220000;
      27975: inst = 32'h10408000;
      27976: inst = 32'hc405447;
      27977: inst = 32'h8220000;
      27978: inst = 32'h10408000;
      27979: inst = 32'hc405448;
      27980: inst = 32'h8220000;
      27981: inst = 32'h10408000;
      27982: inst = 32'hc405449;
      27983: inst = 32'h8220000;
      27984: inst = 32'h10408000;
      27985: inst = 32'hc40547d;
      27986: inst = 32'h8220000;
      27987: inst = 32'h10408000;
      27988: inst = 32'hc40547e;
      27989: inst = 32'h8220000;
      27990: inst = 32'h10408000;
      27991: inst = 32'hc40547f;
      27992: inst = 32'h8220000;
      27993: inst = 32'h10408000;
      27994: inst = 32'hc405480;
      27995: inst = 32'h8220000;
      27996: inst = 32'h10408000;
      27997: inst = 32'hc405481;
      27998: inst = 32'h8220000;
      27999: inst = 32'h10408000;
      28000: inst = 32'hc405482;
      28001: inst = 32'h8220000;
      28002: inst = 32'h10408000;
      28003: inst = 32'hc405496;
      28004: inst = 32'h8220000;
      28005: inst = 32'h10408000;
      28006: inst = 32'hc405497;
      28007: inst = 32'h8220000;
      28008: inst = 32'h10408000;
      28009: inst = 32'hc405498;
      28010: inst = 32'h8220000;
      28011: inst = 32'h10408000;
      28012: inst = 32'hc405499;
      28013: inst = 32'h8220000;
      28014: inst = 32'h10408000;
      28015: inst = 32'hc40549a;
      28016: inst = 32'h8220000;
      28017: inst = 32'h10408000;
      28018: inst = 32'hc40549b;
      28019: inst = 32'h8220000;
      28020: inst = 32'h10408000;
      28021: inst = 32'hc40549c;
      28022: inst = 32'h8220000;
      28023: inst = 32'h10408000;
      28024: inst = 32'hc40549d;
      28025: inst = 32'h8220000;
      28026: inst = 32'h10408000;
      28027: inst = 32'hc40549e;
      28028: inst = 32'h8220000;
      28029: inst = 32'h10408000;
      28030: inst = 32'hc40549f;
      28031: inst = 32'h8220000;
      28032: inst = 32'h10408000;
      28033: inst = 32'hc4054a0;
      28034: inst = 32'h8220000;
      28035: inst = 32'h10408000;
      28036: inst = 32'hc4054a1;
      28037: inst = 32'h8220000;
      28038: inst = 32'h10408000;
      28039: inst = 32'hc4054a2;
      28040: inst = 32'h8220000;
      28041: inst = 32'h10408000;
      28042: inst = 32'hc4054a3;
      28043: inst = 32'h8220000;
      28044: inst = 32'h10408000;
      28045: inst = 32'hc4054a4;
      28046: inst = 32'h8220000;
      28047: inst = 32'h10408000;
      28048: inst = 32'hc4054a5;
      28049: inst = 32'h8220000;
      28050: inst = 32'h10408000;
      28051: inst = 32'hc4054a6;
      28052: inst = 32'h8220000;
      28053: inst = 32'h10408000;
      28054: inst = 32'hc4054a7;
      28055: inst = 32'h8220000;
      28056: inst = 32'h10408000;
      28057: inst = 32'hc4054a8;
      28058: inst = 32'h8220000;
      28059: inst = 32'h10408000;
      28060: inst = 32'hc4054a9;
      28061: inst = 32'h8220000;
      28062: inst = 32'h10408000;
      28063: inst = 32'hc4054dd;
      28064: inst = 32'h8220000;
      28065: inst = 32'h10408000;
      28066: inst = 32'hc4054de;
      28067: inst = 32'h8220000;
      28068: inst = 32'h10408000;
      28069: inst = 32'hc4054df;
      28070: inst = 32'h8220000;
      28071: inst = 32'h10408000;
      28072: inst = 32'hc4054e0;
      28073: inst = 32'h8220000;
      28074: inst = 32'h10408000;
      28075: inst = 32'hc4054e1;
      28076: inst = 32'h8220000;
      28077: inst = 32'h10408000;
      28078: inst = 32'hc4054e2;
      28079: inst = 32'h8220000;
      28080: inst = 32'h10408000;
      28081: inst = 32'hc4054f6;
      28082: inst = 32'h8220000;
      28083: inst = 32'h10408000;
      28084: inst = 32'hc4054f7;
      28085: inst = 32'h8220000;
      28086: inst = 32'h10408000;
      28087: inst = 32'hc4054f8;
      28088: inst = 32'h8220000;
      28089: inst = 32'h10408000;
      28090: inst = 32'hc4054f9;
      28091: inst = 32'h8220000;
      28092: inst = 32'h10408000;
      28093: inst = 32'hc4054fa;
      28094: inst = 32'h8220000;
      28095: inst = 32'h10408000;
      28096: inst = 32'hc4054fb;
      28097: inst = 32'h8220000;
      28098: inst = 32'h10408000;
      28099: inst = 32'hc4054fc;
      28100: inst = 32'h8220000;
      28101: inst = 32'h10408000;
      28102: inst = 32'hc4054fd;
      28103: inst = 32'h8220000;
      28104: inst = 32'h10408000;
      28105: inst = 32'hc4054fe;
      28106: inst = 32'h8220000;
      28107: inst = 32'h10408000;
      28108: inst = 32'hc4054ff;
      28109: inst = 32'h8220000;
      28110: inst = 32'h10408000;
      28111: inst = 32'hc405500;
      28112: inst = 32'h8220000;
      28113: inst = 32'h10408000;
      28114: inst = 32'hc405501;
      28115: inst = 32'h8220000;
      28116: inst = 32'h10408000;
      28117: inst = 32'hc405502;
      28118: inst = 32'h8220000;
      28119: inst = 32'h10408000;
      28120: inst = 32'hc405503;
      28121: inst = 32'h8220000;
      28122: inst = 32'h10408000;
      28123: inst = 32'hc405504;
      28124: inst = 32'h8220000;
      28125: inst = 32'h10408000;
      28126: inst = 32'hc405505;
      28127: inst = 32'h8220000;
      28128: inst = 32'h10408000;
      28129: inst = 32'hc405506;
      28130: inst = 32'h8220000;
      28131: inst = 32'h10408000;
      28132: inst = 32'hc405507;
      28133: inst = 32'h8220000;
      28134: inst = 32'h10408000;
      28135: inst = 32'hc405508;
      28136: inst = 32'h8220000;
      28137: inst = 32'h10408000;
      28138: inst = 32'hc405509;
      28139: inst = 32'h8220000;
      28140: inst = 32'h10408000;
      28141: inst = 32'hc40553d;
      28142: inst = 32'h8220000;
      28143: inst = 32'h10408000;
      28144: inst = 32'hc40553e;
      28145: inst = 32'h8220000;
      28146: inst = 32'h10408000;
      28147: inst = 32'hc40553f;
      28148: inst = 32'h8220000;
      28149: inst = 32'h10408000;
      28150: inst = 32'hc405540;
      28151: inst = 32'h8220000;
      28152: inst = 32'h10408000;
      28153: inst = 32'hc405541;
      28154: inst = 32'h8220000;
      28155: inst = 32'h10408000;
      28156: inst = 32'hc405542;
      28157: inst = 32'h8220000;
      28158: inst = 32'h10408000;
      28159: inst = 32'hc405556;
      28160: inst = 32'h8220000;
      28161: inst = 32'h10408000;
      28162: inst = 32'hc405557;
      28163: inst = 32'h8220000;
      28164: inst = 32'h10408000;
      28165: inst = 32'hc405558;
      28166: inst = 32'h8220000;
      28167: inst = 32'h10408000;
      28168: inst = 32'hc40559d;
      28169: inst = 32'h8220000;
      28170: inst = 32'h10408000;
      28171: inst = 32'hc40559e;
      28172: inst = 32'h8220000;
      28173: inst = 32'h10408000;
      28174: inst = 32'hc40559f;
      28175: inst = 32'h8220000;
      28176: inst = 32'h10408000;
      28177: inst = 32'hc4055a0;
      28178: inst = 32'h8220000;
      28179: inst = 32'h10408000;
      28180: inst = 32'hc4055a1;
      28181: inst = 32'h8220000;
      28182: inst = 32'h10408000;
      28183: inst = 32'hc4055a2;
      28184: inst = 32'h8220000;
      28185: inst = 32'h10408000;
      28186: inst = 32'hc4055b6;
      28187: inst = 32'h8220000;
      28188: inst = 32'h10408000;
      28189: inst = 32'hc4055b7;
      28190: inst = 32'h8220000;
      28191: inst = 32'h10408000;
      28192: inst = 32'hc4055b8;
      28193: inst = 32'h8220000;
      28194: inst = 32'h10408000;
      28195: inst = 32'hc4055fd;
      28196: inst = 32'h8220000;
      28197: inst = 32'h10408000;
      28198: inst = 32'hc4055fe;
      28199: inst = 32'h8220000;
      28200: inst = 32'h10408000;
      28201: inst = 32'hc4055ff;
      28202: inst = 32'h8220000;
      28203: inst = 32'h10408000;
      28204: inst = 32'hc405600;
      28205: inst = 32'h8220000;
      28206: inst = 32'h10408000;
      28207: inst = 32'hc405601;
      28208: inst = 32'h8220000;
      28209: inst = 32'h10408000;
      28210: inst = 32'hc405602;
      28211: inst = 32'h8220000;
      28212: inst = 32'h10408000;
      28213: inst = 32'hc405616;
      28214: inst = 32'h8220000;
      28215: inst = 32'h10408000;
      28216: inst = 32'hc405617;
      28217: inst = 32'h8220000;
      28218: inst = 32'h10408000;
      28219: inst = 32'hc405618;
      28220: inst = 32'h8220000;
      28221: inst = 32'h10408000;
      28222: inst = 32'hc40565d;
      28223: inst = 32'h8220000;
      28224: inst = 32'h10408000;
      28225: inst = 32'hc40565e;
      28226: inst = 32'h8220000;
      28227: inst = 32'h10408000;
      28228: inst = 32'hc40565f;
      28229: inst = 32'h8220000;
      28230: inst = 32'h10408000;
      28231: inst = 32'hc405660;
      28232: inst = 32'h8220000;
      28233: inst = 32'h10408000;
      28234: inst = 32'hc405661;
      28235: inst = 32'h8220000;
      28236: inst = 32'h10408000;
      28237: inst = 32'hc405662;
      28238: inst = 32'h8220000;
      28239: inst = 32'h10408000;
      28240: inst = 32'hc405676;
      28241: inst = 32'h8220000;
      28242: inst = 32'h10408000;
      28243: inst = 32'hc405677;
      28244: inst = 32'h8220000;
      28245: inst = 32'h10408000;
      28246: inst = 32'hc405678;
      28247: inst = 32'h8220000;
      28248: inst = 32'h10408000;
      28249: inst = 32'hc4056b7;
      28250: inst = 32'h8220000;
      28251: inst = 32'h10408000;
      28252: inst = 32'hc4056b8;
      28253: inst = 32'h8220000;
      28254: inst = 32'h10408000;
      28255: inst = 32'hc4056b9;
      28256: inst = 32'h8220000;
      28257: inst = 32'h10408000;
      28258: inst = 32'hc4056bd;
      28259: inst = 32'h8220000;
      28260: inst = 32'h10408000;
      28261: inst = 32'hc4056be;
      28262: inst = 32'h8220000;
      28263: inst = 32'h10408000;
      28264: inst = 32'hc4056bf;
      28265: inst = 32'h8220000;
      28266: inst = 32'h10408000;
      28267: inst = 32'hc4056c0;
      28268: inst = 32'h8220000;
      28269: inst = 32'h10408000;
      28270: inst = 32'hc4056c1;
      28271: inst = 32'h8220000;
      28272: inst = 32'h10408000;
      28273: inst = 32'hc4056c2;
      28274: inst = 32'h8220000;
      28275: inst = 32'h10408000;
      28276: inst = 32'hc4056c3;
      28277: inst = 32'h8220000;
      28278: inst = 32'h10408000;
      28279: inst = 32'hc4056c4;
      28280: inst = 32'h8220000;
      28281: inst = 32'h10408000;
      28282: inst = 32'hc4056c5;
      28283: inst = 32'h8220000;
      28284: inst = 32'h10408000;
      28285: inst = 32'hc4056c6;
      28286: inst = 32'h8220000;
      28287: inst = 32'h10408000;
      28288: inst = 32'hc4056c7;
      28289: inst = 32'h8220000;
      28290: inst = 32'h10408000;
      28291: inst = 32'hc4056c8;
      28292: inst = 32'h8220000;
      28293: inst = 32'h10408000;
      28294: inst = 32'hc4056c9;
      28295: inst = 32'h8220000;
      28296: inst = 32'h10408000;
      28297: inst = 32'hc4056d4;
      28298: inst = 32'h8220000;
      28299: inst = 32'h10408000;
      28300: inst = 32'hc4056d5;
      28301: inst = 32'h8220000;
      28302: inst = 32'h10408000;
      28303: inst = 32'hc4056d6;
      28304: inst = 32'h8220000;
      28305: inst = 32'h10408000;
      28306: inst = 32'hc4056d7;
      28307: inst = 32'h8220000;
      28308: inst = 32'h10408000;
      28309: inst = 32'hc4056d8;
      28310: inst = 32'h8220000;
      28311: inst = 32'h10408000;
      28312: inst = 32'hc4056d9;
      28313: inst = 32'h8220000;
      28314: inst = 32'h10408000;
      28315: inst = 32'hc4056da;
      28316: inst = 32'h8220000;
      28317: inst = 32'h10408000;
      28318: inst = 32'hc4056db;
      28319: inst = 32'h8220000;
      28320: inst = 32'h10408000;
      28321: inst = 32'hc4056dc;
      28322: inst = 32'h8220000;
      28323: inst = 32'h10408000;
      28324: inst = 32'hc4056dd;
      28325: inst = 32'h8220000;
      28326: inst = 32'h10408000;
      28327: inst = 32'hc4056de;
      28328: inst = 32'h8220000;
      28329: inst = 32'h10408000;
      28330: inst = 32'hc4056df;
      28331: inst = 32'h8220000;
      28332: inst = 32'h10408000;
      28333: inst = 32'hc4056e0;
      28334: inst = 32'h8220000;
      28335: inst = 32'h10408000;
      28336: inst = 32'hc4056e1;
      28337: inst = 32'h8220000;
      28338: inst = 32'h10408000;
      28339: inst = 32'hc4056e2;
      28340: inst = 32'h8220000;
      28341: inst = 32'h10408000;
      28342: inst = 32'hc4056e3;
      28343: inst = 32'h8220000;
      28344: inst = 32'h10408000;
      28345: inst = 32'hc4056e4;
      28346: inst = 32'h8220000;
      28347: inst = 32'h10408000;
      28348: inst = 32'hc4056e5;
      28349: inst = 32'h8220000;
      28350: inst = 32'h10408000;
      28351: inst = 32'hc4056e6;
      28352: inst = 32'h8220000;
      28353: inst = 32'h10408000;
      28354: inst = 32'hc4056e7;
      28355: inst = 32'h8220000;
      28356: inst = 32'h10408000;
      28357: inst = 32'hc4056e8;
      28358: inst = 32'h8220000;
      28359: inst = 32'h10408000;
      28360: inst = 32'hc4056e9;
      28361: inst = 32'h8220000;
      28362: inst = 32'h10408000;
      28363: inst = 32'hc4056ea;
      28364: inst = 32'h8220000;
      28365: inst = 32'h10408000;
      28366: inst = 32'hc4056eb;
      28367: inst = 32'h8220000;
      28368: inst = 32'h10408000;
      28369: inst = 32'hc4056ec;
      28370: inst = 32'h8220000;
      28371: inst = 32'h10408000;
      28372: inst = 32'hc4056ed;
      28373: inst = 32'h8220000;
      28374: inst = 32'h10408000;
      28375: inst = 32'hc4056ee;
      28376: inst = 32'h8220000;
      28377: inst = 32'h10408000;
      28378: inst = 32'hc4056ef;
      28379: inst = 32'h8220000;
      28380: inst = 32'h10408000;
      28381: inst = 32'hc4056f0;
      28382: inst = 32'h8220000;
      28383: inst = 32'h10408000;
      28384: inst = 32'hc4056f1;
      28385: inst = 32'h8220000;
      28386: inst = 32'h10408000;
      28387: inst = 32'hc4056f2;
      28388: inst = 32'h8220000;
      28389: inst = 32'h10408000;
      28390: inst = 32'hc4056f3;
      28391: inst = 32'h8220000;
      28392: inst = 32'h10408000;
      28393: inst = 32'hc4056f4;
      28394: inst = 32'h8220000;
      28395: inst = 32'h10408000;
      28396: inst = 32'hc4056f5;
      28397: inst = 32'h8220000;
      28398: inst = 32'h10408000;
      28399: inst = 32'hc4056f6;
      28400: inst = 32'h8220000;
      28401: inst = 32'h10408000;
      28402: inst = 32'hc4056f7;
      28403: inst = 32'h8220000;
      28404: inst = 32'h10408000;
      28405: inst = 32'hc4056f8;
      28406: inst = 32'h8220000;
      28407: inst = 32'h10408000;
      28408: inst = 32'hc4056f9;
      28409: inst = 32'h8220000;
      28410: inst = 32'h10408000;
      28411: inst = 32'hc4056fa;
      28412: inst = 32'h8220000;
      28413: inst = 32'h10408000;
      28414: inst = 32'hc4056fb;
      28415: inst = 32'h8220000;
      28416: inst = 32'h10408000;
      28417: inst = 32'hc4056fc;
      28418: inst = 32'h8220000;
      28419: inst = 32'h10408000;
      28420: inst = 32'hc4056fd;
      28421: inst = 32'h8220000;
      28422: inst = 32'h10408000;
      28423: inst = 32'hc405701;
      28424: inst = 32'h8220000;
      28425: inst = 32'h10408000;
      28426: inst = 32'hc405702;
      28427: inst = 32'h8220000;
      28428: inst = 32'h10408000;
      28429: inst = 32'hc405703;
      28430: inst = 32'h8220000;
      28431: inst = 32'h10408000;
      28432: inst = 32'hc405704;
      28433: inst = 32'h8220000;
      28434: inst = 32'h10408000;
      28435: inst = 32'hc405705;
      28436: inst = 32'h8220000;
      28437: inst = 32'h10408000;
      28438: inst = 32'hc405706;
      28439: inst = 32'h8220000;
      28440: inst = 32'h10408000;
      28441: inst = 32'hc405707;
      28442: inst = 32'h8220000;
      28443: inst = 32'h10408000;
      28444: inst = 32'hc405708;
      28445: inst = 32'h8220000;
      28446: inst = 32'h10408000;
      28447: inst = 32'hc405709;
      28448: inst = 32'h8220000;
      28449: inst = 32'h10408000;
      28450: inst = 32'hc40570a;
      28451: inst = 32'h8220000;
      28452: inst = 32'h10408000;
      28453: inst = 32'hc40570b;
      28454: inst = 32'h8220000;
      28455: inst = 32'h10408000;
      28456: inst = 32'hc40570c;
      28457: inst = 32'h8220000;
      28458: inst = 32'h10408000;
      28459: inst = 32'hc40570d;
      28460: inst = 32'h8220000;
      28461: inst = 32'h10408000;
      28462: inst = 32'hc40570e;
      28463: inst = 32'h8220000;
      28464: inst = 32'h10408000;
      28465: inst = 32'hc40570f;
      28466: inst = 32'h8220000;
      28467: inst = 32'h10408000;
      28468: inst = 32'hc405710;
      28469: inst = 32'h8220000;
      28470: inst = 32'h10408000;
      28471: inst = 32'hc405717;
      28472: inst = 32'h8220000;
      28473: inst = 32'h10408000;
      28474: inst = 32'hc405718;
      28475: inst = 32'h8220000;
      28476: inst = 32'h10408000;
      28477: inst = 32'hc405719;
      28478: inst = 32'h8220000;
      28479: inst = 32'h10408000;
      28480: inst = 32'hc40571d;
      28481: inst = 32'h8220000;
      28482: inst = 32'h10408000;
      28483: inst = 32'hc40571e;
      28484: inst = 32'h8220000;
      28485: inst = 32'h10408000;
      28486: inst = 32'hc40571f;
      28487: inst = 32'h8220000;
      28488: inst = 32'h10408000;
      28489: inst = 32'hc405720;
      28490: inst = 32'h8220000;
      28491: inst = 32'h10408000;
      28492: inst = 32'hc405721;
      28493: inst = 32'h8220000;
      28494: inst = 32'h10408000;
      28495: inst = 32'hc405722;
      28496: inst = 32'h8220000;
      28497: inst = 32'h10408000;
      28498: inst = 32'hc405723;
      28499: inst = 32'h8220000;
      28500: inst = 32'h10408000;
      28501: inst = 32'hc405724;
      28502: inst = 32'h8220000;
      28503: inst = 32'h10408000;
      28504: inst = 32'hc405725;
      28505: inst = 32'h8220000;
      28506: inst = 32'h10408000;
      28507: inst = 32'hc405726;
      28508: inst = 32'h8220000;
      28509: inst = 32'h10408000;
      28510: inst = 32'hc405727;
      28511: inst = 32'h8220000;
      28512: inst = 32'h10408000;
      28513: inst = 32'hc405728;
      28514: inst = 32'h8220000;
      28515: inst = 32'h10408000;
      28516: inst = 32'hc405729;
      28517: inst = 32'h8220000;
      28518: inst = 32'h10408000;
      28519: inst = 32'hc40572a;
      28520: inst = 32'h8220000;
      28521: inst = 32'h10408000;
      28522: inst = 32'hc40572b;
      28523: inst = 32'h8220000;
      28524: inst = 32'h10408000;
      28525: inst = 32'hc40572c;
      28526: inst = 32'h8220000;
      28527: inst = 32'h10408000;
      28528: inst = 32'hc40572d;
      28529: inst = 32'h8220000;
      28530: inst = 32'h10408000;
      28531: inst = 32'hc40572e;
      28532: inst = 32'h8220000;
      28533: inst = 32'h10408000;
      28534: inst = 32'hc40572f;
      28535: inst = 32'h8220000;
      28536: inst = 32'h10408000;
      28537: inst = 32'hc405730;
      28538: inst = 32'h8220000;
      28539: inst = 32'h10408000;
      28540: inst = 32'hc405731;
      28541: inst = 32'h8220000;
      28542: inst = 32'h10408000;
      28543: inst = 32'hc405732;
      28544: inst = 32'h8220000;
      28545: inst = 32'h10408000;
      28546: inst = 32'hc405733;
      28547: inst = 32'h8220000;
      28548: inst = 32'h10408000;
      28549: inst = 32'hc405734;
      28550: inst = 32'h8220000;
      28551: inst = 32'h10408000;
      28552: inst = 32'hc405735;
      28553: inst = 32'h8220000;
      28554: inst = 32'h10408000;
      28555: inst = 32'hc405736;
      28556: inst = 32'h8220000;
      28557: inst = 32'h10408000;
      28558: inst = 32'hc405737;
      28559: inst = 32'h8220000;
      28560: inst = 32'h10408000;
      28561: inst = 32'hc405738;
      28562: inst = 32'h8220000;
      28563: inst = 32'h10408000;
      28564: inst = 32'hc405739;
      28565: inst = 32'h8220000;
      28566: inst = 32'h10408000;
      28567: inst = 32'hc40573a;
      28568: inst = 32'h8220000;
      28569: inst = 32'h10408000;
      28570: inst = 32'hc40573b;
      28571: inst = 32'h8220000;
      28572: inst = 32'h10408000;
      28573: inst = 32'hc40573c;
      28574: inst = 32'h8220000;
      28575: inst = 32'h10408000;
      28576: inst = 32'hc40573d;
      28577: inst = 32'h8220000;
      28578: inst = 32'h10408000;
      28579: inst = 32'hc40573e;
      28580: inst = 32'h8220000;
      28581: inst = 32'h10408000;
      28582: inst = 32'hc40573f;
      28583: inst = 32'h8220000;
      28584: inst = 32'h10408000;
      28585: inst = 32'hc405740;
      28586: inst = 32'h8220000;
      28587: inst = 32'h10408000;
      28588: inst = 32'hc405741;
      28589: inst = 32'h8220000;
      28590: inst = 32'h10408000;
      28591: inst = 32'hc405742;
      28592: inst = 32'h8220000;
      28593: inst = 32'h10408000;
      28594: inst = 32'hc405743;
      28595: inst = 32'h8220000;
      28596: inst = 32'h10408000;
      28597: inst = 32'hc405744;
      28598: inst = 32'h8220000;
      28599: inst = 32'h10408000;
      28600: inst = 32'hc405745;
      28601: inst = 32'h8220000;
      28602: inst = 32'h10408000;
      28603: inst = 32'hc405746;
      28604: inst = 32'h8220000;
      28605: inst = 32'h10408000;
      28606: inst = 32'hc405747;
      28607: inst = 32'h8220000;
      28608: inst = 32'h10408000;
      28609: inst = 32'hc405748;
      28610: inst = 32'h8220000;
      28611: inst = 32'h10408000;
      28612: inst = 32'hc405749;
      28613: inst = 32'h8220000;
      28614: inst = 32'h10408000;
      28615: inst = 32'hc40574a;
      28616: inst = 32'h8220000;
      28617: inst = 32'h10408000;
      28618: inst = 32'hc40574b;
      28619: inst = 32'h8220000;
      28620: inst = 32'h10408000;
      28621: inst = 32'hc40574c;
      28622: inst = 32'h8220000;
      28623: inst = 32'h10408000;
      28624: inst = 32'hc40574d;
      28625: inst = 32'h8220000;
      28626: inst = 32'h10408000;
      28627: inst = 32'hc40574e;
      28628: inst = 32'h8220000;
      28629: inst = 32'h10408000;
      28630: inst = 32'hc40574f;
      28631: inst = 32'h8220000;
      28632: inst = 32'h10408000;
      28633: inst = 32'hc405750;
      28634: inst = 32'h8220000;
      28635: inst = 32'h10408000;
      28636: inst = 32'hc405751;
      28637: inst = 32'h8220000;
      28638: inst = 32'h10408000;
      28639: inst = 32'hc405752;
      28640: inst = 32'h8220000;
      28641: inst = 32'h10408000;
      28642: inst = 32'hc405753;
      28643: inst = 32'h8220000;
      28644: inst = 32'h10408000;
      28645: inst = 32'hc405754;
      28646: inst = 32'h8220000;
      28647: inst = 32'h10408000;
      28648: inst = 32'hc405755;
      28649: inst = 32'h8220000;
      28650: inst = 32'h10408000;
      28651: inst = 32'hc405756;
      28652: inst = 32'h8220000;
      28653: inst = 32'h10408000;
      28654: inst = 32'hc405757;
      28655: inst = 32'h8220000;
      28656: inst = 32'h10408000;
      28657: inst = 32'hc405758;
      28658: inst = 32'h8220000;
      28659: inst = 32'h10408000;
      28660: inst = 32'hc405759;
      28661: inst = 32'h8220000;
      28662: inst = 32'h10408000;
      28663: inst = 32'hc40575a;
      28664: inst = 32'h8220000;
      28665: inst = 32'h10408000;
      28666: inst = 32'hc40575b;
      28667: inst = 32'h8220000;
      28668: inst = 32'h10408000;
      28669: inst = 32'hc40575c;
      28670: inst = 32'h8220000;
      28671: inst = 32'h10408000;
      28672: inst = 32'hc40575d;
      28673: inst = 32'h8220000;
      28674: inst = 32'h10408000;
      28675: inst = 32'hc40575e;
      28676: inst = 32'h8220000;
      28677: inst = 32'h10408000;
      28678: inst = 32'hc405761;
      28679: inst = 32'h8220000;
      28680: inst = 32'h10408000;
      28681: inst = 32'hc405762;
      28682: inst = 32'h8220000;
      28683: inst = 32'h10408000;
      28684: inst = 32'hc405763;
      28685: inst = 32'h8220000;
      28686: inst = 32'h10408000;
      28687: inst = 32'hc405764;
      28688: inst = 32'h8220000;
      28689: inst = 32'h10408000;
      28690: inst = 32'hc405765;
      28691: inst = 32'h8220000;
      28692: inst = 32'h10408000;
      28693: inst = 32'hc405766;
      28694: inst = 32'h8220000;
      28695: inst = 32'h10408000;
      28696: inst = 32'hc405767;
      28697: inst = 32'h8220000;
      28698: inst = 32'h10408000;
      28699: inst = 32'hc405768;
      28700: inst = 32'h8220000;
      28701: inst = 32'h10408000;
      28702: inst = 32'hc405769;
      28703: inst = 32'h8220000;
      28704: inst = 32'h10408000;
      28705: inst = 32'hc40576a;
      28706: inst = 32'h8220000;
      28707: inst = 32'h10408000;
      28708: inst = 32'hc40576b;
      28709: inst = 32'h8220000;
      28710: inst = 32'h10408000;
      28711: inst = 32'hc40576c;
      28712: inst = 32'h8220000;
      28713: inst = 32'h10408000;
      28714: inst = 32'hc40576d;
      28715: inst = 32'h8220000;
      28716: inst = 32'h10408000;
      28717: inst = 32'hc40576e;
      28718: inst = 32'h8220000;
      28719: inst = 32'h10408000;
      28720: inst = 32'hc40576f;
      28721: inst = 32'h8220000;
      28722: inst = 32'h10408000;
      28723: inst = 32'hc405770;
      28724: inst = 32'h8220000;
      28725: inst = 32'h10408000;
      28726: inst = 32'hc40577d;
      28727: inst = 32'h8220000;
      28728: inst = 32'h10408000;
      28729: inst = 32'hc40577e;
      28730: inst = 32'h8220000;
      28731: inst = 32'h10408000;
      28732: inst = 32'hc40577f;
      28733: inst = 32'h8220000;
      28734: inst = 32'h10408000;
      28735: inst = 32'hc405780;
      28736: inst = 32'h8220000;
      28737: inst = 32'h10408000;
      28738: inst = 32'hc405781;
      28739: inst = 32'h8220000;
      28740: inst = 32'h10408000;
      28741: inst = 32'hc405782;
      28742: inst = 32'h8220000;
      28743: inst = 32'h10408000;
      28744: inst = 32'hc405783;
      28745: inst = 32'h8220000;
      28746: inst = 32'h10408000;
      28747: inst = 32'hc405784;
      28748: inst = 32'h8220000;
      28749: inst = 32'h10408000;
      28750: inst = 32'hc405785;
      28751: inst = 32'h8220000;
      28752: inst = 32'h10408000;
      28753: inst = 32'hc405786;
      28754: inst = 32'h8220000;
      28755: inst = 32'h10408000;
      28756: inst = 32'hc405787;
      28757: inst = 32'h8220000;
      28758: inst = 32'h10408000;
      28759: inst = 32'hc405788;
      28760: inst = 32'h8220000;
      28761: inst = 32'h10408000;
      28762: inst = 32'hc405789;
      28763: inst = 32'h8220000;
      28764: inst = 32'h10408000;
      28765: inst = 32'hc40578a;
      28766: inst = 32'h8220000;
      28767: inst = 32'h10408000;
      28768: inst = 32'hc40578b;
      28769: inst = 32'h8220000;
      28770: inst = 32'h10408000;
      28771: inst = 32'hc40578c;
      28772: inst = 32'h8220000;
      28773: inst = 32'h10408000;
      28774: inst = 32'hc40578d;
      28775: inst = 32'h8220000;
      28776: inst = 32'h10408000;
      28777: inst = 32'hc40578e;
      28778: inst = 32'h8220000;
      28779: inst = 32'h10408000;
      28780: inst = 32'hc40578f;
      28781: inst = 32'h8220000;
      28782: inst = 32'h10408000;
      28783: inst = 32'hc405790;
      28784: inst = 32'h8220000;
      28785: inst = 32'h10408000;
      28786: inst = 32'hc405791;
      28787: inst = 32'h8220000;
      28788: inst = 32'h10408000;
      28789: inst = 32'hc405792;
      28790: inst = 32'h8220000;
      28791: inst = 32'h10408000;
      28792: inst = 32'hc405793;
      28793: inst = 32'h8220000;
      28794: inst = 32'h10408000;
      28795: inst = 32'hc405794;
      28796: inst = 32'h8220000;
      28797: inst = 32'h10408000;
      28798: inst = 32'hc405795;
      28799: inst = 32'h8220000;
      28800: inst = 32'h10408000;
      28801: inst = 32'hc405796;
      28802: inst = 32'h8220000;
      28803: inst = 32'h10408000;
      28804: inst = 32'hc405797;
      28805: inst = 32'h8220000;
      28806: inst = 32'h10408000;
      28807: inst = 32'hc405798;
      28808: inst = 32'h8220000;
      28809: inst = 32'h10408000;
      28810: inst = 32'hc405799;
      28811: inst = 32'h8220000;
      28812: inst = 32'h10408000;
      28813: inst = 32'hc40579a;
      28814: inst = 32'h8220000;
      28815: inst = 32'h10408000;
      28816: inst = 32'hc40579b;
      28817: inst = 32'h8220000;
      28818: inst = 32'h10408000;
      28819: inst = 32'hc40579c;
      28820: inst = 32'h8220000;
      28821: inst = 32'h10408000;
      28822: inst = 32'hc40579d;
      28823: inst = 32'h8220000;
      28824: inst = 32'h10408000;
      28825: inst = 32'hc40579e;
      28826: inst = 32'h8220000;
      28827: inst = 32'h10408000;
      28828: inst = 32'hc40579f;
      28829: inst = 32'h8220000;
      28830: inst = 32'h10408000;
      28831: inst = 32'hc4057a0;
      28832: inst = 32'h8220000;
      28833: inst = 32'h10408000;
      28834: inst = 32'hc4057a1;
      28835: inst = 32'h8220000;
      28836: inst = 32'h10408000;
      28837: inst = 32'hc4057a2;
      28838: inst = 32'h8220000;
      28839: inst = 32'h10408000;
      28840: inst = 32'hc4057a3;
      28841: inst = 32'h8220000;
      28842: inst = 32'h10408000;
      28843: inst = 32'hc4057a4;
      28844: inst = 32'h8220000;
      28845: inst = 32'h10408000;
      28846: inst = 32'hc4057a5;
      28847: inst = 32'h8220000;
      28848: inst = 32'h10408000;
      28849: inst = 32'hc4057a6;
      28850: inst = 32'h8220000;
      28851: inst = 32'h10408000;
      28852: inst = 32'hc4057a7;
      28853: inst = 32'h8220000;
      28854: inst = 32'h10408000;
      28855: inst = 32'hc4057a8;
      28856: inst = 32'h8220000;
      28857: inst = 32'h10408000;
      28858: inst = 32'hc4057a9;
      28859: inst = 32'h8220000;
      28860: inst = 32'h10408000;
      28861: inst = 32'hc4057aa;
      28862: inst = 32'h8220000;
      28863: inst = 32'h10408000;
      28864: inst = 32'hc4057ab;
      28865: inst = 32'h8220000;
      28866: inst = 32'h10408000;
      28867: inst = 32'hc4057ac;
      28868: inst = 32'h8220000;
      28869: inst = 32'h10408000;
      28870: inst = 32'hc4057ad;
      28871: inst = 32'h8220000;
      28872: inst = 32'h10408000;
      28873: inst = 32'hc4057ae;
      28874: inst = 32'h8220000;
      28875: inst = 32'h10408000;
      28876: inst = 32'hc4057af;
      28877: inst = 32'h8220000;
      28878: inst = 32'h10408000;
      28879: inst = 32'hc4057b0;
      28880: inst = 32'h8220000;
      28881: inst = 32'h10408000;
      28882: inst = 32'hc4057b1;
      28883: inst = 32'h8220000;
      28884: inst = 32'h10408000;
      28885: inst = 32'hc4057b2;
      28886: inst = 32'h8220000;
      28887: inst = 32'h10408000;
      28888: inst = 32'hc4057b3;
      28889: inst = 32'h8220000;
      28890: inst = 32'h10408000;
      28891: inst = 32'hc4057b4;
      28892: inst = 32'h8220000;
      28893: inst = 32'h10408000;
      28894: inst = 32'hc4057b5;
      28895: inst = 32'h8220000;
      28896: inst = 32'h10408000;
      28897: inst = 32'hc4057b6;
      28898: inst = 32'h8220000;
      28899: inst = 32'h10408000;
      28900: inst = 32'hc4057b7;
      28901: inst = 32'h8220000;
      28902: inst = 32'h10408000;
      28903: inst = 32'hc4057b8;
      28904: inst = 32'h8220000;
      28905: inst = 32'h10408000;
      28906: inst = 32'hc4057b9;
      28907: inst = 32'h8220000;
      28908: inst = 32'h10408000;
      28909: inst = 32'hc4057ba;
      28910: inst = 32'h8220000;
      28911: inst = 32'h10408000;
      28912: inst = 32'hc4057bb;
      28913: inst = 32'h8220000;
      28914: inst = 32'h10408000;
      28915: inst = 32'hc4057bc;
      28916: inst = 32'h8220000;
      28917: inst = 32'h10408000;
      28918: inst = 32'hc4057bd;
      28919: inst = 32'h8220000;
      28920: inst = 32'h10408000;
      28921: inst = 32'hc4057be;
      28922: inst = 32'h8220000;
      28923: inst = 32'h10408000;
      28924: inst = 32'hc4057c1;
      28925: inst = 32'h8220000;
      28926: inst = 32'h10408000;
      28927: inst = 32'hc4057c2;
      28928: inst = 32'h8220000;
      28929: inst = 32'h10408000;
      28930: inst = 32'hc4057c3;
      28931: inst = 32'h8220000;
      28932: inst = 32'h10408000;
      28933: inst = 32'hc4057c4;
      28934: inst = 32'h8220000;
      28935: inst = 32'h10408000;
      28936: inst = 32'hc4057c5;
      28937: inst = 32'h8220000;
      28938: inst = 32'h10408000;
      28939: inst = 32'hc4057c6;
      28940: inst = 32'h8220000;
      28941: inst = 32'h10408000;
      28942: inst = 32'hc4057c7;
      28943: inst = 32'h8220000;
      28944: inst = 32'h10408000;
      28945: inst = 32'hc4057c8;
      28946: inst = 32'h8220000;
      28947: inst = 32'h10408000;
      28948: inst = 32'hc4057c9;
      28949: inst = 32'h8220000;
      28950: inst = 32'h10408000;
      28951: inst = 32'hc4057ca;
      28952: inst = 32'h8220000;
      28953: inst = 32'h10408000;
      28954: inst = 32'hc4057cb;
      28955: inst = 32'h8220000;
      28956: inst = 32'h10408000;
      28957: inst = 32'hc4057cc;
      28958: inst = 32'h8220000;
      28959: inst = 32'h10408000;
      28960: inst = 32'hc4057cd;
      28961: inst = 32'h8220000;
      28962: inst = 32'h10408000;
      28963: inst = 32'hc4057ce;
      28964: inst = 32'h8220000;
      28965: inst = 32'h10408000;
      28966: inst = 32'hc4057cf;
      28967: inst = 32'h8220000;
      28968: inst = 32'h10408000;
      28969: inst = 32'hc4057d0;
      28970: inst = 32'h8220000;
      28971: inst = 32'h10408000;
      28972: inst = 32'hc4057dd;
      28973: inst = 32'h8220000;
      28974: inst = 32'h10408000;
      28975: inst = 32'hc4057de;
      28976: inst = 32'h8220000;
      28977: inst = 32'h10408000;
      28978: inst = 32'hc4057df;
      28979: inst = 32'h8220000;
      28980: inst = 32'hc20eeb6;
      28981: inst = 32'h10408000;
      28982: inst = 32'hc403fe3;
      28983: inst = 32'h8220000;
      28984: inst = 32'h10408000;
      28985: inst = 32'hc404043;
      28986: inst = 32'h8220000;
      28987: inst = 32'h10408000;
      28988: inst = 32'hc4040a3;
      28989: inst = 32'h8220000;
      28990: inst = 32'h10408000;
      28991: inst = 32'hc404103;
      28992: inst = 32'h8220000;
      28993: inst = 32'h10408000;
      28994: inst = 32'hc40410e;
      28995: inst = 32'h8220000;
      28996: inst = 32'h10408000;
      28997: inst = 32'hc40410f;
      28998: inst = 32'h8220000;
      28999: inst = 32'h10408000;
      29000: inst = 32'hc404110;
      29001: inst = 32'h8220000;
      29002: inst = 32'h10408000;
      29003: inst = 32'hc404111;
      29004: inst = 32'h8220000;
      29005: inst = 32'h10408000;
      29006: inst = 32'hc404112;
      29007: inst = 32'h8220000;
      29008: inst = 32'h10408000;
      29009: inst = 32'hc404115;
      29010: inst = 32'h8220000;
      29011: inst = 32'h10408000;
      29012: inst = 32'hc404118;
      29013: inst = 32'h8220000;
      29014: inst = 32'h10408000;
      29015: inst = 32'hc404119;
      29016: inst = 32'h8220000;
      29017: inst = 32'h10408000;
      29018: inst = 32'hc40411a;
      29019: inst = 32'h8220000;
      29020: inst = 32'h10408000;
      29021: inst = 32'hc40411b;
      29022: inst = 32'h8220000;
      29023: inst = 32'h10408000;
      29024: inst = 32'hc40411c;
      29025: inst = 32'h8220000;
      29026: inst = 32'h10408000;
      29027: inst = 32'hc40411d;
      29028: inst = 32'h8220000;
      29029: inst = 32'h10408000;
      29030: inst = 32'hc40411e;
      29031: inst = 32'h8220000;
      29032: inst = 32'h10408000;
      29033: inst = 32'hc40411f;
      29034: inst = 32'h8220000;
      29035: inst = 32'h10408000;
      29036: inst = 32'hc404120;
      29037: inst = 32'h8220000;
      29038: inst = 32'h10408000;
      29039: inst = 32'hc404121;
      29040: inst = 32'h8220000;
      29041: inst = 32'h10408000;
      29042: inst = 32'hc404122;
      29043: inst = 32'h8220000;
      29044: inst = 32'h10408000;
      29045: inst = 32'hc404123;
      29046: inst = 32'h8220000;
      29047: inst = 32'h10408000;
      29048: inst = 32'hc404124;
      29049: inst = 32'h8220000;
      29050: inst = 32'h10408000;
      29051: inst = 32'hc404125;
      29052: inst = 32'h8220000;
      29053: inst = 32'h10408000;
      29054: inst = 32'hc404126;
      29055: inst = 32'h8220000;
      29056: inst = 32'h10408000;
      29057: inst = 32'hc404127;
      29058: inst = 32'h8220000;
      29059: inst = 32'h10408000;
      29060: inst = 32'hc404128;
      29061: inst = 32'h8220000;
      29062: inst = 32'h10408000;
      29063: inst = 32'hc404129;
      29064: inst = 32'h8220000;
      29065: inst = 32'h10408000;
      29066: inst = 32'hc40412a;
      29067: inst = 32'h8220000;
      29068: inst = 32'h10408000;
      29069: inst = 32'hc40412b;
      29070: inst = 32'h8220000;
      29071: inst = 32'h10408000;
      29072: inst = 32'hc40412c;
      29073: inst = 32'h8220000;
      29074: inst = 32'h10408000;
      29075: inst = 32'hc40412d;
      29076: inst = 32'h8220000;
      29077: inst = 32'h10408000;
      29078: inst = 32'hc40412e;
      29079: inst = 32'h8220000;
      29080: inst = 32'h10408000;
      29081: inst = 32'hc40412f;
      29082: inst = 32'h8220000;
      29083: inst = 32'h10408000;
      29084: inst = 32'hc404130;
      29085: inst = 32'h8220000;
      29086: inst = 32'h10408000;
      29087: inst = 32'hc404131;
      29088: inst = 32'h8220000;
      29089: inst = 32'h10408000;
      29090: inst = 32'hc404132;
      29091: inst = 32'h8220000;
      29092: inst = 32'h10408000;
      29093: inst = 32'hc404133;
      29094: inst = 32'h8220000;
      29095: inst = 32'h10408000;
      29096: inst = 32'hc404134;
      29097: inst = 32'h8220000;
      29098: inst = 32'h10408000;
      29099: inst = 32'hc404135;
      29100: inst = 32'h8220000;
      29101: inst = 32'h10408000;
      29102: inst = 32'hc404136;
      29103: inst = 32'h8220000;
      29104: inst = 32'h10408000;
      29105: inst = 32'hc404137;
      29106: inst = 32'h8220000;
      29107: inst = 32'h10408000;
      29108: inst = 32'hc404138;
      29109: inst = 32'h8220000;
      29110: inst = 32'h10408000;
      29111: inst = 32'hc404139;
      29112: inst = 32'h8220000;
      29113: inst = 32'h10408000;
      29114: inst = 32'hc40413a;
      29115: inst = 32'h8220000;
      29116: inst = 32'h10408000;
      29117: inst = 32'hc40413b;
      29118: inst = 32'h8220000;
      29119: inst = 32'h10408000;
      29120: inst = 32'hc40413c;
      29121: inst = 32'h8220000;
      29122: inst = 32'h10408000;
      29123: inst = 32'hc40413d;
      29124: inst = 32'h8220000;
      29125: inst = 32'h10408000;
      29126: inst = 32'hc40413e;
      29127: inst = 32'h8220000;
      29128: inst = 32'h10408000;
      29129: inst = 32'hc40413f;
      29130: inst = 32'h8220000;
      29131: inst = 32'h10408000;
      29132: inst = 32'hc404140;
      29133: inst = 32'h8220000;
      29134: inst = 32'h10408000;
      29135: inst = 32'hc404141;
      29136: inst = 32'h8220000;
      29137: inst = 32'h10408000;
      29138: inst = 32'hc404142;
      29139: inst = 32'h8220000;
      29140: inst = 32'h10408000;
      29141: inst = 32'hc404143;
      29142: inst = 32'h8220000;
      29143: inst = 32'h10408000;
      29144: inst = 32'hc404144;
      29145: inst = 32'h8220000;
      29146: inst = 32'h10408000;
      29147: inst = 32'hc404145;
      29148: inst = 32'h8220000;
      29149: inst = 32'h10408000;
      29150: inst = 32'hc404146;
      29151: inst = 32'h8220000;
      29152: inst = 32'h10408000;
      29153: inst = 32'hc404147;
      29154: inst = 32'h8220000;
      29155: inst = 32'h10408000;
      29156: inst = 32'hc404148;
      29157: inst = 32'h8220000;
      29158: inst = 32'h10408000;
      29159: inst = 32'hc404149;
      29160: inst = 32'h8220000;
      29161: inst = 32'h10408000;
      29162: inst = 32'hc40414a;
      29163: inst = 32'h8220000;
      29164: inst = 32'h10408000;
      29165: inst = 32'hc40414b;
      29166: inst = 32'h8220000;
      29167: inst = 32'h10408000;
      29168: inst = 32'hc40414f;
      29169: inst = 32'h8220000;
      29170: inst = 32'h10408000;
      29171: inst = 32'hc404150;
      29172: inst = 32'h8220000;
      29173: inst = 32'h10408000;
      29174: inst = 32'hc404163;
      29175: inst = 32'h8220000;
      29176: inst = 32'h10408000;
      29177: inst = 32'hc40416e;
      29178: inst = 32'h8220000;
      29179: inst = 32'h10408000;
      29180: inst = 32'hc40416f;
      29181: inst = 32'h8220000;
      29182: inst = 32'h10408000;
      29183: inst = 32'hc404170;
      29184: inst = 32'h8220000;
      29185: inst = 32'h10408000;
      29186: inst = 32'hc404171;
      29187: inst = 32'h8220000;
      29188: inst = 32'h10408000;
      29189: inst = 32'hc404172;
      29190: inst = 32'h8220000;
      29191: inst = 32'h10408000;
      29192: inst = 32'hc404173;
      29193: inst = 32'h8220000;
      29194: inst = 32'h10408000;
      29195: inst = 32'hc404174;
      29196: inst = 32'h8220000;
      29197: inst = 32'h10408000;
      29198: inst = 32'hc404175;
      29199: inst = 32'h8220000;
      29200: inst = 32'h10408000;
      29201: inst = 32'hc404178;
      29202: inst = 32'h8220000;
      29203: inst = 32'h10408000;
      29204: inst = 32'hc404179;
      29205: inst = 32'h8220000;
      29206: inst = 32'h10408000;
      29207: inst = 32'hc40417a;
      29208: inst = 32'h8220000;
      29209: inst = 32'h10408000;
      29210: inst = 32'hc40417c;
      29211: inst = 32'h8220000;
      29212: inst = 32'h10408000;
      29213: inst = 32'hc40417d;
      29214: inst = 32'h8220000;
      29215: inst = 32'h10408000;
      29216: inst = 32'hc40417e;
      29217: inst = 32'h8220000;
      29218: inst = 32'h10408000;
      29219: inst = 32'hc40417f;
      29220: inst = 32'h8220000;
      29221: inst = 32'h10408000;
      29222: inst = 32'hc404180;
      29223: inst = 32'h8220000;
      29224: inst = 32'h10408000;
      29225: inst = 32'hc404181;
      29226: inst = 32'h8220000;
      29227: inst = 32'h10408000;
      29228: inst = 32'hc404182;
      29229: inst = 32'h8220000;
      29230: inst = 32'h10408000;
      29231: inst = 32'hc404183;
      29232: inst = 32'h8220000;
      29233: inst = 32'h10408000;
      29234: inst = 32'hc404184;
      29235: inst = 32'h8220000;
      29236: inst = 32'h10408000;
      29237: inst = 32'hc404185;
      29238: inst = 32'h8220000;
      29239: inst = 32'h10408000;
      29240: inst = 32'hc404186;
      29241: inst = 32'h8220000;
      29242: inst = 32'h10408000;
      29243: inst = 32'hc404187;
      29244: inst = 32'h8220000;
      29245: inst = 32'h10408000;
      29246: inst = 32'hc404188;
      29247: inst = 32'h8220000;
      29248: inst = 32'h10408000;
      29249: inst = 32'hc404189;
      29250: inst = 32'h8220000;
      29251: inst = 32'h10408000;
      29252: inst = 32'hc40418a;
      29253: inst = 32'h8220000;
      29254: inst = 32'h10408000;
      29255: inst = 32'hc40418b;
      29256: inst = 32'h8220000;
      29257: inst = 32'h10408000;
      29258: inst = 32'hc40418c;
      29259: inst = 32'h8220000;
      29260: inst = 32'h10408000;
      29261: inst = 32'hc40418d;
      29262: inst = 32'h8220000;
      29263: inst = 32'h10408000;
      29264: inst = 32'hc40418e;
      29265: inst = 32'h8220000;
      29266: inst = 32'h10408000;
      29267: inst = 32'hc40418f;
      29268: inst = 32'h8220000;
      29269: inst = 32'h10408000;
      29270: inst = 32'hc404190;
      29271: inst = 32'h8220000;
      29272: inst = 32'h10408000;
      29273: inst = 32'hc404191;
      29274: inst = 32'h8220000;
      29275: inst = 32'h10408000;
      29276: inst = 32'hc404192;
      29277: inst = 32'h8220000;
      29278: inst = 32'h10408000;
      29279: inst = 32'hc404193;
      29280: inst = 32'h8220000;
      29281: inst = 32'h10408000;
      29282: inst = 32'hc404194;
      29283: inst = 32'h8220000;
      29284: inst = 32'h10408000;
      29285: inst = 32'hc404195;
      29286: inst = 32'h8220000;
      29287: inst = 32'h10408000;
      29288: inst = 32'hc404196;
      29289: inst = 32'h8220000;
      29290: inst = 32'h10408000;
      29291: inst = 32'hc404197;
      29292: inst = 32'h8220000;
      29293: inst = 32'h10408000;
      29294: inst = 32'hc404198;
      29295: inst = 32'h8220000;
      29296: inst = 32'h10408000;
      29297: inst = 32'hc404199;
      29298: inst = 32'h8220000;
      29299: inst = 32'h10408000;
      29300: inst = 32'hc40419a;
      29301: inst = 32'h8220000;
      29302: inst = 32'h10408000;
      29303: inst = 32'hc40419b;
      29304: inst = 32'h8220000;
      29305: inst = 32'h10408000;
      29306: inst = 32'hc40419c;
      29307: inst = 32'h8220000;
      29308: inst = 32'h10408000;
      29309: inst = 32'hc40419d;
      29310: inst = 32'h8220000;
      29311: inst = 32'h10408000;
      29312: inst = 32'hc40419e;
      29313: inst = 32'h8220000;
      29314: inst = 32'h10408000;
      29315: inst = 32'hc40419f;
      29316: inst = 32'h8220000;
      29317: inst = 32'h10408000;
      29318: inst = 32'hc4041a0;
      29319: inst = 32'h8220000;
      29320: inst = 32'h10408000;
      29321: inst = 32'hc4041a1;
      29322: inst = 32'h8220000;
      29323: inst = 32'h10408000;
      29324: inst = 32'hc4041a2;
      29325: inst = 32'h8220000;
      29326: inst = 32'h10408000;
      29327: inst = 32'hc4041a3;
      29328: inst = 32'h8220000;
      29329: inst = 32'h10408000;
      29330: inst = 32'hc4041a4;
      29331: inst = 32'h8220000;
      29332: inst = 32'h10408000;
      29333: inst = 32'hc4041a5;
      29334: inst = 32'h8220000;
      29335: inst = 32'h10408000;
      29336: inst = 32'hc4041a6;
      29337: inst = 32'h8220000;
      29338: inst = 32'h10408000;
      29339: inst = 32'hc4041a7;
      29340: inst = 32'h8220000;
      29341: inst = 32'h10408000;
      29342: inst = 32'hc4041a8;
      29343: inst = 32'h8220000;
      29344: inst = 32'h10408000;
      29345: inst = 32'hc4041a9;
      29346: inst = 32'h8220000;
      29347: inst = 32'h10408000;
      29348: inst = 32'hc4041aa;
      29349: inst = 32'h8220000;
      29350: inst = 32'h10408000;
      29351: inst = 32'hc4041ab;
      29352: inst = 32'h8220000;
      29353: inst = 32'h10408000;
      29354: inst = 32'hc4041af;
      29355: inst = 32'h8220000;
      29356: inst = 32'h10408000;
      29357: inst = 32'hc4041b5;
      29358: inst = 32'h8220000;
      29359: inst = 32'h10408000;
      29360: inst = 32'hc4041c3;
      29361: inst = 32'h8220000;
      29362: inst = 32'h10408000;
      29363: inst = 32'hc4041cd;
      29364: inst = 32'h8220000;
      29365: inst = 32'h10408000;
      29366: inst = 32'hc4041ce;
      29367: inst = 32'h8220000;
      29368: inst = 32'h10408000;
      29369: inst = 32'hc4041cf;
      29370: inst = 32'h8220000;
      29371: inst = 32'h10408000;
      29372: inst = 32'hc4041d2;
      29373: inst = 32'h8220000;
      29374: inst = 32'h10408000;
      29375: inst = 32'hc4041d3;
      29376: inst = 32'h8220000;
      29377: inst = 32'h10408000;
      29378: inst = 32'hc4041d4;
      29379: inst = 32'h8220000;
      29380: inst = 32'h10408000;
      29381: inst = 32'hc4041d5;
      29382: inst = 32'h8220000;
      29383: inst = 32'h10408000;
      29384: inst = 32'hc4041d9;
      29385: inst = 32'h8220000;
      29386: inst = 32'h10408000;
      29387: inst = 32'hc4041da;
      29388: inst = 32'h8220000;
      29389: inst = 32'h10408000;
      29390: inst = 32'hc4041dd;
      29391: inst = 32'h8220000;
      29392: inst = 32'h10408000;
      29393: inst = 32'hc4041de;
      29394: inst = 32'h8220000;
      29395: inst = 32'h10408000;
      29396: inst = 32'hc4041df;
      29397: inst = 32'h8220000;
      29398: inst = 32'h10408000;
      29399: inst = 32'hc4041e0;
      29400: inst = 32'h8220000;
      29401: inst = 32'h10408000;
      29402: inst = 32'hc4041e1;
      29403: inst = 32'h8220000;
      29404: inst = 32'h10408000;
      29405: inst = 32'hc4041e2;
      29406: inst = 32'h8220000;
      29407: inst = 32'h10408000;
      29408: inst = 32'hc4041e3;
      29409: inst = 32'h8220000;
      29410: inst = 32'h10408000;
      29411: inst = 32'hc4041e4;
      29412: inst = 32'h8220000;
      29413: inst = 32'h10408000;
      29414: inst = 32'hc4041e5;
      29415: inst = 32'h8220000;
      29416: inst = 32'h10408000;
      29417: inst = 32'hc4041e6;
      29418: inst = 32'h8220000;
      29419: inst = 32'h10408000;
      29420: inst = 32'hc4041e7;
      29421: inst = 32'h8220000;
      29422: inst = 32'h10408000;
      29423: inst = 32'hc4041e8;
      29424: inst = 32'h8220000;
      29425: inst = 32'h10408000;
      29426: inst = 32'hc4041e9;
      29427: inst = 32'h8220000;
      29428: inst = 32'h10408000;
      29429: inst = 32'hc4041ea;
      29430: inst = 32'h8220000;
      29431: inst = 32'h10408000;
      29432: inst = 32'hc4041eb;
      29433: inst = 32'h8220000;
      29434: inst = 32'h10408000;
      29435: inst = 32'hc4041ec;
      29436: inst = 32'h8220000;
      29437: inst = 32'h10408000;
      29438: inst = 32'hc4041ed;
      29439: inst = 32'h8220000;
      29440: inst = 32'h10408000;
      29441: inst = 32'hc4041ee;
      29442: inst = 32'h8220000;
      29443: inst = 32'h10408000;
      29444: inst = 32'hc4041ef;
      29445: inst = 32'h8220000;
      29446: inst = 32'h10408000;
      29447: inst = 32'hc4041f0;
      29448: inst = 32'h8220000;
      29449: inst = 32'h10408000;
      29450: inst = 32'hc4041f1;
      29451: inst = 32'h8220000;
      29452: inst = 32'h10408000;
      29453: inst = 32'hc4041f2;
      29454: inst = 32'h8220000;
      29455: inst = 32'h10408000;
      29456: inst = 32'hc4041f3;
      29457: inst = 32'h8220000;
      29458: inst = 32'h10408000;
      29459: inst = 32'hc4041f4;
      29460: inst = 32'h8220000;
      29461: inst = 32'h10408000;
      29462: inst = 32'hc4041f5;
      29463: inst = 32'h8220000;
      29464: inst = 32'h10408000;
      29465: inst = 32'hc4041f6;
      29466: inst = 32'h8220000;
      29467: inst = 32'h10408000;
      29468: inst = 32'hc4041f7;
      29469: inst = 32'h8220000;
      29470: inst = 32'h10408000;
      29471: inst = 32'hc4041f8;
      29472: inst = 32'h8220000;
      29473: inst = 32'h10408000;
      29474: inst = 32'hc4041f9;
      29475: inst = 32'h8220000;
      29476: inst = 32'h10408000;
      29477: inst = 32'hc4041fa;
      29478: inst = 32'h8220000;
      29479: inst = 32'h10408000;
      29480: inst = 32'hc4041fb;
      29481: inst = 32'h8220000;
      29482: inst = 32'h10408000;
      29483: inst = 32'hc4041fc;
      29484: inst = 32'h8220000;
      29485: inst = 32'h10408000;
      29486: inst = 32'hc4041fd;
      29487: inst = 32'h8220000;
      29488: inst = 32'h10408000;
      29489: inst = 32'hc4041fe;
      29490: inst = 32'h8220000;
      29491: inst = 32'h10408000;
      29492: inst = 32'hc4041ff;
      29493: inst = 32'h8220000;
      29494: inst = 32'h10408000;
      29495: inst = 32'hc404200;
      29496: inst = 32'h8220000;
      29497: inst = 32'h10408000;
      29498: inst = 32'hc404201;
      29499: inst = 32'h8220000;
      29500: inst = 32'h10408000;
      29501: inst = 32'hc404202;
      29502: inst = 32'h8220000;
      29503: inst = 32'h10408000;
      29504: inst = 32'hc404203;
      29505: inst = 32'h8220000;
      29506: inst = 32'h10408000;
      29507: inst = 32'hc404204;
      29508: inst = 32'h8220000;
      29509: inst = 32'h10408000;
      29510: inst = 32'hc404205;
      29511: inst = 32'h8220000;
      29512: inst = 32'h10408000;
      29513: inst = 32'hc404206;
      29514: inst = 32'h8220000;
      29515: inst = 32'h10408000;
      29516: inst = 32'hc404207;
      29517: inst = 32'h8220000;
      29518: inst = 32'h10408000;
      29519: inst = 32'hc404208;
      29520: inst = 32'h8220000;
      29521: inst = 32'h10408000;
      29522: inst = 32'hc404209;
      29523: inst = 32'h8220000;
      29524: inst = 32'h10408000;
      29525: inst = 32'hc40420a;
      29526: inst = 32'h8220000;
      29527: inst = 32'h10408000;
      29528: inst = 32'hc40420b;
      29529: inst = 32'h8220000;
      29530: inst = 32'h10408000;
      29531: inst = 32'hc40420f;
      29532: inst = 32'h8220000;
      29533: inst = 32'h10408000;
      29534: inst = 32'hc404214;
      29535: inst = 32'h8220000;
      29536: inst = 32'h10408000;
      29537: inst = 32'hc404223;
      29538: inst = 32'h8220000;
      29539: inst = 32'h10408000;
      29540: inst = 32'hc40422d;
      29541: inst = 32'h8220000;
      29542: inst = 32'h10408000;
      29543: inst = 32'hc40422e;
      29544: inst = 32'h8220000;
      29545: inst = 32'h10408000;
      29546: inst = 32'hc404232;
      29547: inst = 32'h8220000;
      29548: inst = 32'h10408000;
      29549: inst = 32'hc404233;
      29550: inst = 32'h8220000;
      29551: inst = 32'h10408000;
      29552: inst = 32'hc404234;
      29553: inst = 32'h8220000;
      29554: inst = 32'h10408000;
      29555: inst = 32'hc404235;
      29556: inst = 32'h8220000;
      29557: inst = 32'h10408000;
      29558: inst = 32'hc404236;
      29559: inst = 32'h8220000;
      29560: inst = 32'h10408000;
      29561: inst = 32'hc404237;
      29562: inst = 32'h8220000;
      29563: inst = 32'h10408000;
      29564: inst = 32'hc404238;
      29565: inst = 32'h8220000;
      29566: inst = 32'h10408000;
      29567: inst = 32'hc404239;
      29568: inst = 32'h8220000;
      29569: inst = 32'h10408000;
      29570: inst = 32'hc40423a;
      29571: inst = 32'h8220000;
      29572: inst = 32'h10408000;
      29573: inst = 32'hc40423d;
      29574: inst = 32'h8220000;
      29575: inst = 32'h10408000;
      29576: inst = 32'hc40423e;
      29577: inst = 32'h8220000;
      29578: inst = 32'h10408000;
      29579: inst = 32'hc40423f;
      29580: inst = 32'h8220000;
      29581: inst = 32'h10408000;
      29582: inst = 32'hc404240;
      29583: inst = 32'h8220000;
      29584: inst = 32'h10408000;
      29585: inst = 32'hc404241;
      29586: inst = 32'h8220000;
      29587: inst = 32'h10408000;
      29588: inst = 32'hc404242;
      29589: inst = 32'h8220000;
      29590: inst = 32'h10408000;
      29591: inst = 32'hc404243;
      29592: inst = 32'h8220000;
      29593: inst = 32'h10408000;
      29594: inst = 32'hc404244;
      29595: inst = 32'h8220000;
      29596: inst = 32'h10408000;
      29597: inst = 32'hc404245;
      29598: inst = 32'h8220000;
      29599: inst = 32'h10408000;
      29600: inst = 32'hc404246;
      29601: inst = 32'h8220000;
      29602: inst = 32'h10408000;
      29603: inst = 32'hc404247;
      29604: inst = 32'h8220000;
      29605: inst = 32'h10408000;
      29606: inst = 32'hc404248;
      29607: inst = 32'h8220000;
      29608: inst = 32'h10408000;
      29609: inst = 32'hc404249;
      29610: inst = 32'h8220000;
      29611: inst = 32'h10408000;
      29612: inst = 32'hc40424a;
      29613: inst = 32'h8220000;
      29614: inst = 32'h10408000;
      29615: inst = 32'hc40424b;
      29616: inst = 32'h8220000;
      29617: inst = 32'h10408000;
      29618: inst = 32'hc40424c;
      29619: inst = 32'h8220000;
      29620: inst = 32'h10408000;
      29621: inst = 32'hc40424d;
      29622: inst = 32'h8220000;
      29623: inst = 32'h10408000;
      29624: inst = 32'hc40424e;
      29625: inst = 32'h8220000;
      29626: inst = 32'h10408000;
      29627: inst = 32'hc40424f;
      29628: inst = 32'h8220000;
      29629: inst = 32'h10408000;
      29630: inst = 32'hc404250;
      29631: inst = 32'h8220000;
      29632: inst = 32'h10408000;
      29633: inst = 32'hc404251;
      29634: inst = 32'h8220000;
      29635: inst = 32'h10408000;
      29636: inst = 32'hc404252;
      29637: inst = 32'h8220000;
      29638: inst = 32'h10408000;
      29639: inst = 32'hc404253;
      29640: inst = 32'h8220000;
      29641: inst = 32'h10408000;
      29642: inst = 32'hc404254;
      29643: inst = 32'h8220000;
      29644: inst = 32'h10408000;
      29645: inst = 32'hc404255;
      29646: inst = 32'h8220000;
      29647: inst = 32'h10408000;
      29648: inst = 32'hc404256;
      29649: inst = 32'h8220000;
      29650: inst = 32'h10408000;
      29651: inst = 32'hc404257;
      29652: inst = 32'h8220000;
      29653: inst = 32'h10408000;
      29654: inst = 32'hc404258;
      29655: inst = 32'h8220000;
      29656: inst = 32'h10408000;
      29657: inst = 32'hc404259;
      29658: inst = 32'h8220000;
      29659: inst = 32'h10408000;
      29660: inst = 32'hc40425a;
      29661: inst = 32'h8220000;
      29662: inst = 32'h10408000;
      29663: inst = 32'hc40425b;
      29664: inst = 32'h8220000;
      29665: inst = 32'h10408000;
      29666: inst = 32'hc40425c;
      29667: inst = 32'h8220000;
      29668: inst = 32'h10408000;
      29669: inst = 32'hc40425d;
      29670: inst = 32'h8220000;
      29671: inst = 32'h10408000;
      29672: inst = 32'hc40425e;
      29673: inst = 32'h8220000;
      29674: inst = 32'h10408000;
      29675: inst = 32'hc40425f;
      29676: inst = 32'h8220000;
      29677: inst = 32'h10408000;
      29678: inst = 32'hc404260;
      29679: inst = 32'h8220000;
      29680: inst = 32'h10408000;
      29681: inst = 32'hc404261;
      29682: inst = 32'h8220000;
      29683: inst = 32'h10408000;
      29684: inst = 32'hc404262;
      29685: inst = 32'h8220000;
      29686: inst = 32'h10408000;
      29687: inst = 32'hc404263;
      29688: inst = 32'h8220000;
      29689: inst = 32'h10408000;
      29690: inst = 32'hc404264;
      29691: inst = 32'h8220000;
      29692: inst = 32'h10408000;
      29693: inst = 32'hc404265;
      29694: inst = 32'h8220000;
      29695: inst = 32'h10408000;
      29696: inst = 32'hc404266;
      29697: inst = 32'h8220000;
      29698: inst = 32'h10408000;
      29699: inst = 32'hc404267;
      29700: inst = 32'h8220000;
      29701: inst = 32'h10408000;
      29702: inst = 32'hc404268;
      29703: inst = 32'h8220000;
      29704: inst = 32'h10408000;
      29705: inst = 32'hc404269;
      29706: inst = 32'h8220000;
      29707: inst = 32'h10408000;
      29708: inst = 32'hc40426a;
      29709: inst = 32'h8220000;
      29710: inst = 32'h10408000;
      29711: inst = 32'hc40426b;
      29712: inst = 32'h8220000;
      29713: inst = 32'h10408000;
      29714: inst = 32'hc40426f;
      29715: inst = 32'h8220000;
      29716: inst = 32'h10408000;
      29717: inst = 32'hc404283;
      29718: inst = 32'h8220000;
      29719: inst = 32'h10408000;
      29720: inst = 32'hc40428d;
      29721: inst = 32'h8220000;
      29722: inst = 32'h10408000;
      29723: inst = 32'hc40428e;
      29724: inst = 32'h8220000;
      29725: inst = 32'h10408000;
      29726: inst = 32'hc404291;
      29727: inst = 32'h8220000;
      29728: inst = 32'h10408000;
      29729: inst = 32'hc404292;
      29730: inst = 32'h8220000;
      29731: inst = 32'h10408000;
      29732: inst = 32'hc404293;
      29733: inst = 32'h8220000;
      29734: inst = 32'h10408000;
      29735: inst = 32'hc404294;
      29736: inst = 32'h8220000;
      29737: inst = 32'h10408000;
      29738: inst = 32'hc404295;
      29739: inst = 32'h8220000;
      29740: inst = 32'h10408000;
      29741: inst = 32'hc404296;
      29742: inst = 32'h8220000;
      29743: inst = 32'h10408000;
      29744: inst = 32'hc404297;
      29745: inst = 32'h8220000;
      29746: inst = 32'h10408000;
      29747: inst = 32'hc404298;
      29748: inst = 32'h8220000;
      29749: inst = 32'h10408000;
      29750: inst = 32'hc404299;
      29751: inst = 32'h8220000;
      29752: inst = 32'h10408000;
      29753: inst = 32'hc40429a;
      29754: inst = 32'h8220000;
      29755: inst = 32'h10408000;
      29756: inst = 32'hc40429d;
      29757: inst = 32'h8220000;
      29758: inst = 32'h10408000;
      29759: inst = 32'hc40429e;
      29760: inst = 32'h8220000;
      29761: inst = 32'h10408000;
      29762: inst = 32'hc40429f;
      29763: inst = 32'h8220000;
      29764: inst = 32'h10408000;
      29765: inst = 32'hc4042a0;
      29766: inst = 32'h8220000;
      29767: inst = 32'h10408000;
      29768: inst = 32'hc4042a1;
      29769: inst = 32'h8220000;
      29770: inst = 32'h10408000;
      29771: inst = 32'hc4042a2;
      29772: inst = 32'h8220000;
      29773: inst = 32'h10408000;
      29774: inst = 32'hc4042a3;
      29775: inst = 32'h8220000;
      29776: inst = 32'h10408000;
      29777: inst = 32'hc4042a4;
      29778: inst = 32'h8220000;
      29779: inst = 32'h10408000;
      29780: inst = 32'hc4042a5;
      29781: inst = 32'h8220000;
      29782: inst = 32'h10408000;
      29783: inst = 32'hc4042a6;
      29784: inst = 32'h8220000;
      29785: inst = 32'h10408000;
      29786: inst = 32'hc4042a7;
      29787: inst = 32'h8220000;
      29788: inst = 32'h10408000;
      29789: inst = 32'hc4042a8;
      29790: inst = 32'h8220000;
      29791: inst = 32'h10408000;
      29792: inst = 32'hc4042a9;
      29793: inst = 32'h8220000;
      29794: inst = 32'h10408000;
      29795: inst = 32'hc4042aa;
      29796: inst = 32'h8220000;
      29797: inst = 32'h10408000;
      29798: inst = 32'hc4042ab;
      29799: inst = 32'h8220000;
      29800: inst = 32'h10408000;
      29801: inst = 32'hc4042ac;
      29802: inst = 32'h8220000;
      29803: inst = 32'h10408000;
      29804: inst = 32'hc4042ad;
      29805: inst = 32'h8220000;
      29806: inst = 32'h10408000;
      29807: inst = 32'hc4042ae;
      29808: inst = 32'h8220000;
      29809: inst = 32'h10408000;
      29810: inst = 32'hc4042af;
      29811: inst = 32'h8220000;
      29812: inst = 32'h10408000;
      29813: inst = 32'hc4042b0;
      29814: inst = 32'h8220000;
      29815: inst = 32'h10408000;
      29816: inst = 32'hc4042b1;
      29817: inst = 32'h8220000;
      29818: inst = 32'h10408000;
      29819: inst = 32'hc4042b2;
      29820: inst = 32'h8220000;
      29821: inst = 32'h10408000;
      29822: inst = 32'hc4042b3;
      29823: inst = 32'h8220000;
      29824: inst = 32'h10408000;
      29825: inst = 32'hc4042b4;
      29826: inst = 32'h8220000;
      29827: inst = 32'h10408000;
      29828: inst = 32'hc4042b5;
      29829: inst = 32'h8220000;
      29830: inst = 32'h10408000;
      29831: inst = 32'hc4042b6;
      29832: inst = 32'h8220000;
      29833: inst = 32'h10408000;
      29834: inst = 32'hc4042b7;
      29835: inst = 32'h8220000;
      29836: inst = 32'h10408000;
      29837: inst = 32'hc4042b8;
      29838: inst = 32'h8220000;
      29839: inst = 32'h10408000;
      29840: inst = 32'hc4042b9;
      29841: inst = 32'h8220000;
      29842: inst = 32'h10408000;
      29843: inst = 32'hc4042ba;
      29844: inst = 32'h8220000;
      29845: inst = 32'h10408000;
      29846: inst = 32'hc4042bb;
      29847: inst = 32'h8220000;
      29848: inst = 32'h10408000;
      29849: inst = 32'hc4042bc;
      29850: inst = 32'h8220000;
      29851: inst = 32'h10408000;
      29852: inst = 32'hc4042bd;
      29853: inst = 32'h8220000;
      29854: inst = 32'h10408000;
      29855: inst = 32'hc4042be;
      29856: inst = 32'h8220000;
      29857: inst = 32'h10408000;
      29858: inst = 32'hc4042bf;
      29859: inst = 32'h8220000;
      29860: inst = 32'h10408000;
      29861: inst = 32'hc4042c0;
      29862: inst = 32'h8220000;
      29863: inst = 32'h10408000;
      29864: inst = 32'hc4042c1;
      29865: inst = 32'h8220000;
      29866: inst = 32'h10408000;
      29867: inst = 32'hc4042c2;
      29868: inst = 32'h8220000;
      29869: inst = 32'h10408000;
      29870: inst = 32'hc4042c3;
      29871: inst = 32'h8220000;
      29872: inst = 32'h10408000;
      29873: inst = 32'hc4042c4;
      29874: inst = 32'h8220000;
      29875: inst = 32'h10408000;
      29876: inst = 32'hc4042c5;
      29877: inst = 32'h8220000;
      29878: inst = 32'h10408000;
      29879: inst = 32'hc4042c6;
      29880: inst = 32'h8220000;
      29881: inst = 32'h10408000;
      29882: inst = 32'hc4042c7;
      29883: inst = 32'h8220000;
      29884: inst = 32'h10408000;
      29885: inst = 32'hc4042c8;
      29886: inst = 32'h8220000;
      29887: inst = 32'h10408000;
      29888: inst = 32'hc4042c9;
      29889: inst = 32'h8220000;
      29890: inst = 32'h10408000;
      29891: inst = 32'hc4042ca;
      29892: inst = 32'h8220000;
      29893: inst = 32'h10408000;
      29894: inst = 32'hc4042cb;
      29895: inst = 32'h8220000;
      29896: inst = 32'h10408000;
      29897: inst = 32'hc4042cf;
      29898: inst = 32'h8220000;
      29899: inst = 32'h10408000;
      29900: inst = 32'hc4042d3;
      29901: inst = 32'h8220000;
      29902: inst = 32'h10408000;
      29903: inst = 32'hc4042da;
      29904: inst = 32'h8220000;
      29905: inst = 32'h10408000;
      29906: inst = 32'hc4042db;
      29907: inst = 32'h8220000;
      29908: inst = 32'h10408000;
      29909: inst = 32'hc4042e3;
      29910: inst = 32'h8220000;
      29911: inst = 32'h10408000;
      29912: inst = 32'hc4042ed;
      29913: inst = 32'h8220000;
      29914: inst = 32'h10408000;
      29915: inst = 32'hc4042ee;
      29916: inst = 32'h8220000;
      29917: inst = 32'h10408000;
      29918: inst = 32'hc4042ef;
      29919: inst = 32'h8220000;
      29920: inst = 32'h10408000;
      29921: inst = 32'hc4042f0;
      29922: inst = 32'h8220000;
      29923: inst = 32'h10408000;
      29924: inst = 32'hc4042f1;
      29925: inst = 32'h8220000;
      29926: inst = 32'h10408000;
      29927: inst = 32'hc4042f2;
      29928: inst = 32'h8220000;
      29929: inst = 32'h10408000;
      29930: inst = 32'hc4042f3;
      29931: inst = 32'h8220000;
      29932: inst = 32'h10408000;
      29933: inst = 32'hc4042f4;
      29934: inst = 32'h8220000;
      29935: inst = 32'h10408000;
      29936: inst = 32'hc4042f5;
      29937: inst = 32'h8220000;
      29938: inst = 32'h10408000;
      29939: inst = 32'hc4042f6;
      29940: inst = 32'h8220000;
      29941: inst = 32'h10408000;
      29942: inst = 32'hc4042f7;
      29943: inst = 32'h8220000;
      29944: inst = 32'h10408000;
      29945: inst = 32'hc4042f8;
      29946: inst = 32'h8220000;
      29947: inst = 32'h10408000;
      29948: inst = 32'hc4042f9;
      29949: inst = 32'h8220000;
      29950: inst = 32'h10408000;
      29951: inst = 32'hc4042fa;
      29952: inst = 32'h8220000;
      29953: inst = 32'h10408000;
      29954: inst = 32'hc4042fb;
      29955: inst = 32'h8220000;
      29956: inst = 32'h10408000;
      29957: inst = 32'hc4042fc;
      29958: inst = 32'h8220000;
      29959: inst = 32'h10408000;
      29960: inst = 32'hc4042fd;
      29961: inst = 32'h8220000;
      29962: inst = 32'h10408000;
      29963: inst = 32'hc4042fe;
      29964: inst = 32'h8220000;
      29965: inst = 32'h10408000;
      29966: inst = 32'hc4042ff;
      29967: inst = 32'h8220000;
      29968: inst = 32'h10408000;
      29969: inst = 32'hc404300;
      29970: inst = 32'h8220000;
      29971: inst = 32'h10408000;
      29972: inst = 32'hc404301;
      29973: inst = 32'h8220000;
      29974: inst = 32'h10408000;
      29975: inst = 32'hc404302;
      29976: inst = 32'h8220000;
      29977: inst = 32'h10408000;
      29978: inst = 32'hc404303;
      29979: inst = 32'h8220000;
      29980: inst = 32'h10408000;
      29981: inst = 32'hc404304;
      29982: inst = 32'h8220000;
      29983: inst = 32'h10408000;
      29984: inst = 32'hc404305;
      29985: inst = 32'h8220000;
      29986: inst = 32'h10408000;
      29987: inst = 32'hc404306;
      29988: inst = 32'h8220000;
      29989: inst = 32'h10408000;
      29990: inst = 32'hc404307;
      29991: inst = 32'h8220000;
      29992: inst = 32'h10408000;
      29993: inst = 32'hc404308;
      29994: inst = 32'h8220000;
      29995: inst = 32'h10408000;
      29996: inst = 32'hc404309;
      29997: inst = 32'h8220000;
      29998: inst = 32'h10408000;
      29999: inst = 32'hc40430a;
      30000: inst = 32'h8220000;
      30001: inst = 32'h10408000;
      30002: inst = 32'hc40430b;
      30003: inst = 32'h8220000;
      30004: inst = 32'h10408000;
      30005: inst = 32'hc40430c;
      30006: inst = 32'h8220000;
      30007: inst = 32'h10408000;
      30008: inst = 32'hc40430d;
      30009: inst = 32'h8220000;
      30010: inst = 32'h10408000;
      30011: inst = 32'hc40430e;
      30012: inst = 32'h8220000;
      30013: inst = 32'h10408000;
      30014: inst = 32'hc40430f;
      30015: inst = 32'h8220000;
      30016: inst = 32'h10408000;
      30017: inst = 32'hc404310;
      30018: inst = 32'h8220000;
      30019: inst = 32'h10408000;
      30020: inst = 32'hc404311;
      30021: inst = 32'h8220000;
      30022: inst = 32'h10408000;
      30023: inst = 32'hc404312;
      30024: inst = 32'h8220000;
      30025: inst = 32'h10408000;
      30026: inst = 32'hc404313;
      30027: inst = 32'h8220000;
      30028: inst = 32'h10408000;
      30029: inst = 32'hc404314;
      30030: inst = 32'h8220000;
      30031: inst = 32'h10408000;
      30032: inst = 32'hc404315;
      30033: inst = 32'h8220000;
      30034: inst = 32'h10408000;
      30035: inst = 32'hc404316;
      30036: inst = 32'h8220000;
      30037: inst = 32'h10408000;
      30038: inst = 32'hc404317;
      30039: inst = 32'h8220000;
      30040: inst = 32'h10408000;
      30041: inst = 32'hc404318;
      30042: inst = 32'h8220000;
      30043: inst = 32'h10408000;
      30044: inst = 32'hc404319;
      30045: inst = 32'h8220000;
      30046: inst = 32'h10408000;
      30047: inst = 32'hc40431a;
      30048: inst = 32'h8220000;
      30049: inst = 32'h10408000;
      30050: inst = 32'hc40431b;
      30051: inst = 32'h8220000;
      30052: inst = 32'h10408000;
      30053: inst = 32'hc40431c;
      30054: inst = 32'h8220000;
      30055: inst = 32'h10408000;
      30056: inst = 32'hc40431d;
      30057: inst = 32'h8220000;
      30058: inst = 32'h10408000;
      30059: inst = 32'hc40431e;
      30060: inst = 32'h8220000;
      30061: inst = 32'h10408000;
      30062: inst = 32'hc40431f;
      30063: inst = 32'h8220000;
      30064: inst = 32'h10408000;
      30065: inst = 32'hc404320;
      30066: inst = 32'h8220000;
      30067: inst = 32'h10408000;
      30068: inst = 32'hc404321;
      30069: inst = 32'h8220000;
      30070: inst = 32'h10408000;
      30071: inst = 32'hc404322;
      30072: inst = 32'h8220000;
      30073: inst = 32'h10408000;
      30074: inst = 32'hc404323;
      30075: inst = 32'h8220000;
      30076: inst = 32'h10408000;
      30077: inst = 32'hc404324;
      30078: inst = 32'h8220000;
      30079: inst = 32'h10408000;
      30080: inst = 32'hc404325;
      30081: inst = 32'h8220000;
      30082: inst = 32'h10408000;
      30083: inst = 32'hc404326;
      30084: inst = 32'h8220000;
      30085: inst = 32'h10408000;
      30086: inst = 32'hc404327;
      30087: inst = 32'h8220000;
      30088: inst = 32'h10408000;
      30089: inst = 32'hc404328;
      30090: inst = 32'h8220000;
      30091: inst = 32'h10408000;
      30092: inst = 32'hc404329;
      30093: inst = 32'h8220000;
      30094: inst = 32'h10408000;
      30095: inst = 32'hc40432a;
      30096: inst = 32'h8220000;
      30097: inst = 32'h10408000;
      30098: inst = 32'hc40432b;
      30099: inst = 32'h8220000;
      30100: inst = 32'h10408000;
      30101: inst = 32'hc40432f;
      30102: inst = 32'h8220000;
      30103: inst = 32'h10408000;
      30104: inst = 32'hc404330;
      30105: inst = 32'h8220000;
      30106: inst = 32'h10408000;
      30107: inst = 32'hc404333;
      30108: inst = 32'h8220000;
      30109: inst = 32'h10408000;
      30110: inst = 32'hc404334;
      30111: inst = 32'h8220000;
      30112: inst = 32'h10408000;
      30113: inst = 32'hc404343;
      30114: inst = 32'h8220000;
      30115: inst = 32'h10408000;
      30116: inst = 32'hc40434d;
      30117: inst = 32'h8220000;
      30118: inst = 32'h10408000;
      30119: inst = 32'hc40434e;
      30120: inst = 32'h8220000;
      30121: inst = 32'h10408000;
      30122: inst = 32'hc40434f;
      30123: inst = 32'h8220000;
      30124: inst = 32'h10408000;
      30125: inst = 32'hc404350;
      30126: inst = 32'h8220000;
      30127: inst = 32'h10408000;
      30128: inst = 32'hc404351;
      30129: inst = 32'h8220000;
      30130: inst = 32'h10408000;
      30131: inst = 32'hc404352;
      30132: inst = 32'h8220000;
      30133: inst = 32'h10408000;
      30134: inst = 32'hc404353;
      30135: inst = 32'h8220000;
      30136: inst = 32'h10408000;
      30137: inst = 32'hc404354;
      30138: inst = 32'h8220000;
      30139: inst = 32'h10408000;
      30140: inst = 32'hc404355;
      30141: inst = 32'h8220000;
      30142: inst = 32'h10408000;
      30143: inst = 32'hc404356;
      30144: inst = 32'h8220000;
      30145: inst = 32'h10408000;
      30146: inst = 32'hc404357;
      30147: inst = 32'h8220000;
      30148: inst = 32'h10408000;
      30149: inst = 32'hc404358;
      30150: inst = 32'h8220000;
      30151: inst = 32'h10408000;
      30152: inst = 32'hc404359;
      30153: inst = 32'h8220000;
      30154: inst = 32'h10408000;
      30155: inst = 32'hc40435a;
      30156: inst = 32'h8220000;
      30157: inst = 32'h10408000;
      30158: inst = 32'hc40435b;
      30159: inst = 32'h8220000;
      30160: inst = 32'h10408000;
      30161: inst = 32'hc40435c;
      30162: inst = 32'h8220000;
      30163: inst = 32'h10408000;
      30164: inst = 32'hc40435d;
      30165: inst = 32'h8220000;
      30166: inst = 32'h10408000;
      30167: inst = 32'hc40435e;
      30168: inst = 32'h8220000;
      30169: inst = 32'h10408000;
      30170: inst = 32'hc40435f;
      30171: inst = 32'h8220000;
      30172: inst = 32'h10408000;
      30173: inst = 32'hc404360;
      30174: inst = 32'h8220000;
      30175: inst = 32'h10408000;
      30176: inst = 32'hc404361;
      30177: inst = 32'h8220000;
      30178: inst = 32'h10408000;
      30179: inst = 32'hc404362;
      30180: inst = 32'h8220000;
      30181: inst = 32'h10408000;
      30182: inst = 32'hc404363;
      30183: inst = 32'h8220000;
      30184: inst = 32'h10408000;
      30185: inst = 32'hc404364;
      30186: inst = 32'h8220000;
      30187: inst = 32'h10408000;
      30188: inst = 32'hc404365;
      30189: inst = 32'h8220000;
      30190: inst = 32'h10408000;
      30191: inst = 32'hc404366;
      30192: inst = 32'h8220000;
      30193: inst = 32'h10408000;
      30194: inst = 32'hc404367;
      30195: inst = 32'h8220000;
      30196: inst = 32'h10408000;
      30197: inst = 32'hc404368;
      30198: inst = 32'h8220000;
      30199: inst = 32'h10408000;
      30200: inst = 32'hc404369;
      30201: inst = 32'h8220000;
      30202: inst = 32'h10408000;
      30203: inst = 32'hc40436a;
      30204: inst = 32'h8220000;
      30205: inst = 32'h10408000;
      30206: inst = 32'hc40436b;
      30207: inst = 32'h8220000;
      30208: inst = 32'h10408000;
      30209: inst = 32'hc40436c;
      30210: inst = 32'h8220000;
      30211: inst = 32'h10408000;
      30212: inst = 32'hc40436d;
      30213: inst = 32'h8220000;
      30214: inst = 32'h10408000;
      30215: inst = 32'hc40436e;
      30216: inst = 32'h8220000;
      30217: inst = 32'h10408000;
      30218: inst = 32'hc40436f;
      30219: inst = 32'h8220000;
      30220: inst = 32'h10408000;
      30221: inst = 32'hc404370;
      30222: inst = 32'h8220000;
      30223: inst = 32'h10408000;
      30224: inst = 32'hc404371;
      30225: inst = 32'h8220000;
      30226: inst = 32'h10408000;
      30227: inst = 32'hc404372;
      30228: inst = 32'h8220000;
      30229: inst = 32'h10408000;
      30230: inst = 32'hc404373;
      30231: inst = 32'h8220000;
      30232: inst = 32'h10408000;
      30233: inst = 32'hc404374;
      30234: inst = 32'h8220000;
      30235: inst = 32'h10408000;
      30236: inst = 32'hc404375;
      30237: inst = 32'h8220000;
      30238: inst = 32'h10408000;
      30239: inst = 32'hc404376;
      30240: inst = 32'h8220000;
      30241: inst = 32'h10408000;
      30242: inst = 32'hc404377;
      30243: inst = 32'h8220000;
      30244: inst = 32'h10408000;
      30245: inst = 32'hc404378;
      30246: inst = 32'h8220000;
      30247: inst = 32'h10408000;
      30248: inst = 32'hc404379;
      30249: inst = 32'h8220000;
      30250: inst = 32'h10408000;
      30251: inst = 32'hc40437a;
      30252: inst = 32'h8220000;
      30253: inst = 32'h10408000;
      30254: inst = 32'hc40437b;
      30255: inst = 32'h8220000;
      30256: inst = 32'h10408000;
      30257: inst = 32'hc40437c;
      30258: inst = 32'h8220000;
      30259: inst = 32'h10408000;
      30260: inst = 32'hc40437d;
      30261: inst = 32'h8220000;
      30262: inst = 32'h10408000;
      30263: inst = 32'hc40437e;
      30264: inst = 32'h8220000;
      30265: inst = 32'h10408000;
      30266: inst = 32'hc40437f;
      30267: inst = 32'h8220000;
      30268: inst = 32'h10408000;
      30269: inst = 32'hc404380;
      30270: inst = 32'h8220000;
      30271: inst = 32'h10408000;
      30272: inst = 32'hc404381;
      30273: inst = 32'h8220000;
      30274: inst = 32'h10408000;
      30275: inst = 32'hc404382;
      30276: inst = 32'h8220000;
      30277: inst = 32'h10408000;
      30278: inst = 32'hc404383;
      30279: inst = 32'h8220000;
      30280: inst = 32'h10408000;
      30281: inst = 32'hc404384;
      30282: inst = 32'h8220000;
      30283: inst = 32'h10408000;
      30284: inst = 32'hc404385;
      30285: inst = 32'h8220000;
      30286: inst = 32'h10408000;
      30287: inst = 32'hc404386;
      30288: inst = 32'h8220000;
      30289: inst = 32'h10408000;
      30290: inst = 32'hc404387;
      30291: inst = 32'h8220000;
      30292: inst = 32'h10408000;
      30293: inst = 32'hc404388;
      30294: inst = 32'h8220000;
      30295: inst = 32'h10408000;
      30296: inst = 32'hc404389;
      30297: inst = 32'h8220000;
      30298: inst = 32'h10408000;
      30299: inst = 32'hc40438a;
      30300: inst = 32'h8220000;
      30301: inst = 32'h10408000;
      30302: inst = 32'hc40438b;
      30303: inst = 32'h8220000;
      30304: inst = 32'h10408000;
      30305: inst = 32'hc40438f;
      30306: inst = 32'h8220000;
      30307: inst = 32'h10408000;
      30308: inst = 32'hc404390;
      30309: inst = 32'h8220000;
      30310: inst = 32'h10408000;
      30311: inst = 32'hc4043a3;
      30312: inst = 32'h8220000;
      30313: inst = 32'h10408000;
      30314: inst = 32'hc4043ad;
      30315: inst = 32'h8220000;
      30316: inst = 32'h10408000;
      30317: inst = 32'hc4043ae;
      30318: inst = 32'h8220000;
      30319: inst = 32'h10408000;
      30320: inst = 32'hc4043af;
      30321: inst = 32'h8220000;
      30322: inst = 32'h10408000;
      30323: inst = 32'hc4043b0;
      30324: inst = 32'h8220000;
      30325: inst = 32'h10408000;
      30326: inst = 32'hc4043b1;
      30327: inst = 32'h8220000;
      30328: inst = 32'h10408000;
      30329: inst = 32'hc4043b2;
      30330: inst = 32'h8220000;
      30331: inst = 32'h10408000;
      30332: inst = 32'hc4043b3;
      30333: inst = 32'h8220000;
      30334: inst = 32'h10408000;
      30335: inst = 32'hc4043b4;
      30336: inst = 32'h8220000;
      30337: inst = 32'h10408000;
      30338: inst = 32'hc4043b5;
      30339: inst = 32'h8220000;
      30340: inst = 32'h10408000;
      30341: inst = 32'hc4043b6;
      30342: inst = 32'h8220000;
      30343: inst = 32'h10408000;
      30344: inst = 32'hc4043b7;
      30345: inst = 32'h8220000;
      30346: inst = 32'h10408000;
      30347: inst = 32'hc4043b8;
      30348: inst = 32'h8220000;
      30349: inst = 32'h10408000;
      30350: inst = 32'hc4043b9;
      30351: inst = 32'h8220000;
      30352: inst = 32'h10408000;
      30353: inst = 32'hc4043ba;
      30354: inst = 32'h8220000;
      30355: inst = 32'h10408000;
      30356: inst = 32'hc4043bb;
      30357: inst = 32'h8220000;
      30358: inst = 32'h10408000;
      30359: inst = 32'hc4043bc;
      30360: inst = 32'h8220000;
      30361: inst = 32'h10408000;
      30362: inst = 32'hc4043bd;
      30363: inst = 32'h8220000;
      30364: inst = 32'h10408000;
      30365: inst = 32'hc4043be;
      30366: inst = 32'h8220000;
      30367: inst = 32'h10408000;
      30368: inst = 32'hc4043bf;
      30369: inst = 32'h8220000;
      30370: inst = 32'h10408000;
      30371: inst = 32'hc4043c0;
      30372: inst = 32'h8220000;
      30373: inst = 32'h10408000;
      30374: inst = 32'hc4043c1;
      30375: inst = 32'h8220000;
      30376: inst = 32'h10408000;
      30377: inst = 32'hc4043c2;
      30378: inst = 32'h8220000;
      30379: inst = 32'h10408000;
      30380: inst = 32'hc4043c3;
      30381: inst = 32'h8220000;
      30382: inst = 32'h10408000;
      30383: inst = 32'hc4043c4;
      30384: inst = 32'h8220000;
      30385: inst = 32'h10408000;
      30386: inst = 32'hc4043c5;
      30387: inst = 32'h8220000;
      30388: inst = 32'h10408000;
      30389: inst = 32'hc4043c6;
      30390: inst = 32'h8220000;
      30391: inst = 32'h10408000;
      30392: inst = 32'hc4043c7;
      30393: inst = 32'h8220000;
      30394: inst = 32'h10408000;
      30395: inst = 32'hc4043c8;
      30396: inst = 32'h8220000;
      30397: inst = 32'h10408000;
      30398: inst = 32'hc4043c9;
      30399: inst = 32'h8220000;
      30400: inst = 32'h10408000;
      30401: inst = 32'hc4043ca;
      30402: inst = 32'h8220000;
      30403: inst = 32'h10408000;
      30404: inst = 32'hc4043cb;
      30405: inst = 32'h8220000;
      30406: inst = 32'h10408000;
      30407: inst = 32'hc4043cc;
      30408: inst = 32'h8220000;
      30409: inst = 32'h10408000;
      30410: inst = 32'hc4043cd;
      30411: inst = 32'h8220000;
      30412: inst = 32'h10408000;
      30413: inst = 32'hc4043ce;
      30414: inst = 32'h8220000;
      30415: inst = 32'h10408000;
      30416: inst = 32'hc4043cf;
      30417: inst = 32'h8220000;
      30418: inst = 32'h10408000;
      30419: inst = 32'hc4043d0;
      30420: inst = 32'h8220000;
      30421: inst = 32'h10408000;
      30422: inst = 32'hc4043d1;
      30423: inst = 32'h8220000;
      30424: inst = 32'h10408000;
      30425: inst = 32'hc4043d2;
      30426: inst = 32'h8220000;
      30427: inst = 32'h10408000;
      30428: inst = 32'hc4043d3;
      30429: inst = 32'h8220000;
      30430: inst = 32'h10408000;
      30431: inst = 32'hc4043d4;
      30432: inst = 32'h8220000;
      30433: inst = 32'h10408000;
      30434: inst = 32'hc4043d5;
      30435: inst = 32'h8220000;
      30436: inst = 32'h10408000;
      30437: inst = 32'hc4043d6;
      30438: inst = 32'h8220000;
      30439: inst = 32'h10408000;
      30440: inst = 32'hc4043d7;
      30441: inst = 32'h8220000;
      30442: inst = 32'h10408000;
      30443: inst = 32'hc4043d8;
      30444: inst = 32'h8220000;
      30445: inst = 32'h10408000;
      30446: inst = 32'hc4043d9;
      30447: inst = 32'h8220000;
      30448: inst = 32'h10408000;
      30449: inst = 32'hc4043da;
      30450: inst = 32'h8220000;
      30451: inst = 32'h10408000;
      30452: inst = 32'hc4043db;
      30453: inst = 32'h8220000;
      30454: inst = 32'h10408000;
      30455: inst = 32'hc4043dc;
      30456: inst = 32'h8220000;
      30457: inst = 32'h10408000;
      30458: inst = 32'hc4043dd;
      30459: inst = 32'h8220000;
      30460: inst = 32'h10408000;
      30461: inst = 32'hc4043de;
      30462: inst = 32'h8220000;
      30463: inst = 32'h10408000;
      30464: inst = 32'hc4043df;
      30465: inst = 32'h8220000;
      30466: inst = 32'h10408000;
      30467: inst = 32'hc4043e0;
      30468: inst = 32'h8220000;
      30469: inst = 32'h10408000;
      30470: inst = 32'hc4043e1;
      30471: inst = 32'h8220000;
      30472: inst = 32'h10408000;
      30473: inst = 32'hc4043e2;
      30474: inst = 32'h8220000;
      30475: inst = 32'h10408000;
      30476: inst = 32'hc4043e3;
      30477: inst = 32'h8220000;
      30478: inst = 32'h10408000;
      30479: inst = 32'hc4043e4;
      30480: inst = 32'h8220000;
      30481: inst = 32'h10408000;
      30482: inst = 32'hc4043e5;
      30483: inst = 32'h8220000;
      30484: inst = 32'h10408000;
      30485: inst = 32'hc4043e6;
      30486: inst = 32'h8220000;
      30487: inst = 32'h10408000;
      30488: inst = 32'hc4043e7;
      30489: inst = 32'h8220000;
      30490: inst = 32'h10408000;
      30491: inst = 32'hc4043e8;
      30492: inst = 32'h8220000;
      30493: inst = 32'h10408000;
      30494: inst = 32'hc4043e9;
      30495: inst = 32'h8220000;
      30496: inst = 32'h10408000;
      30497: inst = 32'hc4043ea;
      30498: inst = 32'h8220000;
      30499: inst = 32'h10408000;
      30500: inst = 32'hc4043eb;
      30501: inst = 32'h8220000;
      30502: inst = 32'h10408000;
      30503: inst = 32'hc4043ef;
      30504: inst = 32'h8220000;
      30505: inst = 32'h10408000;
      30506: inst = 32'hc4043f9;
      30507: inst = 32'h8220000;
      30508: inst = 32'h10408000;
      30509: inst = 32'hc404403;
      30510: inst = 32'h8220000;
      30511: inst = 32'h10408000;
      30512: inst = 32'hc404404;
      30513: inst = 32'h8220000;
      30514: inst = 32'h10408000;
      30515: inst = 32'hc404405;
      30516: inst = 32'h8220000;
      30517: inst = 32'h10408000;
      30518: inst = 32'hc404406;
      30519: inst = 32'h8220000;
      30520: inst = 32'h10408000;
      30521: inst = 32'hc404407;
      30522: inst = 32'h8220000;
      30523: inst = 32'h10408000;
      30524: inst = 32'hc404408;
      30525: inst = 32'h8220000;
      30526: inst = 32'h10408000;
      30527: inst = 32'hc404409;
      30528: inst = 32'h8220000;
      30529: inst = 32'h10408000;
      30530: inst = 32'hc40440a;
      30531: inst = 32'h8220000;
      30532: inst = 32'h10408000;
      30533: inst = 32'hc40440b;
      30534: inst = 32'h8220000;
      30535: inst = 32'h10408000;
      30536: inst = 32'hc40440c;
      30537: inst = 32'h8220000;
      30538: inst = 32'h10408000;
      30539: inst = 32'hc40440d;
      30540: inst = 32'h8220000;
      30541: inst = 32'h10408000;
      30542: inst = 32'hc40440e;
      30543: inst = 32'h8220000;
      30544: inst = 32'h10408000;
      30545: inst = 32'hc40440f;
      30546: inst = 32'h8220000;
      30547: inst = 32'h10408000;
      30548: inst = 32'hc404410;
      30549: inst = 32'h8220000;
      30550: inst = 32'h10408000;
      30551: inst = 32'hc404411;
      30552: inst = 32'h8220000;
      30553: inst = 32'h10408000;
      30554: inst = 32'hc404412;
      30555: inst = 32'h8220000;
      30556: inst = 32'h10408000;
      30557: inst = 32'hc404413;
      30558: inst = 32'h8220000;
      30559: inst = 32'h10408000;
      30560: inst = 32'hc404414;
      30561: inst = 32'h8220000;
      30562: inst = 32'h10408000;
      30563: inst = 32'hc404415;
      30564: inst = 32'h8220000;
      30565: inst = 32'h10408000;
      30566: inst = 32'hc404416;
      30567: inst = 32'h8220000;
      30568: inst = 32'h10408000;
      30569: inst = 32'hc404417;
      30570: inst = 32'h8220000;
      30571: inst = 32'h10408000;
      30572: inst = 32'hc404418;
      30573: inst = 32'h8220000;
      30574: inst = 32'h10408000;
      30575: inst = 32'hc404419;
      30576: inst = 32'h8220000;
      30577: inst = 32'h10408000;
      30578: inst = 32'hc40441a;
      30579: inst = 32'h8220000;
      30580: inst = 32'h10408000;
      30581: inst = 32'hc40441b;
      30582: inst = 32'h8220000;
      30583: inst = 32'h10408000;
      30584: inst = 32'hc40441c;
      30585: inst = 32'h8220000;
      30586: inst = 32'h10408000;
      30587: inst = 32'hc40441d;
      30588: inst = 32'h8220000;
      30589: inst = 32'h10408000;
      30590: inst = 32'hc40441e;
      30591: inst = 32'h8220000;
      30592: inst = 32'h10408000;
      30593: inst = 32'hc40441f;
      30594: inst = 32'h8220000;
      30595: inst = 32'h10408000;
      30596: inst = 32'hc404420;
      30597: inst = 32'h8220000;
      30598: inst = 32'h10408000;
      30599: inst = 32'hc404421;
      30600: inst = 32'h8220000;
      30601: inst = 32'h10408000;
      30602: inst = 32'hc404422;
      30603: inst = 32'h8220000;
      30604: inst = 32'h10408000;
      30605: inst = 32'hc404423;
      30606: inst = 32'h8220000;
      30607: inst = 32'h10408000;
      30608: inst = 32'hc404424;
      30609: inst = 32'h8220000;
      30610: inst = 32'h10408000;
      30611: inst = 32'hc404425;
      30612: inst = 32'h8220000;
      30613: inst = 32'h10408000;
      30614: inst = 32'hc404426;
      30615: inst = 32'h8220000;
      30616: inst = 32'h10408000;
      30617: inst = 32'hc404427;
      30618: inst = 32'h8220000;
      30619: inst = 32'h10408000;
      30620: inst = 32'hc404428;
      30621: inst = 32'h8220000;
      30622: inst = 32'h10408000;
      30623: inst = 32'hc404429;
      30624: inst = 32'h8220000;
      30625: inst = 32'h10408000;
      30626: inst = 32'hc40442a;
      30627: inst = 32'h8220000;
      30628: inst = 32'h10408000;
      30629: inst = 32'hc40442b;
      30630: inst = 32'h8220000;
      30631: inst = 32'h10408000;
      30632: inst = 32'hc40442c;
      30633: inst = 32'h8220000;
      30634: inst = 32'h10408000;
      30635: inst = 32'hc40442d;
      30636: inst = 32'h8220000;
      30637: inst = 32'h10408000;
      30638: inst = 32'hc40442e;
      30639: inst = 32'h8220000;
      30640: inst = 32'h10408000;
      30641: inst = 32'hc40442f;
      30642: inst = 32'h8220000;
      30643: inst = 32'h10408000;
      30644: inst = 32'hc404430;
      30645: inst = 32'h8220000;
      30646: inst = 32'h10408000;
      30647: inst = 32'hc404431;
      30648: inst = 32'h8220000;
      30649: inst = 32'h10408000;
      30650: inst = 32'hc404432;
      30651: inst = 32'h8220000;
      30652: inst = 32'h10408000;
      30653: inst = 32'hc404433;
      30654: inst = 32'h8220000;
      30655: inst = 32'h10408000;
      30656: inst = 32'hc404434;
      30657: inst = 32'h8220000;
      30658: inst = 32'h10408000;
      30659: inst = 32'hc404435;
      30660: inst = 32'h8220000;
      30661: inst = 32'h10408000;
      30662: inst = 32'hc404436;
      30663: inst = 32'h8220000;
      30664: inst = 32'h10408000;
      30665: inst = 32'hc404437;
      30666: inst = 32'h8220000;
      30667: inst = 32'h10408000;
      30668: inst = 32'hc404438;
      30669: inst = 32'h8220000;
      30670: inst = 32'h10408000;
      30671: inst = 32'hc404439;
      30672: inst = 32'h8220000;
      30673: inst = 32'h10408000;
      30674: inst = 32'hc40443a;
      30675: inst = 32'h8220000;
      30676: inst = 32'h10408000;
      30677: inst = 32'hc40443b;
      30678: inst = 32'h8220000;
      30679: inst = 32'h10408000;
      30680: inst = 32'hc40443c;
      30681: inst = 32'h8220000;
      30682: inst = 32'h10408000;
      30683: inst = 32'hc40443d;
      30684: inst = 32'h8220000;
      30685: inst = 32'h10408000;
      30686: inst = 32'hc40443e;
      30687: inst = 32'h8220000;
      30688: inst = 32'h10408000;
      30689: inst = 32'hc40443f;
      30690: inst = 32'h8220000;
      30691: inst = 32'h10408000;
      30692: inst = 32'hc404440;
      30693: inst = 32'h8220000;
      30694: inst = 32'h10408000;
      30695: inst = 32'hc404441;
      30696: inst = 32'h8220000;
      30697: inst = 32'h10408000;
      30698: inst = 32'hc404442;
      30699: inst = 32'h8220000;
      30700: inst = 32'h10408000;
      30701: inst = 32'hc404443;
      30702: inst = 32'h8220000;
      30703: inst = 32'h10408000;
      30704: inst = 32'hc404444;
      30705: inst = 32'h8220000;
      30706: inst = 32'h10408000;
      30707: inst = 32'hc404445;
      30708: inst = 32'h8220000;
      30709: inst = 32'h10408000;
      30710: inst = 32'hc404446;
      30711: inst = 32'h8220000;
      30712: inst = 32'h10408000;
      30713: inst = 32'hc404447;
      30714: inst = 32'h8220000;
      30715: inst = 32'h10408000;
      30716: inst = 32'hc404448;
      30717: inst = 32'h8220000;
      30718: inst = 32'h10408000;
      30719: inst = 32'hc404449;
      30720: inst = 32'h8220000;
      30721: inst = 32'h10408000;
      30722: inst = 32'hc40444a;
      30723: inst = 32'h8220000;
      30724: inst = 32'h10408000;
      30725: inst = 32'hc40444b;
      30726: inst = 32'h8220000;
      30727: inst = 32'h10408000;
      30728: inst = 32'hc40444f;
      30729: inst = 32'h8220000;
      30730: inst = 32'h10408000;
      30731: inst = 32'hc404455;
      30732: inst = 32'h8220000;
      30733: inst = 32'h10408000;
      30734: inst = 32'hc404463;
      30735: inst = 32'h8220000;
      30736: inst = 32'h10408000;
      30737: inst = 32'hc404464;
      30738: inst = 32'h8220000;
      30739: inst = 32'h10408000;
      30740: inst = 32'hc404465;
      30741: inst = 32'h8220000;
      30742: inst = 32'h10408000;
      30743: inst = 32'hc404466;
      30744: inst = 32'h8220000;
      30745: inst = 32'h10408000;
      30746: inst = 32'hc404467;
      30747: inst = 32'h8220000;
      30748: inst = 32'h10408000;
      30749: inst = 32'hc404468;
      30750: inst = 32'h8220000;
      30751: inst = 32'h10408000;
      30752: inst = 32'hc404469;
      30753: inst = 32'h8220000;
      30754: inst = 32'h10408000;
      30755: inst = 32'hc40446a;
      30756: inst = 32'h8220000;
      30757: inst = 32'h10408000;
      30758: inst = 32'hc40446b;
      30759: inst = 32'h8220000;
      30760: inst = 32'h10408000;
      30761: inst = 32'hc40446c;
      30762: inst = 32'h8220000;
      30763: inst = 32'h10408000;
      30764: inst = 32'hc40446d;
      30765: inst = 32'h8220000;
      30766: inst = 32'h10408000;
      30767: inst = 32'hc40446e;
      30768: inst = 32'h8220000;
      30769: inst = 32'h10408000;
      30770: inst = 32'hc40446f;
      30771: inst = 32'h8220000;
      30772: inst = 32'h10408000;
      30773: inst = 32'hc404470;
      30774: inst = 32'h8220000;
      30775: inst = 32'h10408000;
      30776: inst = 32'hc404471;
      30777: inst = 32'h8220000;
      30778: inst = 32'h10408000;
      30779: inst = 32'hc404472;
      30780: inst = 32'h8220000;
      30781: inst = 32'h10408000;
      30782: inst = 32'hc404473;
      30783: inst = 32'h8220000;
      30784: inst = 32'h10408000;
      30785: inst = 32'hc404474;
      30786: inst = 32'h8220000;
      30787: inst = 32'h10408000;
      30788: inst = 32'hc404475;
      30789: inst = 32'h8220000;
      30790: inst = 32'h10408000;
      30791: inst = 32'hc404476;
      30792: inst = 32'h8220000;
      30793: inst = 32'h10408000;
      30794: inst = 32'hc404477;
      30795: inst = 32'h8220000;
      30796: inst = 32'h10408000;
      30797: inst = 32'hc404478;
      30798: inst = 32'h8220000;
      30799: inst = 32'h10408000;
      30800: inst = 32'hc404479;
      30801: inst = 32'h8220000;
      30802: inst = 32'h10408000;
      30803: inst = 32'hc40447a;
      30804: inst = 32'h8220000;
      30805: inst = 32'h10408000;
      30806: inst = 32'hc40447b;
      30807: inst = 32'h8220000;
      30808: inst = 32'h10408000;
      30809: inst = 32'hc40447c;
      30810: inst = 32'h8220000;
      30811: inst = 32'h10408000;
      30812: inst = 32'hc40447d;
      30813: inst = 32'h8220000;
      30814: inst = 32'h10408000;
      30815: inst = 32'hc40447e;
      30816: inst = 32'h8220000;
      30817: inst = 32'h10408000;
      30818: inst = 32'hc40447f;
      30819: inst = 32'h8220000;
      30820: inst = 32'h10408000;
      30821: inst = 32'hc404480;
      30822: inst = 32'h8220000;
      30823: inst = 32'h10408000;
      30824: inst = 32'hc404481;
      30825: inst = 32'h8220000;
      30826: inst = 32'h10408000;
      30827: inst = 32'hc404482;
      30828: inst = 32'h8220000;
      30829: inst = 32'h10408000;
      30830: inst = 32'hc404483;
      30831: inst = 32'h8220000;
      30832: inst = 32'h10408000;
      30833: inst = 32'hc404484;
      30834: inst = 32'h8220000;
      30835: inst = 32'h10408000;
      30836: inst = 32'hc404485;
      30837: inst = 32'h8220000;
      30838: inst = 32'h10408000;
      30839: inst = 32'hc404486;
      30840: inst = 32'h8220000;
      30841: inst = 32'h10408000;
      30842: inst = 32'hc404487;
      30843: inst = 32'h8220000;
      30844: inst = 32'h10408000;
      30845: inst = 32'hc404488;
      30846: inst = 32'h8220000;
      30847: inst = 32'h10408000;
      30848: inst = 32'hc404489;
      30849: inst = 32'h8220000;
      30850: inst = 32'h10408000;
      30851: inst = 32'hc40448a;
      30852: inst = 32'h8220000;
      30853: inst = 32'h10408000;
      30854: inst = 32'hc40448b;
      30855: inst = 32'h8220000;
      30856: inst = 32'h10408000;
      30857: inst = 32'hc40448c;
      30858: inst = 32'h8220000;
      30859: inst = 32'h10408000;
      30860: inst = 32'hc40448d;
      30861: inst = 32'h8220000;
      30862: inst = 32'h10408000;
      30863: inst = 32'hc40448e;
      30864: inst = 32'h8220000;
      30865: inst = 32'h10408000;
      30866: inst = 32'hc40448f;
      30867: inst = 32'h8220000;
      30868: inst = 32'h10408000;
      30869: inst = 32'hc404490;
      30870: inst = 32'h8220000;
      30871: inst = 32'h10408000;
      30872: inst = 32'hc404491;
      30873: inst = 32'h8220000;
      30874: inst = 32'h10408000;
      30875: inst = 32'hc404492;
      30876: inst = 32'h8220000;
      30877: inst = 32'h10408000;
      30878: inst = 32'hc404493;
      30879: inst = 32'h8220000;
      30880: inst = 32'h10408000;
      30881: inst = 32'hc404494;
      30882: inst = 32'h8220000;
      30883: inst = 32'h10408000;
      30884: inst = 32'hc404495;
      30885: inst = 32'h8220000;
      30886: inst = 32'h10408000;
      30887: inst = 32'hc404496;
      30888: inst = 32'h8220000;
      30889: inst = 32'h10408000;
      30890: inst = 32'hc404497;
      30891: inst = 32'h8220000;
      30892: inst = 32'h10408000;
      30893: inst = 32'hc404498;
      30894: inst = 32'h8220000;
      30895: inst = 32'h10408000;
      30896: inst = 32'hc404499;
      30897: inst = 32'h8220000;
      30898: inst = 32'h10408000;
      30899: inst = 32'hc40449a;
      30900: inst = 32'h8220000;
      30901: inst = 32'h10408000;
      30902: inst = 32'hc40449b;
      30903: inst = 32'h8220000;
      30904: inst = 32'h10408000;
      30905: inst = 32'hc40449c;
      30906: inst = 32'h8220000;
      30907: inst = 32'h10408000;
      30908: inst = 32'hc40449d;
      30909: inst = 32'h8220000;
      30910: inst = 32'h10408000;
      30911: inst = 32'hc40449e;
      30912: inst = 32'h8220000;
      30913: inst = 32'h10408000;
      30914: inst = 32'hc40449f;
      30915: inst = 32'h8220000;
      30916: inst = 32'h10408000;
      30917: inst = 32'hc4044a0;
      30918: inst = 32'h8220000;
      30919: inst = 32'h10408000;
      30920: inst = 32'hc4044a1;
      30921: inst = 32'h8220000;
      30922: inst = 32'h10408000;
      30923: inst = 32'hc4044a2;
      30924: inst = 32'h8220000;
      30925: inst = 32'h10408000;
      30926: inst = 32'hc4044a3;
      30927: inst = 32'h8220000;
      30928: inst = 32'h10408000;
      30929: inst = 32'hc4044a4;
      30930: inst = 32'h8220000;
      30931: inst = 32'h10408000;
      30932: inst = 32'hc4044a5;
      30933: inst = 32'h8220000;
      30934: inst = 32'h10408000;
      30935: inst = 32'hc4044a6;
      30936: inst = 32'h8220000;
      30937: inst = 32'h10408000;
      30938: inst = 32'hc4044a7;
      30939: inst = 32'h8220000;
      30940: inst = 32'h10408000;
      30941: inst = 32'hc4044a8;
      30942: inst = 32'h8220000;
      30943: inst = 32'h10408000;
      30944: inst = 32'hc4044a9;
      30945: inst = 32'h8220000;
      30946: inst = 32'h10408000;
      30947: inst = 32'hc4044aa;
      30948: inst = 32'h8220000;
      30949: inst = 32'h10408000;
      30950: inst = 32'hc4044ab;
      30951: inst = 32'h8220000;
      30952: inst = 32'h10408000;
      30953: inst = 32'hc4044af;
      30954: inst = 32'h8220000;
      30955: inst = 32'h10408000;
      30956: inst = 32'hc4044b0;
      30957: inst = 32'h8220000;
      30958: inst = 32'h10408000;
      30959: inst = 32'hc4044b1;
      30960: inst = 32'h8220000;
      30961: inst = 32'h10408000;
      30962: inst = 32'hc4044b2;
      30963: inst = 32'h8220000;
      30964: inst = 32'h10408000;
      30965: inst = 32'hc4044b7;
      30966: inst = 32'h8220000;
      30967: inst = 32'h10408000;
      30968: inst = 32'hc4044c3;
      30969: inst = 32'h8220000;
      30970: inst = 32'h10408000;
      30971: inst = 32'hc4044c4;
      30972: inst = 32'h8220000;
      30973: inst = 32'h10408000;
      30974: inst = 32'hc4044c5;
      30975: inst = 32'h8220000;
      30976: inst = 32'h10408000;
      30977: inst = 32'hc4044c6;
      30978: inst = 32'h8220000;
      30979: inst = 32'h10408000;
      30980: inst = 32'hc4044c7;
      30981: inst = 32'h8220000;
      30982: inst = 32'h10408000;
      30983: inst = 32'hc4044c8;
      30984: inst = 32'h8220000;
      30985: inst = 32'h10408000;
      30986: inst = 32'hc4044c9;
      30987: inst = 32'h8220000;
      30988: inst = 32'h10408000;
      30989: inst = 32'hc4044ca;
      30990: inst = 32'h8220000;
      30991: inst = 32'h10408000;
      30992: inst = 32'hc4044cb;
      30993: inst = 32'h8220000;
      30994: inst = 32'h10408000;
      30995: inst = 32'hc4044cc;
      30996: inst = 32'h8220000;
      30997: inst = 32'h10408000;
      30998: inst = 32'hc4044cd;
      30999: inst = 32'h8220000;
      31000: inst = 32'h10408000;
      31001: inst = 32'hc4044ce;
      31002: inst = 32'h8220000;
      31003: inst = 32'h10408000;
      31004: inst = 32'hc4044cf;
      31005: inst = 32'h8220000;
      31006: inst = 32'h10408000;
      31007: inst = 32'hc4044d0;
      31008: inst = 32'h8220000;
      31009: inst = 32'h10408000;
      31010: inst = 32'hc4044d1;
      31011: inst = 32'h8220000;
      31012: inst = 32'h10408000;
      31013: inst = 32'hc4044d2;
      31014: inst = 32'h8220000;
      31015: inst = 32'h10408000;
      31016: inst = 32'hc4044d3;
      31017: inst = 32'h8220000;
      31018: inst = 32'h10408000;
      31019: inst = 32'hc4044d4;
      31020: inst = 32'h8220000;
      31021: inst = 32'h10408000;
      31022: inst = 32'hc4044d5;
      31023: inst = 32'h8220000;
      31024: inst = 32'h10408000;
      31025: inst = 32'hc4044d6;
      31026: inst = 32'h8220000;
      31027: inst = 32'h10408000;
      31028: inst = 32'hc4044d7;
      31029: inst = 32'h8220000;
      31030: inst = 32'h10408000;
      31031: inst = 32'hc4044d8;
      31032: inst = 32'h8220000;
      31033: inst = 32'h10408000;
      31034: inst = 32'hc4044d9;
      31035: inst = 32'h8220000;
      31036: inst = 32'h10408000;
      31037: inst = 32'hc4044da;
      31038: inst = 32'h8220000;
      31039: inst = 32'h10408000;
      31040: inst = 32'hc4044db;
      31041: inst = 32'h8220000;
      31042: inst = 32'h10408000;
      31043: inst = 32'hc4044dc;
      31044: inst = 32'h8220000;
      31045: inst = 32'h10408000;
      31046: inst = 32'hc4044dd;
      31047: inst = 32'h8220000;
      31048: inst = 32'h10408000;
      31049: inst = 32'hc4044de;
      31050: inst = 32'h8220000;
      31051: inst = 32'h10408000;
      31052: inst = 32'hc4044df;
      31053: inst = 32'h8220000;
      31054: inst = 32'h10408000;
      31055: inst = 32'hc4044e0;
      31056: inst = 32'h8220000;
      31057: inst = 32'h10408000;
      31058: inst = 32'hc4044e1;
      31059: inst = 32'h8220000;
      31060: inst = 32'h10408000;
      31061: inst = 32'hc4044e2;
      31062: inst = 32'h8220000;
      31063: inst = 32'h10408000;
      31064: inst = 32'hc4044e3;
      31065: inst = 32'h8220000;
      31066: inst = 32'h10408000;
      31067: inst = 32'hc4044e4;
      31068: inst = 32'h8220000;
      31069: inst = 32'h10408000;
      31070: inst = 32'hc4044e5;
      31071: inst = 32'h8220000;
      31072: inst = 32'h10408000;
      31073: inst = 32'hc4044e6;
      31074: inst = 32'h8220000;
      31075: inst = 32'h10408000;
      31076: inst = 32'hc4044e7;
      31077: inst = 32'h8220000;
      31078: inst = 32'h10408000;
      31079: inst = 32'hc4044e8;
      31080: inst = 32'h8220000;
      31081: inst = 32'h10408000;
      31082: inst = 32'hc4044e9;
      31083: inst = 32'h8220000;
      31084: inst = 32'h10408000;
      31085: inst = 32'hc4044ea;
      31086: inst = 32'h8220000;
      31087: inst = 32'h10408000;
      31088: inst = 32'hc4044eb;
      31089: inst = 32'h8220000;
      31090: inst = 32'h10408000;
      31091: inst = 32'hc4044ec;
      31092: inst = 32'h8220000;
      31093: inst = 32'h10408000;
      31094: inst = 32'hc4044ed;
      31095: inst = 32'h8220000;
      31096: inst = 32'h10408000;
      31097: inst = 32'hc4044ee;
      31098: inst = 32'h8220000;
      31099: inst = 32'h10408000;
      31100: inst = 32'hc4044ef;
      31101: inst = 32'h8220000;
      31102: inst = 32'h10408000;
      31103: inst = 32'hc4044f0;
      31104: inst = 32'h8220000;
      31105: inst = 32'h10408000;
      31106: inst = 32'hc4044f1;
      31107: inst = 32'h8220000;
      31108: inst = 32'h10408000;
      31109: inst = 32'hc4044f2;
      31110: inst = 32'h8220000;
      31111: inst = 32'h10408000;
      31112: inst = 32'hc4044f3;
      31113: inst = 32'h8220000;
      31114: inst = 32'h10408000;
      31115: inst = 32'hc4044f4;
      31116: inst = 32'h8220000;
      31117: inst = 32'h10408000;
      31118: inst = 32'hc4044f5;
      31119: inst = 32'h8220000;
      31120: inst = 32'h10408000;
      31121: inst = 32'hc4044f6;
      31122: inst = 32'h8220000;
      31123: inst = 32'h10408000;
      31124: inst = 32'hc4044f7;
      31125: inst = 32'h8220000;
      31126: inst = 32'h10408000;
      31127: inst = 32'hc4044f8;
      31128: inst = 32'h8220000;
      31129: inst = 32'h10408000;
      31130: inst = 32'hc4044f9;
      31131: inst = 32'h8220000;
      31132: inst = 32'h10408000;
      31133: inst = 32'hc4044fa;
      31134: inst = 32'h8220000;
      31135: inst = 32'h10408000;
      31136: inst = 32'hc4044fb;
      31137: inst = 32'h8220000;
      31138: inst = 32'h10408000;
      31139: inst = 32'hc4044fc;
      31140: inst = 32'h8220000;
      31141: inst = 32'h10408000;
      31142: inst = 32'hc4044fd;
      31143: inst = 32'h8220000;
      31144: inst = 32'h10408000;
      31145: inst = 32'hc4044fe;
      31146: inst = 32'h8220000;
      31147: inst = 32'h10408000;
      31148: inst = 32'hc4044ff;
      31149: inst = 32'h8220000;
      31150: inst = 32'h10408000;
      31151: inst = 32'hc404500;
      31152: inst = 32'h8220000;
      31153: inst = 32'h10408000;
      31154: inst = 32'hc404501;
      31155: inst = 32'h8220000;
      31156: inst = 32'h10408000;
      31157: inst = 32'hc404502;
      31158: inst = 32'h8220000;
      31159: inst = 32'h10408000;
      31160: inst = 32'hc404503;
      31161: inst = 32'h8220000;
      31162: inst = 32'h10408000;
      31163: inst = 32'hc404504;
      31164: inst = 32'h8220000;
      31165: inst = 32'h10408000;
      31166: inst = 32'hc404505;
      31167: inst = 32'h8220000;
      31168: inst = 32'h10408000;
      31169: inst = 32'hc404506;
      31170: inst = 32'h8220000;
      31171: inst = 32'h10408000;
      31172: inst = 32'hc404507;
      31173: inst = 32'h8220000;
      31174: inst = 32'h10408000;
      31175: inst = 32'hc404508;
      31176: inst = 32'h8220000;
      31177: inst = 32'h10408000;
      31178: inst = 32'hc404509;
      31179: inst = 32'h8220000;
      31180: inst = 32'h10408000;
      31181: inst = 32'hc40450a;
      31182: inst = 32'h8220000;
      31183: inst = 32'h10408000;
      31184: inst = 32'hc40450b;
      31185: inst = 32'h8220000;
      31186: inst = 32'h10408000;
      31187: inst = 32'hc40450f;
      31188: inst = 32'h8220000;
      31189: inst = 32'h10408000;
      31190: inst = 32'hc404512;
      31191: inst = 32'h8220000;
      31192: inst = 32'h10408000;
      31193: inst = 32'hc404513;
      31194: inst = 32'h8220000;
      31195: inst = 32'h10408000;
      31196: inst = 32'hc404523;
      31197: inst = 32'h8220000;
      31198: inst = 32'h10408000;
      31199: inst = 32'hc404524;
      31200: inst = 32'h8220000;
      31201: inst = 32'h10408000;
      31202: inst = 32'hc404525;
      31203: inst = 32'h8220000;
      31204: inst = 32'h10408000;
      31205: inst = 32'hc404526;
      31206: inst = 32'h8220000;
      31207: inst = 32'h10408000;
      31208: inst = 32'hc404527;
      31209: inst = 32'h8220000;
      31210: inst = 32'h10408000;
      31211: inst = 32'hc404528;
      31212: inst = 32'h8220000;
      31213: inst = 32'h10408000;
      31214: inst = 32'hc404529;
      31215: inst = 32'h8220000;
      31216: inst = 32'h10408000;
      31217: inst = 32'hc40452a;
      31218: inst = 32'h8220000;
      31219: inst = 32'h10408000;
      31220: inst = 32'hc40452b;
      31221: inst = 32'h8220000;
      31222: inst = 32'h10408000;
      31223: inst = 32'hc40452c;
      31224: inst = 32'h8220000;
      31225: inst = 32'h10408000;
      31226: inst = 32'hc40452d;
      31227: inst = 32'h8220000;
      31228: inst = 32'h10408000;
      31229: inst = 32'hc40452e;
      31230: inst = 32'h8220000;
      31231: inst = 32'h10408000;
      31232: inst = 32'hc40452f;
      31233: inst = 32'h8220000;
      31234: inst = 32'h10408000;
      31235: inst = 32'hc404530;
      31236: inst = 32'h8220000;
      31237: inst = 32'h10408000;
      31238: inst = 32'hc404531;
      31239: inst = 32'h8220000;
      31240: inst = 32'h10408000;
      31241: inst = 32'hc404532;
      31242: inst = 32'h8220000;
      31243: inst = 32'h10408000;
      31244: inst = 32'hc404533;
      31245: inst = 32'h8220000;
      31246: inst = 32'h10408000;
      31247: inst = 32'hc404534;
      31248: inst = 32'h8220000;
      31249: inst = 32'h10408000;
      31250: inst = 32'hc404535;
      31251: inst = 32'h8220000;
      31252: inst = 32'h10408000;
      31253: inst = 32'hc404536;
      31254: inst = 32'h8220000;
      31255: inst = 32'h10408000;
      31256: inst = 32'hc404537;
      31257: inst = 32'h8220000;
      31258: inst = 32'h10408000;
      31259: inst = 32'hc404538;
      31260: inst = 32'h8220000;
      31261: inst = 32'h10408000;
      31262: inst = 32'hc404539;
      31263: inst = 32'h8220000;
      31264: inst = 32'h10408000;
      31265: inst = 32'hc40453a;
      31266: inst = 32'h8220000;
      31267: inst = 32'h10408000;
      31268: inst = 32'hc40453b;
      31269: inst = 32'h8220000;
      31270: inst = 32'h10408000;
      31271: inst = 32'hc40453c;
      31272: inst = 32'h8220000;
      31273: inst = 32'h10408000;
      31274: inst = 32'hc40453d;
      31275: inst = 32'h8220000;
      31276: inst = 32'h10408000;
      31277: inst = 32'hc40453e;
      31278: inst = 32'h8220000;
      31279: inst = 32'h10408000;
      31280: inst = 32'hc40453f;
      31281: inst = 32'h8220000;
      31282: inst = 32'h10408000;
      31283: inst = 32'hc404540;
      31284: inst = 32'h8220000;
      31285: inst = 32'h10408000;
      31286: inst = 32'hc404541;
      31287: inst = 32'h8220000;
      31288: inst = 32'h10408000;
      31289: inst = 32'hc404542;
      31290: inst = 32'h8220000;
      31291: inst = 32'h10408000;
      31292: inst = 32'hc404543;
      31293: inst = 32'h8220000;
      31294: inst = 32'h10408000;
      31295: inst = 32'hc404544;
      31296: inst = 32'h8220000;
      31297: inst = 32'h10408000;
      31298: inst = 32'hc404545;
      31299: inst = 32'h8220000;
      31300: inst = 32'h10408000;
      31301: inst = 32'hc404546;
      31302: inst = 32'h8220000;
      31303: inst = 32'h10408000;
      31304: inst = 32'hc404547;
      31305: inst = 32'h8220000;
      31306: inst = 32'h10408000;
      31307: inst = 32'hc404548;
      31308: inst = 32'h8220000;
      31309: inst = 32'h10408000;
      31310: inst = 32'hc404549;
      31311: inst = 32'h8220000;
      31312: inst = 32'h10408000;
      31313: inst = 32'hc40454a;
      31314: inst = 32'h8220000;
      31315: inst = 32'h10408000;
      31316: inst = 32'hc40454b;
      31317: inst = 32'h8220000;
      31318: inst = 32'h10408000;
      31319: inst = 32'hc40454c;
      31320: inst = 32'h8220000;
      31321: inst = 32'h10408000;
      31322: inst = 32'hc40454d;
      31323: inst = 32'h8220000;
      31324: inst = 32'h10408000;
      31325: inst = 32'hc40454e;
      31326: inst = 32'h8220000;
      31327: inst = 32'h10408000;
      31328: inst = 32'hc40454f;
      31329: inst = 32'h8220000;
      31330: inst = 32'h10408000;
      31331: inst = 32'hc404550;
      31332: inst = 32'h8220000;
      31333: inst = 32'h10408000;
      31334: inst = 32'hc404551;
      31335: inst = 32'h8220000;
      31336: inst = 32'h10408000;
      31337: inst = 32'hc404552;
      31338: inst = 32'h8220000;
      31339: inst = 32'h10408000;
      31340: inst = 32'hc404553;
      31341: inst = 32'h8220000;
      31342: inst = 32'h10408000;
      31343: inst = 32'hc404554;
      31344: inst = 32'h8220000;
      31345: inst = 32'h10408000;
      31346: inst = 32'hc404555;
      31347: inst = 32'h8220000;
      31348: inst = 32'h10408000;
      31349: inst = 32'hc404556;
      31350: inst = 32'h8220000;
      31351: inst = 32'h10408000;
      31352: inst = 32'hc404557;
      31353: inst = 32'h8220000;
      31354: inst = 32'h10408000;
      31355: inst = 32'hc404558;
      31356: inst = 32'h8220000;
      31357: inst = 32'h10408000;
      31358: inst = 32'hc404559;
      31359: inst = 32'h8220000;
      31360: inst = 32'h10408000;
      31361: inst = 32'hc40455a;
      31362: inst = 32'h8220000;
      31363: inst = 32'h10408000;
      31364: inst = 32'hc40455b;
      31365: inst = 32'h8220000;
      31366: inst = 32'h10408000;
      31367: inst = 32'hc40455c;
      31368: inst = 32'h8220000;
      31369: inst = 32'h10408000;
      31370: inst = 32'hc40455d;
      31371: inst = 32'h8220000;
      31372: inst = 32'h10408000;
      31373: inst = 32'hc40455e;
      31374: inst = 32'h8220000;
      31375: inst = 32'h10408000;
      31376: inst = 32'hc40455f;
      31377: inst = 32'h8220000;
      31378: inst = 32'h10408000;
      31379: inst = 32'hc404560;
      31380: inst = 32'h8220000;
      31381: inst = 32'h10408000;
      31382: inst = 32'hc404561;
      31383: inst = 32'h8220000;
      31384: inst = 32'h10408000;
      31385: inst = 32'hc404562;
      31386: inst = 32'h8220000;
      31387: inst = 32'h10408000;
      31388: inst = 32'hc404563;
      31389: inst = 32'h8220000;
      31390: inst = 32'h10408000;
      31391: inst = 32'hc404564;
      31392: inst = 32'h8220000;
      31393: inst = 32'h10408000;
      31394: inst = 32'hc404565;
      31395: inst = 32'h8220000;
      31396: inst = 32'h10408000;
      31397: inst = 32'hc404566;
      31398: inst = 32'h8220000;
      31399: inst = 32'h10408000;
      31400: inst = 32'hc404567;
      31401: inst = 32'h8220000;
      31402: inst = 32'h10408000;
      31403: inst = 32'hc404568;
      31404: inst = 32'h8220000;
      31405: inst = 32'h10408000;
      31406: inst = 32'hc404569;
      31407: inst = 32'h8220000;
      31408: inst = 32'h10408000;
      31409: inst = 32'hc40456a;
      31410: inst = 32'h8220000;
      31411: inst = 32'h10408000;
      31412: inst = 32'hc40456b;
      31413: inst = 32'h8220000;
      31414: inst = 32'h10408000;
      31415: inst = 32'hc40456f;
      31416: inst = 32'h8220000;
      31417: inst = 32'h10408000;
      31418: inst = 32'hc40457a;
      31419: inst = 32'h8220000;
      31420: inst = 32'h10408000;
      31421: inst = 32'hc40457b;
      31422: inst = 32'h8220000;
      31423: inst = 32'h10408000;
      31424: inst = 32'hc40457c;
      31425: inst = 32'h8220000;
      31426: inst = 32'h10408000;
      31427: inst = 32'hc404583;
      31428: inst = 32'h8220000;
      31429: inst = 32'h10408000;
      31430: inst = 32'hc404584;
      31431: inst = 32'h8220000;
      31432: inst = 32'h10408000;
      31433: inst = 32'hc404585;
      31434: inst = 32'h8220000;
      31435: inst = 32'h10408000;
      31436: inst = 32'hc404586;
      31437: inst = 32'h8220000;
      31438: inst = 32'h10408000;
      31439: inst = 32'hc404587;
      31440: inst = 32'h8220000;
      31441: inst = 32'h10408000;
      31442: inst = 32'hc404588;
      31443: inst = 32'h8220000;
      31444: inst = 32'h10408000;
      31445: inst = 32'hc404589;
      31446: inst = 32'h8220000;
      31447: inst = 32'h10408000;
      31448: inst = 32'hc40458a;
      31449: inst = 32'h8220000;
      31450: inst = 32'h10408000;
      31451: inst = 32'hc40458b;
      31452: inst = 32'h8220000;
      31453: inst = 32'h10408000;
      31454: inst = 32'hc40458c;
      31455: inst = 32'h8220000;
      31456: inst = 32'h10408000;
      31457: inst = 32'hc40458d;
      31458: inst = 32'h8220000;
      31459: inst = 32'h10408000;
      31460: inst = 32'hc40458e;
      31461: inst = 32'h8220000;
      31462: inst = 32'h10408000;
      31463: inst = 32'hc40458f;
      31464: inst = 32'h8220000;
      31465: inst = 32'h10408000;
      31466: inst = 32'hc404590;
      31467: inst = 32'h8220000;
      31468: inst = 32'h10408000;
      31469: inst = 32'hc404591;
      31470: inst = 32'h8220000;
      31471: inst = 32'h10408000;
      31472: inst = 32'hc404592;
      31473: inst = 32'h8220000;
      31474: inst = 32'h10408000;
      31475: inst = 32'hc404593;
      31476: inst = 32'h8220000;
      31477: inst = 32'h10408000;
      31478: inst = 32'hc404594;
      31479: inst = 32'h8220000;
      31480: inst = 32'h10408000;
      31481: inst = 32'hc404595;
      31482: inst = 32'h8220000;
      31483: inst = 32'h10408000;
      31484: inst = 32'hc404596;
      31485: inst = 32'h8220000;
      31486: inst = 32'h10408000;
      31487: inst = 32'hc404597;
      31488: inst = 32'h8220000;
      31489: inst = 32'h10408000;
      31490: inst = 32'hc404598;
      31491: inst = 32'h8220000;
      31492: inst = 32'h10408000;
      31493: inst = 32'hc404599;
      31494: inst = 32'h8220000;
      31495: inst = 32'h10408000;
      31496: inst = 32'hc40459a;
      31497: inst = 32'h8220000;
      31498: inst = 32'h10408000;
      31499: inst = 32'hc40459b;
      31500: inst = 32'h8220000;
      31501: inst = 32'h10408000;
      31502: inst = 32'hc40459c;
      31503: inst = 32'h8220000;
      31504: inst = 32'h10408000;
      31505: inst = 32'hc40459d;
      31506: inst = 32'h8220000;
      31507: inst = 32'h10408000;
      31508: inst = 32'hc40459e;
      31509: inst = 32'h8220000;
      31510: inst = 32'h10408000;
      31511: inst = 32'hc40459f;
      31512: inst = 32'h8220000;
      31513: inst = 32'h10408000;
      31514: inst = 32'hc4045a0;
      31515: inst = 32'h8220000;
      31516: inst = 32'h10408000;
      31517: inst = 32'hc4045a1;
      31518: inst = 32'h8220000;
      31519: inst = 32'h10408000;
      31520: inst = 32'hc4045a2;
      31521: inst = 32'h8220000;
      31522: inst = 32'h10408000;
      31523: inst = 32'hc4045a3;
      31524: inst = 32'h8220000;
      31525: inst = 32'h10408000;
      31526: inst = 32'hc4045a4;
      31527: inst = 32'h8220000;
      31528: inst = 32'h10408000;
      31529: inst = 32'hc4045a5;
      31530: inst = 32'h8220000;
      31531: inst = 32'h10408000;
      31532: inst = 32'hc4045a6;
      31533: inst = 32'h8220000;
      31534: inst = 32'h10408000;
      31535: inst = 32'hc4045a7;
      31536: inst = 32'h8220000;
      31537: inst = 32'h10408000;
      31538: inst = 32'hc4045a8;
      31539: inst = 32'h8220000;
      31540: inst = 32'h10408000;
      31541: inst = 32'hc4045a9;
      31542: inst = 32'h8220000;
      31543: inst = 32'h10408000;
      31544: inst = 32'hc4045aa;
      31545: inst = 32'h8220000;
      31546: inst = 32'h10408000;
      31547: inst = 32'hc4045ab;
      31548: inst = 32'h8220000;
      31549: inst = 32'h10408000;
      31550: inst = 32'hc4045ac;
      31551: inst = 32'h8220000;
      31552: inst = 32'h10408000;
      31553: inst = 32'hc4045ad;
      31554: inst = 32'h8220000;
      31555: inst = 32'h10408000;
      31556: inst = 32'hc4045ae;
      31557: inst = 32'h8220000;
      31558: inst = 32'h10408000;
      31559: inst = 32'hc4045af;
      31560: inst = 32'h8220000;
      31561: inst = 32'h10408000;
      31562: inst = 32'hc4045b0;
      31563: inst = 32'h8220000;
      31564: inst = 32'h10408000;
      31565: inst = 32'hc4045b1;
      31566: inst = 32'h8220000;
      31567: inst = 32'h10408000;
      31568: inst = 32'hc4045b2;
      31569: inst = 32'h8220000;
      31570: inst = 32'h10408000;
      31571: inst = 32'hc4045b3;
      31572: inst = 32'h8220000;
      31573: inst = 32'h10408000;
      31574: inst = 32'hc4045b4;
      31575: inst = 32'h8220000;
      31576: inst = 32'h10408000;
      31577: inst = 32'hc4045b5;
      31578: inst = 32'h8220000;
      31579: inst = 32'h10408000;
      31580: inst = 32'hc4045b6;
      31581: inst = 32'h8220000;
      31582: inst = 32'h10408000;
      31583: inst = 32'hc4045b7;
      31584: inst = 32'h8220000;
      31585: inst = 32'h10408000;
      31586: inst = 32'hc4045b8;
      31587: inst = 32'h8220000;
      31588: inst = 32'h10408000;
      31589: inst = 32'hc4045b9;
      31590: inst = 32'h8220000;
      31591: inst = 32'h10408000;
      31592: inst = 32'hc4045ba;
      31593: inst = 32'h8220000;
      31594: inst = 32'h10408000;
      31595: inst = 32'hc4045bb;
      31596: inst = 32'h8220000;
      31597: inst = 32'h10408000;
      31598: inst = 32'hc4045bc;
      31599: inst = 32'h8220000;
      31600: inst = 32'h10408000;
      31601: inst = 32'hc4045bd;
      31602: inst = 32'h8220000;
      31603: inst = 32'h10408000;
      31604: inst = 32'hc4045be;
      31605: inst = 32'h8220000;
      31606: inst = 32'h10408000;
      31607: inst = 32'hc4045bf;
      31608: inst = 32'h8220000;
      31609: inst = 32'h10408000;
      31610: inst = 32'hc4045c0;
      31611: inst = 32'h8220000;
      31612: inst = 32'h10408000;
      31613: inst = 32'hc4045c1;
      31614: inst = 32'h8220000;
      31615: inst = 32'h10408000;
      31616: inst = 32'hc4045c2;
      31617: inst = 32'h8220000;
      31618: inst = 32'h10408000;
      31619: inst = 32'hc4045c3;
      31620: inst = 32'h8220000;
      31621: inst = 32'h10408000;
      31622: inst = 32'hc4045c4;
      31623: inst = 32'h8220000;
      31624: inst = 32'h10408000;
      31625: inst = 32'hc4045c5;
      31626: inst = 32'h8220000;
      31627: inst = 32'h10408000;
      31628: inst = 32'hc4045c6;
      31629: inst = 32'h8220000;
      31630: inst = 32'h10408000;
      31631: inst = 32'hc4045c7;
      31632: inst = 32'h8220000;
      31633: inst = 32'h10408000;
      31634: inst = 32'hc4045c8;
      31635: inst = 32'h8220000;
      31636: inst = 32'h10408000;
      31637: inst = 32'hc4045c9;
      31638: inst = 32'h8220000;
      31639: inst = 32'h10408000;
      31640: inst = 32'hc4045ca;
      31641: inst = 32'h8220000;
      31642: inst = 32'h10408000;
      31643: inst = 32'hc4045cb;
      31644: inst = 32'h8220000;
      31645: inst = 32'h10408000;
      31646: inst = 32'hc4045cf;
      31647: inst = 32'h8220000;
      31648: inst = 32'h10408000;
      31649: inst = 32'hc4045d0;
      31650: inst = 32'h8220000;
      31651: inst = 32'h10408000;
      31652: inst = 32'hc4045d4;
      31653: inst = 32'h8220000;
      31654: inst = 32'h10408000;
      31655: inst = 32'hc4045d5;
      31656: inst = 32'h8220000;
      31657: inst = 32'h10408000;
      31658: inst = 32'hc4045d6;
      31659: inst = 32'h8220000;
      31660: inst = 32'h10408000;
      31661: inst = 32'hc4045d7;
      31662: inst = 32'h8220000;
      31663: inst = 32'h10408000;
      31664: inst = 32'hc4045da;
      31665: inst = 32'h8220000;
      31666: inst = 32'h10408000;
      31667: inst = 32'hc4045db;
      31668: inst = 32'h8220000;
      31669: inst = 32'h10408000;
      31670: inst = 32'hc4045e3;
      31671: inst = 32'h8220000;
      31672: inst = 32'h10408000;
      31673: inst = 32'hc4045e4;
      31674: inst = 32'h8220000;
      31675: inst = 32'h10408000;
      31676: inst = 32'hc4045e5;
      31677: inst = 32'h8220000;
      31678: inst = 32'h10408000;
      31679: inst = 32'hc4045e6;
      31680: inst = 32'h8220000;
      31681: inst = 32'h10408000;
      31682: inst = 32'hc4045e7;
      31683: inst = 32'h8220000;
      31684: inst = 32'h10408000;
      31685: inst = 32'hc4045e8;
      31686: inst = 32'h8220000;
      31687: inst = 32'h10408000;
      31688: inst = 32'hc4045e9;
      31689: inst = 32'h8220000;
      31690: inst = 32'h10408000;
      31691: inst = 32'hc4045ea;
      31692: inst = 32'h8220000;
      31693: inst = 32'h10408000;
      31694: inst = 32'hc4045eb;
      31695: inst = 32'h8220000;
      31696: inst = 32'h10408000;
      31697: inst = 32'hc4045ec;
      31698: inst = 32'h8220000;
      31699: inst = 32'h10408000;
      31700: inst = 32'hc4045ed;
      31701: inst = 32'h8220000;
      31702: inst = 32'h10408000;
      31703: inst = 32'hc4045ee;
      31704: inst = 32'h8220000;
      31705: inst = 32'h10408000;
      31706: inst = 32'hc4045ef;
      31707: inst = 32'h8220000;
      31708: inst = 32'h10408000;
      31709: inst = 32'hc4045f0;
      31710: inst = 32'h8220000;
      31711: inst = 32'h10408000;
      31712: inst = 32'hc4045f1;
      31713: inst = 32'h8220000;
      31714: inst = 32'h10408000;
      31715: inst = 32'hc4045f2;
      31716: inst = 32'h8220000;
      31717: inst = 32'h10408000;
      31718: inst = 32'hc4045f3;
      31719: inst = 32'h8220000;
      31720: inst = 32'h10408000;
      31721: inst = 32'hc4045f4;
      31722: inst = 32'h8220000;
      31723: inst = 32'h10408000;
      31724: inst = 32'hc4045f5;
      31725: inst = 32'h8220000;
      31726: inst = 32'h10408000;
      31727: inst = 32'hc4045f6;
      31728: inst = 32'h8220000;
      31729: inst = 32'h10408000;
      31730: inst = 32'hc4045f7;
      31731: inst = 32'h8220000;
      31732: inst = 32'h10408000;
      31733: inst = 32'hc4045f8;
      31734: inst = 32'h8220000;
      31735: inst = 32'h10408000;
      31736: inst = 32'hc4045f9;
      31737: inst = 32'h8220000;
      31738: inst = 32'h10408000;
      31739: inst = 32'hc4045fa;
      31740: inst = 32'h8220000;
      31741: inst = 32'h10408000;
      31742: inst = 32'hc4045fb;
      31743: inst = 32'h8220000;
      31744: inst = 32'h10408000;
      31745: inst = 32'hc4045fc;
      31746: inst = 32'h8220000;
      31747: inst = 32'h10408000;
      31748: inst = 32'hc4045fd;
      31749: inst = 32'h8220000;
      31750: inst = 32'h10408000;
      31751: inst = 32'hc4045fe;
      31752: inst = 32'h8220000;
      31753: inst = 32'h10408000;
      31754: inst = 32'hc4045ff;
      31755: inst = 32'h8220000;
      31756: inst = 32'h10408000;
      31757: inst = 32'hc404600;
      31758: inst = 32'h8220000;
      31759: inst = 32'h10408000;
      31760: inst = 32'hc404601;
      31761: inst = 32'h8220000;
      31762: inst = 32'h10408000;
      31763: inst = 32'hc404602;
      31764: inst = 32'h8220000;
      31765: inst = 32'h10408000;
      31766: inst = 32'hc404603;
      31767: inst = 32'h8220000;
      31768: inst = 32'h10408000;
      31769: inst = 32'hc404604;
      31770: inst = 32'h8220000;
      31771: inst = 32'h10408000;
      31772: inst = 32'hc404605;
      31773: inst = 32'h8220000;
      31774: inst = 32'h10408000;
      31775: inst = 32'hc404606;
      31776: inst = 32'h8220000;
      31777: inst = 32'h10408000;
      31778: inst = 32'hc404607;
      31779: inst = 32'h8220000;
      31780: inst = 32'h10408000;
      31781: inst = 32'hc404608;
      31782: inst = 32'h8220000;
      31783: inst = 32'h10408000;
      31784: inst = 32'hc404609;
      31785: inst = 32'h8220000;
      31786: inst = 32'h10408000;
      31787: inst = 32'hc40460a;
      31788: inst = 32'h8220000;
      31789: inst = 32'h10408000;
      31790: inst = 32'hc40460b;
      31791: inst = 32'h8220000;
      31792: inst = 32'h10408000;
      31793: inst = 32'hc40460c;
      31794: inst = 32'h8220000;
      31795: inst = 32'h10408000;
      31796: inst = 32'hc40460d;
      31797: inst = 32'h8220000;
      31798: inst = 32'h10408000;
      31799: inst = 32'hc40460e;
      31800: inst = 32'h8220000;
      31801: inst = 32'h10408000;
      31802: inst = 32'hc40460f;
      31803: inst = 32'h8220000;
      31804: inst = 32'h10408000;
      31805: inst = 32'hc404610;
      31806: inst = 32'h8220000;
      31807: inst = 32'h10408000;
      31808: inst = 32'hc404611;
      31809: inst = 32'h8220000;
      31810: inst = 32'h10408000;
      31811: inst = 32'hc404612;
      31812: inst = 32'h8220000;
      31813: inst = 32'h10408000;
      31814: inst = 32'hc404613;
      31815: inst = 32'h8220000;
      31816: inst = 32'h10408000;
      31817: inst = 32'hc404614;
      31818: inst = 32'h8220000;
      31819: inst = 32'h10408000;
      31820: inst = 32'hc404615;
      31821: inst = 32'h8220000;
      31822: inst = 32'h10408000;
      31823: inst = 32'hc404616;
      31824: inst = 32'h8220000;
      31825: inst = 32'h10408000;
      31826: inst = 32'hc404617;
      31827: inst = 32'h8220000;
      31828: inst = 32'h10408000;
      31829: inst = 32'hc404618;
      31830: inst = 32'h8220000;
      31831: inst = 32'h10408000;
      31832: inst = 32'hc404619;
      31833: inst = 32'h8220000;
      31834: inst = 32'h10408000;
      31835: inst = 32'hc40461a;
      31836: inst = 32'h8220000;
      31837: inst = 32'h10408000;
      31838: inst = 32'hc40461b;
      31839: inst = 32'h8220000;
      31840: inst = 32'h10408000;
      31841: inst = 32'hc40461c;
      31842: inst = 32'h8220000;
      31843: inst = 32'h10408000;
      31844: inst = 32'hc40461d;
      31845: inst = 32'h8220000;
      31846: inst = 32'h10408000;
      31847: inst = 32'hc40461e;
      31848: inst = 32'h8220000;
      31849: inst = 32'h10408000;
      31850: inst = 32'hc40461f;
      31851: inst = 32'h8220000;
      31852: inst = 32'h10408000;
      31853: inst = 32'hc404620;
      31854: inst = 32'h8220000;
      31855: inst = 32'h10408000;
      31856: inst = 32'hc404621;
      31857: inst = 32'h8220000;
      31858: inst = 32'h10408000;
      31859: inst = 32'hc404622;
      31860: inst = 32'h8220000;
      31861: inst = 32'h10408000;
      31862: inst = 32'hc404623;
      31863: inst = 32'h8220000;
      31864: inst = 32'h10408000;
      31865: inst = 32'hc404624;
      31866: inst = 32'h8220000;
      31867: inst = 32'h10408000;
      31868: inst = 32'hc404625;
      31869: inst = 32'h8220000;
      31870: inst = 32'h10408000;
      31871: inst = 32'hc404626;
      31872: inst = 32'h8220000;
      31873: inst = 32'h10408000;
      31874: inst = 32'hc404627;
      31875: inst = 32'h8220000;
      31876: inst = 32'h10408000;
      31877: inst = 32'hc404628;
      31878: inst = 32'h8220000;
      31879: inst = 32'h10408000;
      31880: inst = 32'hc404629;
      31881: inst = 32'h8220000;
      31882: inst = 32'h10408000;
      31883: inst = 32'hc40462a;
      31884: inst = 32'h8220000;
      31885: inst = 32'h10408000;
      31886: inst = 32'hc40462b;
      31887: inst = 32'h8220000;
      31888: inst = 32'h10408000;
      31889: inst = 32'hc40462f;
      31890: inst = 32'h8220000;
      31891: inst = 32'h10408000;
      31892: inst = 32'hc404630;
      31893: inst = 32'h8220000;
      31894: inst = 32'h10408000;
      31895: inst = 32'hc404631;
      31896: inst = 32'h8220000;
      31897: inst = 32'h10408000;
      31898: inst = 32'hc404632;
      31899: inst = 32'h8220000;
      31900: inst = 32'h10408000;
      31901: inst = 32'hc404633;
      31902: inst = 32'h8220000;
      31903: inst = 32'h10408000;
      31904: inst = 32'hc404634;
      31905: inst = 32'h8220000;
      31906: inst = 32'h10408000;
      31907: inst = 32'hc404635;
      31908: inst = 32'h8220000;
      31909: inst = 32'h10408000;
      31910: inst = 32'hc404636;
      31911: inst = 32'h8220000;
      31912: inst = 32'h10408000;
      31913: inst = 32'hc404637;
      31914: inst = 32'h8220000;
      31915: inst = 32'h10408000;
      31916: inst = 32'hc404638;
      31917: inst = 32'h8220000;
      31918: inst = 32'h10408000;
      31919: inst = 32'hc404639;
      31920: inst = 32'h8220000;
      31921: inst = 32'h10408000;
      31922: inst = 32'hc40463a;
      31923: inst = 32'h8220000;
      31924: inst = 32'h10408000;
      31925: inst = 32'hc40463b;
      31926: inst = 32'h8220000;
      31927: inst = 32'h10408000;
      31928: inst = 32'hc40463c;
      31929: inst = 32'h8220000;
      31930: inst = 32'h10408000;
      31931: inst = 32'hc404643;
      31932: inst = 32'h8220000;
      31933: inst = 32'h10408000;
      31934: inst = 32'hc404644;
      31935: inst = 32'h8220000;
      31936: inst = 32'h10408000;
      31937: inst = 32'hc404645;
      31938: inst = 32'h8220000;
      31939: inst = 32'h10408000;
      31940: inst = 32'hc404646;
      31941: inst = 32'h8220000;
      31942: inst = 32'h10408000;
      31943: inst = 32'hc404647;
      31944: inst = 32'h8220000;
      31945: inst = 32'h10408000;
      31946: inst = 32'hc404648;
      31947: inst = 32'h8220000;
      31948: inst = 32'h10408000;
      31949: inst = 32'hc404649;
      31950: inst = 32'h8220000;
      31951: inst = 32'h10408000;
      31952: inst = 32'hc40464a;
      31953: inst = 32'h8220000;
      31954: inst = 32'h10408000;
      31955: inst = 32'hc40464b;
      31956: inst = 32'h8220000;
      31957: inst = 32'h10408000;
      31958: inst = 32'hc40464c;
      31959: inst = 32'h8220000;
      31960: inst = 32'h10408000;
      31961: inst = 32'hc40464d;
      31962: inst = 32'h8220000;
      31963: inst = 32'h10408000;
      31964: inst = 32'hc40467a;
      31965: inst = 32'h8220000;
      31966: inst = 32'h10408000;
      31967: inst = 32'hc40467b;
      31968: inst = 32'h8220000;
      31969: inst = 32'h10408000;
      31970: inst = 32'hc40467c;
      31971: inst = 32'h8220000;
      31972: inst = 32'h10408000;
      31973: inst = 32'hc40467d;
      31974: inst = 32'h8220000;
      31975: inst = 32'h10408000;
      31976: inst = 32'hc40467e;
      31977: inst = 32'h8220000;
      31978: inst = 32'h10408000;
      31979: inst = 32'hc40467f;
      31980: inst = 32'h8220000;
      31981: inst = 32'h10408000;
      31982: inst = 32'hc404680;
      31983: inst = 32'h8220000;
      31984: inst = 32'h10408000;
      31985: inst = 32'hc404681;
      31986: inst = 32'h8220000;
      31987: inst = 32'h10408000;
      31988: inst = 32'hc404682;
      31989: inst = 32'h8220000;
      31990: inst = 32'h10408000;
      31991: inst = 32'hc404683;
      31992: inst = 32'h8220000;
      31993: inst = 32'h10408000;
      31994: inst = 32'hc404684;
      31995: inst = 32'h8220000;
      31996: inst = 32'h10408000;
      31997: inst = 32'hc404685;
      31998: inst = 32'h8220000;
      31999: inst = 32'h10408000;
      32000: inst = 32'hc404686;
      32001: inst = 32'h8220000;
      32002: inst = 32'h10408000;
      32003: inst = 32'hc404687;
      32004: inst = 32'h8220000;
      32005: inst = 32'h10408000;
      32006: inst = 32'hc404688;
      32007: inst = 32'h8220000;
      32008: inst = 32'h10408000;
      32009: inst = 32'hc404689;
      32010: inst = 32'h8220000;
      32011: inst = 32'h10408000;
      32012: inst = 32'hc40468a;
      32013: inst = 32'h8220000;
      32014: inst = 32'h10408000;
      32015: inst = 32'hc40468b;
      32016: inst = 32'h8220000;
      32017: inst = 32'h10408000;
      32018: inst = 32'hc40468f;
      32019: inst = 32'h8220000;
      32020: inst = 32'h10408000;
      32021: inst = 32'hc404690;
      32022: inst = 32'h8220000;
      32023: inst = 32'h10408000;
      32024: inst = 32'hc404691;
      32025: inst = 32'h8220000;
      32026: inst = 32'h10408000;
      32027: inst = 32'hc404692;
      32028: inst = 32'h8220000;
      32029: inst = 32'h10408000;
      32030: inst = 32'hc404693;
      32031: inst = 32'h8220000;
      32032: inst = 32'h10408000;
      32033: inst = 32'hc404694;
      32034: inst = 32'h8220000;
      32035: inst = 32'h10408000;
      32036: inst = 32'hc404695;
      32037: inst = 32'h8220000;
      32038: inst = 32'h10408000;
      32039: inst = 32'hc404696;
      32040: inst = 32'h8220000;
      32041: inst = 32'h10408000;
      32042: inst = 32'hc404697;
      32043: inst = 32'h8220000;
      32044: inst = 32'h10408000;
      32045: inst = 32'hc404698;
      32046: inst = 32'h8220000;
      32047: inst = 32'h10408000;
      32048: inst = 32'hc404699;
      32049: inst = 32'h8220000;
      32050: inst = 32'h10408000;
      32051: inst = 32'hc40469a;
      32052: inst = 32'h8220000;
      32053: inst = 32'h10408000;
      32054: inst = 32'hc40469b;
      32055: inst = 32'h8220000;
      32056: inst = 32'h10408000;
      32057: inst = 32'hc40469c;
      32058: inst = 32'h8220000;
      32059: inst = 32'h10408000;
      32060: inst = 32'hc4046a3;
      32061: inst = 32'h8220000;
      32062: inst = 32'h10408000;
      32063: inst = 32'hc4046a4;
      32064: inst = 32'h8220000;
      32065: inst = 32'h10408000;
      32066: inst = 32'hc4046a5;
      32067: inst = 32'h8220000;
      32068: inst = 32'h10408000;
      32069: inst = 32'hc4046a6;
      32070: inst = 32'h8220000;
      32071: inst = 32'h10408000;
      32072: inst = 32'hc4046a7;
      32073: inst = 32'h8220000;
      32074: inst = 32'h10408000;
      32075: inst = 32'hc4046a8;
      32076: inst = 32'h8220000;
      32077: inst = 32'h10408000;
      32078: inst = 32'hc4046a9;
      32079: inst = 32'h8220000;
      32080: inst = 32'h10408000;
      32081: inst = 32'hc4046aa;
      32082: inst = 32'h8220000;
      32083: inst = 32'h10408000;
      32084: inst = 32'hc4046ab;
      32085: inst = 32'h8220000;
      32086: inst = 32'h10408000;
      32087: inst = 32'hc4046ac;
      32088: inst = 32'h8220000;
      32089: inst = 32'h10408000;
      32090: inst = 32'hc4046ad;
      32091: inst = 32'h8220000;
      32092: inst = 32'h10408000;
      32093: inst = 32'hc4046da;
      32094: inst = 32'h8220000;
      32095: inst = 32'h10408000;
      32096: inst = 32'hc4046db;
      32097: inst = 32'h8220000;
      32098: inst = 32'h10408000;
      32099: inst = 32'hc4046dc;
      32100: inst = 32'h8220000;
      32101: inst = 32'h10408000;
      32102: inst = 32'hc4046dd;
      32103: inst = 32'h8220000;
      32104: inst = 32'h10408000;
      32105: inst = 32'hc4046de;
      32106: inst = 32'h8220000;
      32107: inst = 32'h10408000;
      32108: inst = 32'hc4046df;
      32109: inst = 32'h8220000;
      32110: inst = 32'h10408000;
      32111: inst = 32'hc4046e0;
      32112: inst = 32'h8220000;
      32113: inst = 32'h10408000;
      32114: inst = 32'hc4046e1;
      32115: inst = 32'h8220000;
      32116: inst = 32'h10408000;
      32117: inst = 32'hc4046e2;
      32118: inst = 32'h8220000;
      32119: inst = 32'h10408000;
      32120: inst = 32'hc4046e3;
      32121: inst = 32'h8220000;
      32122: inst = 32'h10408000;
      32123: inst = 32'hc4046e4;
      32124: inst = 32'h8220000;
      32125: inst = 32'h10408000;
      32126: inst = 32'hc4046e5;
      32127: inst = 32'h8220000;
      32128: inst = 32'h10408000;
      32129: inst = 32'hc4046e6;
      32130: inst = 32'h8220000;
      32131: inst = 32'h10408000;
      32132: inst = 32'hc4046e7;
      32133: inst = 32'h8220000;
      32134: inst = 32'h10408000;
      32135: inst = 32'hc4046e8;
      32136: inst = 32'h8220000;
      32137: inst = 32'h10408000;
      32138: inst = 32'hc4046e9;
      32139: inst = 32'h8220000;
      32140: inst = 32'h10408000;
      32141: inst = 32'hc4046ea;
      32142: inst = 32'h8220000;
      32143: inst = 32'h10408000;
      32144: inst = 32'hc4046eb;
      32145: inst = 32'h8220000;
      32146: inst = 32'h10408000;
      32147: inst = 32'hc4046ef;
      32148: inst = 32'h8220000;
      32149: inst = 32'h10408000;
      32150: inst = 32'hc4046f0;
      32151: inst = 32'h8220000;
      32152: inst = 32'h10408000;
      32153: inst = 32'hc4046f1;
      32154: inst = 32'h8220000;
      32155: inst = 32'h10408000;
      32156: inst = 32'hc4046f2;
      32157: inst = 32'h8220000;
      32158: inst = 32'h10408000;
      32159: inst = 32'hc4046f3;
      32160: inst = 32'h8220000;
      32161: inst = 32'h10408000;
      32162: inst = 32'hc4046f4;
      32163: inst = 32'h8220000;
      32164: inst = 32'h10408000;
      32165: inst = 32'hc4046f5;
      32166: inst = 32'h8220000;
      32167: inst = 32'h10408000;
      32168: inst = 32'hc4046f6;
      32169: inst = 32'h8220000;
      32170: inst = 32'h10408000;
      32171: inst = 32'hc4046f7;
      32172: inst = 32'h8220000;
      32173: inst = 32'h10408000;
      32174: inst = 32'hc4046f8;
      32175: inst = 32'h8220000;
      32176: inst = 32'h10408000;
      32177: inst = 32'hc4046f9;
      32178: inst = 32'h8220000;
      32179: inst = 32'h10408000;
      32180: inst = 32'hc4046fa;
      32181: inst = 32'h8220000;
      32182: inst = 32'h10408000;
      32183: inst = 32'hc4046fb;
      32184: inst = 32'h8220000;
      32185: inst = 32'h10408000;
      32186: inst = 32'hc4046fc;
      32187: inst = 32'h8220000;
      32188: inst = 32'h10408000;
      32189: inst = 32'hc404703;
      32190: inst = 32'h8220000;
      32191: inst = 32'h10408000;
      32192: inst = 32'hc404704;
      32193: inst = 32'h8220000;
      32194: inst = 32'h10408000;
      32195: inst = 32'hc404705;
      32196: inst = 32'h8220000;
      32197: inst = 32'h10408000;
      32198: inst = 32'hc404706;
      32199: inst = 32'h8220000;
      32200: inst = 32'h10408000;
      32201: inst = 32'hc404707;
      32202: inst = 32'h8220000;
      32203: inst = 32'h10408000;
      32204: inst = 32'hc404708;
      32205: inst = 32'h8220000;
      32206: inst = 32'h10408000;
      32207: inst = 32'hc404709;
      32208: inst = 32'h8220000;
      32209: inst = 32'h10408000;
      32210: inst = 32'hc40470a;
      32211: inst = 32'h8220000;
      32212: inst = 32'h10408000;
      32213: inst = 32'hc40470b;
      32214: inst = 32'h8220000;
      32215: inst = 32'h10408000;
      32216: inst = 32'hc40470c;
      32217: inst = 32'h8220000;
      32218: inst = 32'h10408000;
      32219: inst = 32'hc40470d;
      32220: inst = 32'h8220000;
      32221: inst = 32'h10408000;
      32222: inst = 32'hc40473a;
      32223: inst = 32'h8220000;
      32224: inst = 32'h10408000;
      32225: inst = 32'hc40473b;
      32226: inst = 32'h8220000;
      32227: inst = 32'h10408000;
      32228: inst = 32'hc40473c;
      32229: inst = 32'h8220000;
      32230: inst = 32'h10408000;
      32231: inst = 32'hc40473d;
      32232: inst = 32'h8220000;
      32233: inst = 32'h10408000;
      32234: inst = 32'hc40473e;
      32235: inst = 32'h8220000;
      32236: inst = 32'h10408000;
      32237: inst = 32'hc40473f;
      32238: inst = 32'h8220000;
      32239: inst = 32'h10408000;
      32240: inst = 32'hc404740;
      32241: inst = 32'h8220000;
      32242: inst = 32'h10408000;
      32243: inst = 32'hc404741;
      32244: inst = 32'h8220000;
      32245: inst = 32'h10408000;
      32246: inst = 32'hc404742;
      32247: inst = 32'h8220000;
      32248: inst = 32'h10408000;
      32249: inst = 32'hc404743;
      32250: inst = 32'h8220000;
      32251: inst = 32'h10408000;
      32252: inst = 32'hc404744;
      32253: inst = 32'h8220000;
      32254: inst = 32'h10408000;
      32255: inst = 32'hc404745;
      32256: inst = 32'h8220000;
      32257: inst = 32'h10408000;
      32258: inst = 32'hc404746;
      32259: inst = 32'h8220000;
      32260: inst = 32'h10408000;
      32261: inst = 32'hc404747;
      32262: inst = 32'h8220000;
      32263: inst = 32'h10408000;
      32264: inst = 32'hc404748;
      32265: inst = 32'h8220000;
      32266: inst = 32'h10408000;
      32267: inst = 32'hc404749;
      32268: inst = 32'h8220000;
      32269: inst = 32'h10408000;
      32270: inst = 32'hc40474a;
      32271: inst = 32'h8220000;
      32272: inst = 32'h10408000;
      32273: inst = 32'hc40474b;
      32274: inst = 32'h8220000;
      32275: inst = 32'h10408000;
      32276: inst = 32'hc40474f;
      32277: inst = 32'h8220000;
      32278: inst = 32'h10408000;
      32279: inst = 32'hc404750;
      32280: inst = 32'h8220000;
      32281: inst = 32'h10408000;
      32282: inst = 32'hc404751;
      32283: inst = 32'h8220000;
      32284: inst = 32'h10408000;
      32285: inst = 32'hc404752;
      32286: inst = 32'h8220000;
      32287: inst = 32'h10408000;
      32288: inst = 32'hc404753;
      32289: inst = 32'h8220000;
      32290: inst = 32'h10408000;
      32291: inst = 32'hc404754;
      32292: inst = 32'h8220000;
      32293: inst = 32'h10408000;
      32294: inst = 32'hc404755;
      32295: inst = 32'h8220000;
      32296: inst = 32'h10408000;
      32297: inst = 32'hc404756;
      32298: inst = 32'h8220000;
      32299: inst = 32'h10408000;
      32300: inst = 32'hc404757;
      32301: inst = 32'h8220000;
      32302: inst = 32'h10408000;
      32303: inst = 32'hc404758;
      32304: inst = 32'h8220000;
      32305: inst = 32'h10408000;
      32306: inst = 32'hc404759;
      32307: inst = 32'h8220000;
      32308: inst = 32'h10408000;
      32309: inst = 32'hc40475a;
      32310: inst = 32'h8220000;
      32311: inst = 32'h10408000;
      32312: inst = 32'hc40475b;
      32313: inst = 32'h8220000;
      32314: inst = 32'h10408000;
      32315: inst = 32'hc40475c;
      32316: inst = 32'h8220000;
      32317: inst = 32'h10408000;
      32318: inst = 32'hc404763;
      32319: inst = 32'h8220000;
      32320: inst = 32'h10408000;
      32321: inst = 32'hc404764;
      32322: inst = 32'h8220000;
      32323: inst = 32'h10408000;
      32324: inst = 32'hc404765;
      32325: inst = 32'h8220000;
      32326: inst = 32'h10408000;
      32327: inst = 32'hc404766;
      32328: inst = 32'h8220000;
      32329: inst = 32'h10408000;
      32330: inst = 32'hc404767;
      32331: inst = 32'h8220000;
      32332: inst = 32'h10408000;
      32333: inst = 32'hc404768;
      32334: inst = 32'h8220000;
      32335: inst = 32'h10408000;
      32336: inst = 32'hc404769;
      32337: inst = 32'h8220000;
      32338: inst = 32'h10408000;
      32339: inst = 32'hc40476a;
      32340: inst = 32'h8220000;
      32341: inst = 32'h10408000;
      32342: inst = 32'hc40476b;
      32343: inst = 32'h8220000;
      32344: inst = 32'h10408000;
      32345: inst = 32'hc40476c;
      32346: inst = 32'h8220000;
      32347: inst = 32'h10408000;
      32348: inst = 32'hc40476d;
      32349: inst = 32'h8220000;
      32350: inst = 32'h10408000;
      32351: inst = 32'hc404771;
      32352: inst = 32'h8220000;
      32353: inst = 32'h10408000;
      32354: inst = 32'hc404772;
      32355: inst = 32'h8220000;
      32356: inst = 32'h10408000;
      32357: inst = 32'hc404773;
      32358: inst = 32'h8220000;
      32359: inst = 32'h10408000;
      32360: inst = 32'hc404774;
      32361: inst = 32'h8220000;
      32362: inst = 32'h10408000;
      32363: inst = 32'hc404775;
      32364: inst = 32'h8220000;
      32365: inst = 32'h10408000;
      32366: inst = 32'hc404776;
      32367: inst = 32'h8220000;
      32368: inst = 32'h10408000;
      32369: inst = 32'hc404777;
      32370: inst = 32'h8220000;
      32371: inst = 32'h10408000;
      32372: inst = 32'hc404778;
      32373: inst = 32'h8220000;
      32374: inst = 32'h10408000;
      32375: inst = 32'hc404779;
      32376: inst = 32'h8220000;
      32377: inst = 32'h10408000;
      32378: inst = 32'hc40477a;
      32379: inst = 32'h8220000;
      32380: inst = 32'h10408000;
      32381: inst = 32'hc40477b;
      32382: inst = 32'h8220000;
      32383: inst = 32'h10408000;
      32384: inst = 32'hc40477c;
      32385: inst = 32'h8220000;
      32386: inst = 32'h10408000;
      32387: inst = 32'hc40477d;
      32388: inst = 32'h8220000;
      32389: inst = 32'h10408000;
      32390: inst = 32'hc40477e;
      32391: inst = 32'h8220000;
      32392: inst = 32'h10408000;
      32393: inst = 32'hc40477f;
      32394: inst = 32'h8220000;
      32395: inst = 32'h10408000;
      32396: inst = 32'hc404780;
      32397: inst = 32'h8220000;
      32398: inst = 32'h10408000;
      32399: inst = 32'hc404781;
      32400: inst = 32'h8220000;
      32401: inst = 32'h10408000;
      32402: inst = 32'hc404782;
      32403: inst = 32'h8220000;
      32404: inst = 32'h10408000;
      32405: inst = 32'hc404783;
      32406: inst = 32'h8220000;
      32407: inst = 32'h10408000;
      32408: inst = 32'hc404784;
      32409: inst = 32'h8220000;
      32410: inst = 32'h10408000;
      32411: inst = 32'hc404785;
      32412: inst = 32'h8220000;
      32413: inst = 32'h10408000;
      32414: inst = 32'hc404786;
      32415: inst = 32'h8220000;
      32416: inst = 32'h10408000;
      32417: inst = 32'hc404787;
      32418: inst = 32'h8220000;
      32419: inst = 32'h10408000;
      32420: inst = 32'hc404788;
      32421: inst = 32'h8220000;
      32422: inst = 32'h10408000;
      32423: inst = 32'hc404789;
      32424: inst = 32'h8220000;
      32425: inst = 32'h10408000;
      32426: inst = 32'hc40478a;
      32427: inst = 32'h8220000;
      32428: inst = 32'h10408000;
      32429: inst = 32'hc404795;
      32430: inst = 32'h8220000;
      32431: inst = 32'h10408000;
      32432: inst = 32'hc404796;
      32433: inst = 32'h8220000;
      32434: inst = 32'h10408000;
      32435: inst = 32'hc404797;
      32436: inst = 32'h8220000;
      32437: inst = 32'h10408000;
      32438: inst = 32'hc404799;
      32439: inst = 32'h8220000;
      32440: inst = 32'h10408000;
      32441: inst = 32'hc40479a;
      32442: inst = 32'h8220000;
      32443: inst = 32'h10408000;
      32444: inst = 32'hc40479b;
      32445: inst = 32'h8220000;
      32446: inst = 32'h10408000;
      32447: inst = 32'hc40479c;
      32448: inst = 32'h8220000;
      32449: inst = 32'h10408000;
      32450: inst = 32'hc40479d;
      32451: inst = 32'h8220000;
      32452: inst = 32'h10408000;
      32453: inst = 32'hc40479e;
      32454: inst = 32'h8220000;
      32455: inst = 32'h10408000;
      32456: inst = 32'hc40479f;
      32457: inst = 32'h8220000;
      32458: inst = 32'h10408000;
      32459: inst = 32'hc4047a0;
      32460: inst = 32'h8220000;
      32461: inst = 32'h10408000;
      32462: inst = 32'hc4047a1;
      32463: inst = 32'h8220000;
      32464: inst = 32'h10408000;
      32465: inst = 32'hc4047a2;
      32466: inst = 32'h8220000;
      32467: inst = 32'h10408000;
      32468: inst = 32'hc4047a3;
      32469: inst = 32'h8220000;
      32470: inst = 32'h10408000;
      32471: inst = 32'hc4047a4;
      32472: inst = 32'h8220000;
      32473: inst = 32'h10408000;
      32474: inst = 32'hc4047a5;
      32475: inst = 32'h8220000;
      32476: inst = 32'h10408000;
      32477: inst = 32'hc4047a6;
      32478: inst = 32'h8220000;
      32479: inst = 32'h10408000;
      32480: inst = 32'hc4047a7;
      32481: inst = 32'h8220000;
      32482: inst = 32'h10408000;
      32483: inst = 32'hc4047a8;
      32484: inst = 32'h8220000;
      32485: inst = 32'h10408000;
      32486: inst = 32'hc4047a9;
      32487: inst = 32'h8220000;
      32488: inst = 32'h10408000;
      32489: inst = 32'hc4047aa;
      32490: inst = 32'h8220000;
      32491: inst = 32'h10408000;
      32492: inst = 32'hc4047ab;
      32493: inst = 32'h8220000;
      32494: inst = 32'h10408000;
      32495: inst = 32'hc4047af;
      32496: inst = 32'h8220000;
      32497: inst = 32'h10408000;
      32498: inst = 32'hc4047b0;
      32499: inst = 32'h8220000;
      32500: inst = 32'h10408000;
      32501: inst = 32'hc4047b1;
      32502: inst = 32'h8220000;
      32503: inst = 32'h10408000;
      32504: inst = 32'hc4047b2;
      32505: inst = 32'h8220000;
      32506: inst = 32'h10408000;
      32507: inst = 32'hc4047b3;
      32508: inst = 32'h8220000;
      32509: inst = 32'h10408000;
      32510: inst = 32'hc4047b4;
      32511: inst = 32'h8220000;
      32512: inst = 32'h10408000;
      32513: inst = 32'hc4047b5;
      32514: inst = 32'h8220000;
      32515: inst = 32'h10408000;
      32516: inst = 32'hc4047b6;
      32517: inst = 32'h8220000;
      32518: inst = 32'h10408000;
      32519: inst = 32'hc4047b7;
      32520: inst = 32'h8220000;
      32521: inst = 32'h10408000;
      32522: inst = 32'hc4047b8;
      32523: inst = 32'h8220000;
      32524: inst = 32'h10408000;
      32525: inst = 32'hc4047b9;
      32526: inst = 32'h8220000;
      32527: inst = 32'h10408000;
      32528: inst = 32'hc4047ba;
      32529: inst = 32'h8220000;
      32530: inst = 32'h10408000;
      32531: inst = 32'hc4047bb;
      32532: inst = 32'h8220000;
      32533: inst = 32'h10408000;
      32534: inst = 32'hc4047bc;
      32535: inst = 32'h8220000;
      32536: inst = 32'h10408000;
      32537: inst = 32'hc4047c3;
      32538: inst = 32'h8220000;
      32539: inst = 32'h10408000;
      32540: inst = 32'hc4047c4;
      32541: inst = 32'h8220000;
      32542: inst = 32'h10408000;
      32543: inst = 32'hc4047c5;
      32544: inst = 32'h8220000;
      32545: inst = 32'h10408000;
      32546: inst = 32'hc4047c6;
      32547: inst = 32'h8220000;
      32548: inst = 32'h10408000;
      32549: inst = 32'hc4047c7;
      32550: inst = 32'h8220000;
      32551: inst = 32'h10408000;
      32552: inst = 32'hc4047c8;
      32553: inst = 32'h8220000;
      32554: inst = 32'h10408000;
      32555: inst = 32'hc4047c9;
      32556: inst = 32'h8220000;
      32557: inst = 32'h10408000;
      32558: inst = 32'hc4047ca;
      32559: inst = 32'h8220000;
      32560: inst = 32'h10408000;
      32561: inst = 32'hc4047cb;
      32562: inst = 32'h8220000;
      32563: inst = 32'h10408000;
      32564: inst = 32'hc4047cc;
      32565: inst = 32'h8220000;
      32566: inst = 32'h10408000;
      32567: inst = 32'hc4047cd;
      32568: inst = 32'h8220000;
      32569: inst = 32'h10408000;
      32570: inst = 32'hc4047d1;
      32571: inst = 32'h8220000;
      32572: inst = 32'h10408000;
      32573: inst = 32'hc4047d2;
      32574: inst = 32'h8220000;
      32575: inst = 32'h10408000;
      32576: inst = 32'hc4047d3;
      32577: inst = 32'h8220000;
      32578: inst = 32'h10408000;
      32579: inst = 32'hc4047d4;
      32580: inst = 32'h8220000;
      32581: inst = 32'h10408000;
      32582: inst = 32'hc4047d5;
      32583: inst = 32'h8220000;
      32584: inst = 32'h10408000;
      32585: inst = 32'hc4047d6;
      32586: inst = 32'h8220000;
      32587: inst = 32'h10408000;
      32588: inst = 32'hc4047d7;
      32589: inst = 32'h8220000;
      32590: inst = 32'h10408000;
      32591: inst = 32'hc4047d8;
      32592: inst = 32'h8220000;
      32593: inst = 32'h10408000;
      32594: inst = 32'hc4047d9;
      32595: inst = 32'h8220000;
      32596: inst = 32'h10408000;
      32597: inst = 32'hc4047da;
      32598: inst = 32'h8220000;
      32599: inst = 32'h10408000;
      32600: inst = 32'hc4047db;
      32601: inst = 32'h8220000;
      32602: inst = 32'h10408000;
      32603: inst = 32'hc4047dc;
      32604: inst = 32'h8220000;
      32605: inst = 32'h10408000;
      32606: inst = 32'hc4047dd;
      32607: inst = 32'h8220000;
      32608: inst = 32'h10408000;
      32609: inst = 32'hc4047de;
      32610: inst = 32'h8220000;
      32611: inst = 32'h10408000;
      32612: inst = 32'hc4047df;
      32613: inst = 32'h8220000;
      32614: inst = 32'h10408000;
      32615: inst = 32'hc4047e0;
      32616: inst = 32'h8220000;
      32617: inst = 32'h10408000;
      32618: inst = 32'hc4047e1;
      32619: inst = 32'h8220000;
      32620: inst = 32'h10408000;
      32621: inst = 32'hc4047e2;
      32622: inst = 32'h8220000;
      32623: inst = 32'h10408000;
      32624: inst = 32'hc4047e3;
      32625: inst = 32'h8220000;
      32626: inst = 32'h10408000;
      32627: inst = 32'hc4047e4;
      32628: inst = 32'h8220000;
      32629: inst = 32'h10408000;
      32630: inst = 32'hc4047e5;
      32631: inst = 32'h8220000;
      32632: inst = 32'h10408000;
      32633: inst = 32'hc4047e6;
      32634: inst = 32'h8220000;
      32635: inst = 32'h10408000;
      32636: inst = 32'hc4047e7;
      32637: inst = 32'h8220000;
      32638: inst = 32'h10408000;
      32639: inst = 32'hc4047e8;
      32640: inst = 32'h8220000;
      32641: inst = 32'h10408000;
      32642: inst = 32'hc4047e9;
      32643: inst = 32'h8220000;
      32644: inst = 32'h10408000;
      32645: inst = 32'hc4047ea;
      32646: inst = 32'h8220000;
      32647: inst = 32'h10408000;
      32648: inst = 32'hc4047ee;
      32649: inst = 32'h8220000;
      32650: inst = 32'h10408000;
      32651: inst = 32'hc4047ef;
      32652: inst = 32'h8220000;
      32653: inst = 32'h10408000;
      32654: inst = 32'hc4047f6;
      32655: inst = 32'h8220000;
      32656: inst = 32'h10408000;
      32657: inst = 32'hc4047f7;
      32658: inst = 32'h8220000;
      32659: inst = 32'h10408000;
      32660: inst = 32'hc4047fa;
      32661: inst = 32'h8220000;
      32662: inst = 32'h10408000;
      32663: inst = 32'hc4047fb;
      32664: inst = 32'h8220000;
      32665: inst = 32'h10408000;
      32666: inst = 32'hc4047fc;
      32667: inst = 32'h8220000;
      32668: inst = 32'h10408000;
      32669: inst = 32'hc4047fd;
      32670: inst = 32'h8220000;
      32671: inst = 32'h10408000;
      32672: inst = 32'hc4047fe;
      32673: inst = 32'h8220000;
      32674: inst = 32'h10408000;
      32675: inst = 32'hc4047ff;
      32676: inst = 32'h8220000;
      32677: inst = 32'h10408000;
      32678: inst = 32'hc404800;
      32679: inst = 32'h8220000;
      32680: inst = 32'h10408000;
      32681: inst = 32'hc404801;
      32682: inst = 32'h8220000;
      32683: inst = 32'h10408000;
      32684: inst = 32'hc404802;
      32685: inst = 32'h8220000;
      32686: inst = 32'h10408000;
      32687: inst = 32'hc404803;
      32688: inst = 32'h8220000;
      32689: inst = 32'h10408000;
      32690: inst = 32'hc404804;
      32691: inst = 32'h8220000;
      32692: inst = 32'h10408000;
      32693: inst = 32'hc404805;
      32694: inst = 32'h8220000;
      32695: inst = 32'h10408000;
      32696: inst = 32'hc404806;
      32697: inst = 32'h8220000;
      32698: inst = 32'h10408000;
      32699: inst = 32'hc404807;
      32700: inst = 32'h8220000;
      32701: inst = 32'h10408000;
      32702: inst = 32'hc404808;
      32703: inst = 32'h8220000;
      32704: inst = 32'h10408000;
      32705: inst = 32'hc404809;
      32706: inst = 32'h8220000;
      32707: inst = 32'h10408000;
      32708: inst = 32'hc40480a;
      32709: inst = 32'h8220000;
      32710: inst = 32'h10408000;
      32711: inst = 32'hc40480b;
      32712: inst = 32'h8220000;
      32713: inst = 32'h10408000;
      32714: inst = 32'hc40480f;
      32715: inst = 32'h8220000;
      32716: inst = 32'h10408000;
      32717: inst = 32'hc404810;
      32718: inst = 32'h8220000;
      32719: inst = 32'h10408000;
      32720: inst = 32'hc404811;
      32721: inst = 32'h8220000;
      32722: inst = 32'h10408000;
      32723: inst = 32'hc404812;
      32724: inst = 32'h8220000;
      32725: inst = 32'h10408000;
      32726: inst = 32'hc404813;
      32727: inst = 32'h8220000;
      32728: inst = 32'h10408000;
      32729: inst = 32'hc404814;
      32730: inst = 32'h8220000;
      32731: inst = 32'h10408000;
      32732: inst = 32'hc404815;
      32733: inst = 32'h8220000;
      32734: inst = 32'h10408000;
      32735: inst = 32'hc404816;
      32736: inst = 32'h8220000;
      32737: inst = 32'h10408000;
      32738: inst = 32'hc404817;
      32739: inst = 32'h8220000;
      32740: inst = 32'h10408000;
      32741: inst = 32'hc404818;
      32742: inst = 32'h8220000;
      32743: inst = 32'h10408000;
      32744: inst = 32'hc404819;
      32745: inst = 32'h8220000;
      32746: inst = 32'h10408000;
      32747: inst = 32'hc40481a;
      32748: inst = 32'h8220000;
      32749: inst = 32'h10408000;
      32750: inst = 32'hc40481b;
      32751: inst = 32'h8220000;
      32752: inst = 32'h10408000;
      32753: inst = 32'hc40481c;
      32754: inst = 32'h8220000;
      32755: inst = 32'h10408000;
      32756: inst = 32'hc404823;
      32757: inst = 32'h8220000;
      32758: inst = 32'h10408000;
      32759: inst = 32'hc404824;
      32760: inst = 32'h8220000;
      32761: inst = 32'h10408000;
      32762: inst = 32'hc404825;
      32763: inst = 32'h8220000;
      32764: inst = 32'h10408000;
      32765: inst = 32'hc404826;
      32766: inst = 32'h8220000;
      32767: inst = 32'h10408000;
      32768: inst = 32'hc404827;
      32769: inst = 32'h8220000;
      32770: inst = 32'h10408000;
      32771: inst = 32'hc404828;
      32772: inst = 32'h8220000;
      32773: inst = 32'h10408000;
      32774: inst = 32'hc404829;
      32775: inst = 32'h8220000;
      32776: inst = 32'h10408000;
      32777: inst = 32'hc40482a;
      32778: inst = 32'h8220000;
      32779: inst = 32'h10408000;
      32780: inst = 32'hc40482b;
      32781: inst = 32'h8220000;
      32782: inst = 32'h10408000;
      32783: inst = 32'hc40482c;
      32784: inst = 32'h8220000;
      32785: inst = 32'h10408000;
      32786: inst = 32'hc40482d;
      32787: inst = 32'h8220000;
      32788: inst = 32'h10408000;
      32789: inst = 32'hc404831;
      32790: inst = 32'h8220000;
      32791: inst = 32'h10408000;
      32792: inst = 32'hc404832;
      32793: inst = 32'h8220000;
      32794: inst = 32'h10408000;
      32795: inst = 32'hc404833;
      32796: inst = 32'h8220000;
      32797: inst = 32'h10408000;
      32798: inst = 32'hc404834;
      32799: inst = 32'h8220000;
      32800: inst = 32'h10408000;
      32801: inst = 32'hc404835;
      32802: inst = 32'h8220000;
      32803: inst = 32'h10408000;
      32804: inst = 32'hc404836;
      32805: inst = 32'h8220000;
      32806: inst = 32'h10408000;
      32807: inst = 32'hc404837;
      32808: inst = 32'h8220000;
      32809: inst = 32'h10408000;
      32810: inst = 32'hc404838;
      32811: inst = 32'h8220000;
      32812: inst = 32'h10408000;
      32813: inst = 32'hc404839;
      32814: inst = 32'h8220000;
      32815: inst = 32'h10408000;
      32816: inst = 32'hc40483a;
      32817: inst = 32'h8220000;
      32818: inst = 32'h10408000;
      32819: inst = 32'hc40483b;
      32820: inst = 32'h8220000;
      32821: inst = 32'h10408000;
      32822: inst = 32'hc40483c;
      32823: inst = 32'h8220000;
      32824: inst = 32'h10408000;
      32825: inst = 32'hc40483d;
      32826: inst = 32'h8220000;
      32827: inst = 32'h10408000;
      32828: inst = 32'hc40483e;
      32829: inst = 32'h8220000;
      32830: inst = 32'h10408000;
      32831: inst = 32'hc40483f;
      32832: inst = 32'h8220000;
      32833: inst = 32'h10408000;
      32834: inst = 32'hc404840;
      32835: inst = 32'h8220000;
      32836: inst = 32'h10408000;
      32837: inst = 32'hc404841;
      32838: inst = 32'h8220000;
      32839: inst = 32'h10408000;
      32840: inst = 32'hc404842;
      32841: inst = 32'h8220000;
      32842: inst = 32'h10408000;
      32843: inst = 32'hc404843;
      32844: inst = 32'h8220000;
      32845: inst = 32'h10408000;
      32846: inst = 32'hc404844;
      32847: inst = 32'h8220000;
      32848: inst = 32'h10408000;
      32849: inst = 32'hc404845;
      32850: inst = 32'h8220000;
      32851: inst = 32'h10408000;
      32852: inst = 32'hc404846;
      32853: inst = 32'h8220000;
      32854: inst = 32'h10408000;
      32855: inst = 32'hc404847;
      32856: inst = 32'h8220000;
      32857: inst = 32'h10408000;
      32858: inst = 32'hc404848;
      32859: inst = 32'h8220000;
      32860: inst = 32'h10408000;
      32861: inst = 32'hc404849;
      32862: inst = 32'h8220000;
      32863: inst = 32'h10408000;
      32864: inst = 32'hc40484a;
      32865: inst = 32'h8220000;
      32866: inst = 32'h10408000;
      32867: inst = 32'hc40484b;
      32868: inst = 32'h8220000;
      32869: inst = 32'h10408000;
      32870: inst = 32'hc40484c;
      32871: inst = 32'h8220000;
      32872: inst = 32'h10408000;
      32873: inst = 32'hc40484d;
      32874: inst = 32'h8220000;
      32875: inst = 32'h10408000;
      32876: inst = 32'hc40484e;
      32877: inst = 32'h8220000;
      32878: inst = 32'h10408000;
      32879: inst = 32'hc40484f;
      32880: inst = 32'h8220000;
      32881: inst = 32'h10408000;
      32882: inst = 32'hc404850;
      32883: inst = 32'h8220000;
      32884: inst = 32'h10408000;
      32885: inst = 32'hc404851;
      32886: inst = 32'h8220000;
      32887: inst = 32'h10408000;
      32888: inst = 32'hc404852;
      32889: inst = 32'h8220000;
      32890: inst = 32'h10408000;
      32891: inst = 32'hc404853;
      32892: inst = 32'h8220000;
      32893: inst = 32'h10408000;
      32894: inst = 32'hc40485a;
      32895: inst = 32'h8220000;
      32896: inst = 32'h10408000;
      32897: inst = 32'hc40485b;
      32898: inst = 32'h8220000;
      32899: inst = 32'h10408000;
      32900: inst = 32'hc40485c;
      32901: inst = 32'h8220000;
      32902: inst = 32'h10408000;
      32903: inst = 32'hc40485d;
      32904: inst = 32'h8220000;
      32905: inst = 32'h10408000;
      32906: inst = 32'hc40485e;
      32907: inst = 32'h8220000;
      32908: inst = 32'h10408000;
      32909: inst = 32'hc40485f;
      32910: inst = 32'h8220000;
      32911: inst = 32'h10408000;
      32912: inst = 32'hc404860;
      32913: inst = 32'h8220000;
      32914: inst = 32'h10408000;
      32915: inst = 32'hc404861;
      32916: inst = 32'h8220000;
      32917: inst = 32'h10408000;
      32918: inst = 32'hc404862;
      32919: inst = 32'h8220000;
      32920: inst = 32'h10408000;
      32921: inst = 32'hc404863;
      32922: inst = 32'h8220000;
      32923: inst = 32'h10408000;
      32924: inst = 32'hc404864;
      32925: inst = 32'h8220000;
      32926: inst = 32'h10408000;
      32927: inst = 32'hc404865;
      32928: inst = 32'h8220000;
      32929: inst = 32'h10408000;
      32930: inst = 32'hc404866;
      32931: inst = 32'h8220000;
      32932: inst = 32'h10408000;
      32933: inst = 32'hc404867;
      32934: inst = 32'h8220000;
      32935: inst = 32'h10408000;
      32936: inst = 32'hc404868;
      32937: inst = 32'h8220000;
      32938: inst = 32'h10408000;
      32939: inst = 32'hc404869;
      32940: inst = 32'h8220000;
      32941: inst = 32'h10408000;
      32942: inst = 32'hc40486a;
      32943: inst = 32'h8220000;
      32944: inst = 32'h10408000;
      32945: inst = 32'hc40486b;
      32946: inst = 32'h8220000;
      32947: inst = 32'h10408000;
      32948: inst = 32'hc40486f;
      32949: inst = 32'h8220000;
      32950: inst = 32'h10408000;
      32951: inst = 32'hc404870;
      32952: inst = 32'h8220000;
      32953: inst = 32'h10408000;
      32954: inst = 32'hc404871;
      32955: inst = 32'h8220000;
      32956: inst = 32'h10408000;
      32957: inst = 32'hc404872;
      32958: inst = 32'h8220000;
      32959: inst = 32'h10408000;
      32960: inst = 32'hc404873;
      32961: inst = 32'h8220000;
      32962: inst = 32'h10408000;
      32963: inst = 32'hc404874;
      32964: inst = 32'h8220000;
      32965: inst = 32'h10408000;
      32966: inst = 32'hc404875;
      32967: inst = 32'h8220000;
      32968: inst = 32'h10408000;
      32969: inst = 32'hc404876;
      32970: inst = 32'h8220000;
      32971: inst = 32'h10408000;
      32972: inst = 32'hc404877;
      32973: inst = 32'h8220000;
      32974: inst = 32'h10408000;
      32975: inst = 32'hc404878;
      32976: inst = 32'h8220000;
      32977: inst = 32'h10408000;
      32978: inst = 32'hc404879;
      32979: inst = 32'h8220000;
      32980: inst = 32'h10408000;
      32981: inst = 32'hc40487a;
      32982: inst = 32'h8220000;
      32983: inst = 32'h10408000;
      32984: inst = 32'hc40487b;
      32985: inst = 32'h8220000;
      32986: inst = 32'h10408000;
      32987: inst = 32'hc40487c;
      32988: inst = 32'h8220000;
      32989: inst = 32'h10408000;
      32990: inst = 32'hc404883;
      32991: inst = 32'h8220000;
      32992: inst = 32'h10408000;
      32993: inst = 32'hc404884;
      32994: inst = 32'h8220000;
      32995: inst = 32'h10408000;
      32996: inst = 32'hc404885;
      32997: inst = 32'h8220000;
      32998: inst = 32'h10408000;
      32999: inst = 32'hc404886;
      33000: inst = 32'h8220000;
      33001: inst = 32'h10408000;
      33002: inst = 32'hc404887;
      33003: inst = 32'h8220000;
      33004: inst = 32'h10408000;
      33005: inst = 32'hc404888;
      33006: inst = 32'h8220000;
      33007: inst = 32'h10408000;
      33008: inst = 32'hc404889;
      33009: inst = 32'h8220000;
      33010: inst = 32'h10408000;
      33011: inst = 32'hc40488a;
      33012: inst = 32'h8220000;
      33013: inst = 32'h10408000;
      33014: inst = 32'hc40488b;
      33015: inst = 32'h8220000;
      33016: inst = 32'h10408000;
      33017: inst = 32'hc40488c;
      33018: inst = 32'h8220000;
      33019: inst = 32'h10408000;
      33020: inst = 32'hc40488d;
      33021: inst = 32'h8220000;
      33022: inst = 32'h10408000;
      33023: inst = 32'hc404891;
      33024: inst = 32'h8220000;
      33025: inst = 32'h10408000;
      33026: inst = 32'hc404892;
      33027: inst = 32'h8220000;
      33028: inst = 32'h10408000;
      33029: inst = 32'hc404893;
      33030: inst = 32'h8220000;
      33031: inst = 32'h10408000;
      33032: inst = 32'hc404894;
      33033: inst = 32'h8220000;
      33034: inst = 32'h10408000;
      33035: inst = 32'hc404895;
      33036: inst = 32'h8220000;
      33037: inst = 32'h10408000;
      33038: inst = 32'hc404896;
      33039: inst = 32'h8220000;
      33040: inst = 32'h10408000;
      33041: inst = 32'hc404897;
      33042: inst = 32'h8220000;
      33043: inst = 32'h10408000;
      33044: inst = 32'hc404898;
      33045: inst = 32'h8220000;
      33046: inst = 32'h10408000;
      33047: inst = 32'hc404899;
      33048: inst = 32'h8220000;
      33049: inst = 32'h10408000;
      33050: inst = 32'hc40489a;
      33051: inst = 32'h8220000;
      33052: inst = 32'h10408000;
      33053: inst = 32'hc40489b;
      33054: inst = 32'h8220000;
      33055: inst = 32'h10408000;
      33056: inst = 32'hc40489c;
      33057: inst = 32'h8220000;
      33058: inst = 32'h10408000;
      33059: inst = 32'hc40489d;
      33060: inst = 32'h8220000;
      33061: inst = 32'h10408000;
      33062: inst = 32'hc40489e;
      33063: inst = 32'h8220000;
      33064: inst = 32'h10408000;
      33065: inst = 32'hc40489f;
      33066: inst = 32'h8220000;
      33067: inst = 32'h10408000;
      33068: inst = 32'hc4048a0;
      33069: inst = 32'h8220000;
      33070: inst = 32'h10408000;
      33071: inst = 32'hc4048a1;
      33072: inst = 32'h8220000;
      33073: inst = 32'h10408000;
      33074: inst = 32'hc4048a2;
      33075: inst = 32'h8220000;
      33076: inst = 32'h10408000;
      33077: inst = 32'hc4048a3;
      33078: inst = 32'h8220000;
      33079: inst = 32'h10408000;
      33080: inst = 32'hc4048a4;
      33081: inst = 32'h8220000;
      33082: inst = 32'h10408000;
      33083: inst = 32'hc4048a5;
      33084: inst = 32'h8220000;
      33085: inst = 32'h10408000;
      33086: inst = 32'hc4048a6;
      33087: inst = 32'h8220000;
      33088: inst = 32'h10408000;
      33089: inst = 32'hc4048a7;
      33090: inst = 32'h8220000;
      33091: inst = 32'h10408000;
      33092: inst = 32'hc4048a8;
      33093: inst = 32'h8220000;
      33094: inst = 32'h10408000;
      33095: inst = 32'hc4048a9;
      33096: inst = 32'h8220000;
      33097: inst = 32'h10408000;
      33098: inst = 32'hc4048aa;
      33099: inst = 32'h8220000;
      33100: inst = 32'h10408000;
      33101: inst = 32'hc4048ab;
      33102: inst = 32'h8220000;
      33103: inst = 32'h10408000;
      33104: inst = 32'hc4048ac;
      33105: inst = 32'h8220000;
      33106: inst = 32'h10408000;
      33107: inst = 32'hc4048ad;
      33108: inst = 32'h8220000;
      33109: inst = 32'h10408000;
      33110: inst = 32'hc4048ae;
      33111: inst = 32'h8220000;
      33112: inst = 32'h10408000;
      33113: inst = 32'hc4048af;
      33114: inst = 32'h8220000;
      33115: inst = 32'h10408000;
      33116: inst = 32'hc4048b0;
      33117: inst = 32'h8220000;
      33118: inst = 32'h10408000;
      33119: inst = 32'hc4048b1;
      33120: inst = 32'h8220000;
      33121: inst = 32'h10408000;
      33122: inst = 32'hc4048b2;
      33123: inst = 32'h8220000;
      33124: inst = 32'h10408000;
      33125: inst = 32'hc4048b3;
      33126: inst = 32'h8220000;
      33127: inst = 32'h10408000;
      33128: inst = 32'hc4048ba;
      33129: inst = 32'h8220000;
      33130: inst = 32'h10408000;
      33131: inst = 32'hc4048bb;
      33132: inst = 32'h8220000;
      33133: inst = 32'h10408000;
      33134: inst = 32'hc4048bc;
      33135: inst = 32'h8220000;
      33136: inst = 32'h10408000;
      33137: inst = 32'hc4048bd;
      33138: inst = 32'h8220000;
      33139: inst = 32'h10408000;
      33140: inst = 32'hc4048be;
      33141: inst = 32'h8220000;
      33142: inst = 32'h10408000;
      33143: inst = 32'hc4048bf;
      33144: inst = 32'h8220000;
      33145: inst = 32'h10408000;
      33146: inst = 32'hc4048c0;
      33147: inst = 32'h8220000;
      33148: inst = 32'h10408000;
      33149: inst = 32'hc4048c1;
      33150: inst = 32'h8220000;
      33151: inst = 32'h10408000;
      33152: inst = 32'hc4048c2;
      33153: inst = 32'h8220000;
      33154: inst = 32'h10408000;
      33155: inst = 32'hc4048c3;
      33156: inst = 32'h8220000;
      33157: inst = 32'h10408000;
      33158: inst = 32'hc4048c4;
      33159: inst = 32'h8220000;
      33160: inst = 32'h10408000;
      33161: inst = 32'hc4048c5;
      33162: inst = 32'h8220000;
      33163: inst = 32'h10408000;
      33164: inst = 32'hc4048c6;
      33165: inst = 32'h8220000;
      33166: inst = 32'h10408000;
      33167: inst = 32'hc4048c7;
      33168: inst = 32'h8220000;
      33169: inst = 32'h10408000;
      33170: inst = 32'hc4048c8;
      33171: inst = 32'h8220000;
      33172: inst = 32'h10408000;
      33173: inst = 32'hc4048c9;
      33174: inst = 32'h8220000;
      33175: inst = 32'h10408000;
      33176: inst = 32'hc4048ca;
      33177: inst = 32'h8220000;
      33178: inst = 32'h10408000;
      33179: inst = 32'hc4048cb;
      33180: inst = 32'h8220000;
      33181: inst = 32'h10408000;
      33182: inst = 32'hc4048cf;
      33183: inst = 32'h8220000;
      33184: inst = 32'h10408000;
      33185: inst = 32'hc4048d0;
      33186: inst = 32'h8220000;
      33187: inst = 32'h10408000;
      33188: inst = 32'hc4048d1;
      33189: inst = 32'h8220000;
      33190: inst = 32'h10408000;
      33191: inst = 32'hc4048d2;
      33192: inst = 32'h8220000;
      33193: inst = 32'h10408000;
      33194: inst = 32'hc4048d3;
      33195: inst = 32'h8220000;
      33196: inst = 32'h10408000;
      33197: inst = 32'hc4048d4;
      33198: inst = 32'h8220000;
      33199: inst = 32'h10408000;
      33200: inst = 32'hc4048d5;
      33201: inst = 32'h8220000;
      33202: inst = 32'h10408000;
      33203: inst = 32'hc4048d6;
      33204: inst = 32'h8220000;
      33205: inst = 32'h10408000;
      33206: inst = 32'hc4048d7;
      33207: inst = 32'h8220000;
      33208: inst = 32'h10408000;
      33209: inst = 32'hc4048d8;
      33210: inst = 32'h8220000;
      33211: inst = 32'h10408000;
      33212: inst = 32'hc4048d9;
      33213: inst = 32'h8220000;
      33214: inst = 32'h10408000;
      33215: inst = 32'hc4048da;
      33216: inst = 32'h8220000;
      33217: inst = 32'h10408000;
      33218: inst = 32'hc4048db;
      33219: inst = 32'h8220000;
      33220: inst = 32'h10408000;
      33221: inst = 32'hc4048dc;
      33222: inst = 32'h8220000;
      33223: inst = 32'h10408000;
      33224: inst = 32'hc4048e3;
      33225: inst = 32'h8220000;
      33226: inst = 32'h10408000;
      33227: inst = 32'hc4048e4;
      33228: inst = 32'h8220000;
      33229: inst = 32'h10408000;
      33230: inst = 32'hc4048e5;
      33231: inst = 32'h8220000;
      33232: inst = 32'h10408000;
      33233: inst = 32'hc4048e6;
      33234: inst = 32'h8220000;
      33235: inst = 32'h10408000;
      33236: inst = 32'hc4048e7;
      33237: inst = 32'h8220000;
      33238: inst = 32'h10408000;
      33239: inst = 32'hc4048e8;
      33240: inst = 32'h8220000;
      33241: inst = 32'h10408000;
      33242: inst = 32'hc4048e9;
      33243: inst = 32'h8220000;
      33244: inst = 32'h10408000;
      33245: inst = 32'hc4048ea;
      33246: inst = 32'h8220000;
      33247: inst = 32'h10408000;
      33248: inst = 32'hc4048eb;
      33249: inst = 32'h8220000;
      33250: inst = 32'h10408000;
      33251: inst = 32'hc4048ec;
      33252: inst = 32'h8220000;
      33253: inst = 32'h10408000;
      33254: inst = 32'hc4048ed;
      33255: inst = 32'h8220000;
      33256: inst = 32'h10408000;
      33257: inst = 32'hc4048f1;
      33258: inst = 32'h8220000;
      33259: inst = 32'h10408000;
      33260: inst = 32'hc4048f2;
      33261: inst = 32'h8220000;
      33262: inst = 32'h10408000;
      33263: inst = 32'hc4048f3;
      33264: inst = 32'h8220000;
      33265: inst = 32'h10408000;
      33266: inst = 32'hc4048f4;
      33267: inst = 32'h8220000;
      33268: inst = 32'h10408000;
      33269: inst = 32'hc4048f5;
      33270: inst = 32'h8220000;
      33271: inst = 32'h10408000;
      33272: inst = 32'hc4048f6;
      33273: inst = 32'h8220000;
      33274: inst = 32'h10408000;
      33275: inst = 32'hc4048f7;
      33276: inst = 32'h8220000;
      33277: inst = 32'h10408000;
      33278: inst = 32'hc4048f8;
      33279: inst = 32'h8220000;
      33280: inst = 32'h10408000;
      33281: inst = 32'hc4048f9;
      33282: inst = 32'h8220000;
      33283: inst = 32'h10408000;
      33284: inst = 32'hc4048fa;
      33285: inst = 32'h8220000;
      33286: inst = 32'h10408000;
      33287: inst = 32'hc4048fb;
      33288: inst = 32'h8220000;
      33289: inst = 32'h10408000;
      33290: inst = 32'hc4048fc;
      33291: inst = 32'h8220000;
      33292: inst = 32'h10408000;
      33293: inst = 32'hc4048fd;
      33294: inst = 32'h8220000;
      33295: inst = 32'h10408000;
      33296: inst = 32'hc4048fe;
      33297: inst = 32'h8220000;
      33298: inst = 32'h10408000;
      33299: inst = 32'hc4048ff;
      33300: inst = 32'h8220000;
      33301: inst = 32'h10408000;
      33302: inst = 32'hc404900;
      33303: inst = 32'h8220000;
      33304: inst = 32'h10408000;
      33305: inst = 32'hc404901;
      33306: inst = 32'h8220000;
      33307: inst = 32'h10408000;
      33308: inst = 32'hc404902;
      33309: inst = 32'h8220000;
      33310: inst = 32'h10408000;
      33311: inst = 32'hc404903;
      33312: inst = 32'h8220000;
      33313: inst = 32'h10408000;
      33314: inst = 32'hc404904;
      33315: inst = 32'h8220000;
      33316: inst = 32'h10408000;
      33317: inst = 32'hc404905;
      33318: inst = 32'h8220000;
      33319: inst = 32'h10408000;
      33320: inst = 32'hc404906;
      33321: inst = 32'h8220000;
      33322: inst = 32'h10408000;
      33323: inst = 32'hc404907;
      33324: inst = 32'h8220000;
      33325: inst = 32'h10408000;
      33326: inst = 32'hc404908;
      33327: inst = 32'h8220000;
      33328: inst = 32'h10408000;
      33329: inst = 32'hc404909;
      33330: inst = 32'h8220000;
      33331: inst = 32'h10408000;
      33332: inst = 32'hc40490a;
      33333: inst = 32'h8220000;
      33334: inst = 32'h10408000;
      33335: inst = 32'hc40490b;
      33336: inst = 32'h8220000;
      33337: inst = 32'h10408000;
      33338: inst = 32'hc40490c;
      33339: inst = 32'h8220000;
      33340: inst = 32'h10408000;
      33341: inst = 32'hc40490d;
      33342: inst = 32'h8220000;
      33343: inst = 32'h10408000;
      33344: inst = 32'hc40490e;
      33345: inst = 32'h8220000;
      33346: inst = 32'h10408000;
      33347: inst = 32'hc40490f;
      33348: inst = 32'h8220000;
      33349: inst = 32'h10408000;
      33350: inst = 32'hc404910;
      33351: inst = 32'h8220000;
      33352: inst = 32'h10408000;
      33353: inst = 32'hc404911;
      33354: inst = 32'h8220000;
      33355: inst = 32'h10408000;
      33356: inst = 32'hc404912;
      33357: inst = 32'h8220000;
      33358: inst = 32'h10408000;
      33359: inst = 32'hc404913;
      33360: inst = 32'h8220000;
      33361: inst = 32'h10408000;
      33362: inst = 32'hc404916;
      33363: inst = 32'h8220000;
      33364: inst = 32'h10408000;
      33365: inst = 32'hc40491a;
      33366: inst = 32'h8220000;
      33367: inst = 32'h10408000;
      33368: inst = 32'hc40491b;
      33369: inst = 32'h8220000;
      33370: inst = 32'h10408000;
      33371: inst = 32'hc40491c;
      33372: inst = 32'h8220000;
      33373: inst = 32'h10408000;
      33374: inst = 32'hc40491d;
      33375: inst = 32'h8220000;
      33376: inst = 32'h10408000;
      33377: inst = 32'hc40491e;
      33378: inst = 32'h8220000;
      33379: inst = 32'h10408000;
      33380: inst = 32'hc40491f;
      33381: inst = 32'h8220000;
      33382: inst = 32'h10408000;
      33383: inst = 32'hc404920;
      33384: inst = 32'h8220000;
      33385: inst = 32'h10408000;
      33386: inst = 32'hc404921;
      33387: inst = 32'h8220000;
      33388: inst = 32'h10408000;
      33389: inst = 32'hc404922;
      33390: inst = 32'h8220000;
      33391: inst = 32'h10408000;
      33392: inst = 32'hc404923;
      33393: inst = 32'h8220000;
      33394: inst = 32'h10408000;
      33395: inst = 32'hc404924;
      33396: inst = 32'h8220000;
      33397: inst = 32'h10408000;
      33398: inst = 32'hc404925;
      33399: inst = 32'h8220000;
      33400: inst = 32'h10408000;
      33401: inst = 32'hc404926;
      33402: inst = 32'h8220000;
      33403: inst = 32'h10408000;
      33404: inst = 32'hc404927;
      33405: inst = 32'h8220000;
      33406: inst = 32'h10408000;
      33407: inst = 32'hc404928;
      33408: inst = 32'h8220000;
      33409: inst = 32'h10408000;
      33410: inst = 32'hc404929;
      33411: inst = 32'h8220000;
      33412: inst = 32'h10408000;
      33413: inst = 32'hc40492a;
      33414: inst = 32'h8220000;
      33415: inst = 32'h10408000;
      33416: inst = 32'hc40492b;
      33417: inst = 32'h8220000;
      33418: inst = 32'h10408000;
      33419: inst = 32'hc40492f;
      33420: inst = 32'h8220000;
      33421: inst = 32'h10408000;
      33422: inst = 32'hc404930;
      33423: inst = 32'h8220000;
      33424: inst = 32'h10408000;
      33425: inst = 32'hc404931;
      33426: inst = 32'h8220000;
      33427: inst = 32'h10408000;
      33428: inst = 32'hc404932;
      33429: inst = 32'h8220000;
      33430: inst = 32'h10408000;
      33431: inst = 32'hc404933;
      33432: inst = 32'h8220000;
      33433: inst = 32'h10408000;
      33434: inst = 32'hc404934;
      33435: inst = 32'h8220000;
      33436: inst = 32'h10408000;
      33437: inst = 32'hc404935;
      33438: inst = 32'h8220000;
      33439: inst = 32'h10408000;
      33440: inst = 32'hc404936;
      33441: inst = 32'h8220000;
      33442: inst = 32'h10408000;
      33443: inst = 32'hc404937;
      33444: inst = 32'h8220000;
      33445: inst = 32'h10408000;
      33446: inst = 32'hc404938;
      33447: inst = 32'h8220000;
      33448: inst = 32'h10408000;
      33449: inst = 32'hc404939;
      33450: inst = 32'h8220000;
      33451: inst = 32'h10408000;
      33452: inst = 32'hc40493a;
      33453: inst = 32'h8220000;
      33454: inst = 32'h10408000;
      33455: inst = 32'hc40493b;
      33456: inst = 32'h8220000;
      33457: inst = 32'h10408000;
      33458: inst = 32'hc40493c;
      33459: inst = 32'h8220000;
      33460: inst = 32'h10408000;
      33461: inst = 32'hc404943;
      33462: inst = 32'h8220000;
      33463: inst = 32'h10408000;
      33464: inst = 32'hc404944;
      33465: inst = 32'h8220000;
      33466: inst = 32'h10408000;
      33467: inst = 32'hc404945;
      33468: inst = 32'h8220000;
      33469: inst = 32'h10408000;
      33470: inst = 32'hc404946;
      33471: inst = 32'h8220000;
      33472: inst = 32'h10408000;
      33473: inst = 32'hc404947;
      33474: inst = 32'h8220000;
      33475: inst = 32'h10408000;
      33476: inst = 32'hc404948;
      33477: inst = 32'h8220000;
      33478: inst = 32'h10408000;
      33479: inst = 32'hc404949;
      33480: inst = 32'h8220000;
      33481: inst = 32'h10408000;
      33482: inst = 32'hc40494a;
      33483: inst = 32'h8220000;
      33484: inst = 32'h10408000;
      33485: inst = 32'hc40494b;
      33486: inst = 32'h8220000;
      33487: inst = 32'h10408000;
      33488: inst = 32'hc40494c;
      33489: inst = 32'h8220000;
      33490: inst = 32'h10408000;
      33491: inst = 32'hc40494d;
      33492: inst = 32'h8220000;
      33493: inst = 32'h10408000;
      33494: inst = 32'hc404951;
      33495: inst = 32'h8220000;
      33496: inst = 32'h10408000;
      33497: inst = 32'hc404952;
      33498: inst = 32'h8220000;
      33499: inst = 32'h10408000;
      33500: inst = 32'hc404953;
      33501: inst = 32'h8220000;
      33502: inst = 32'h10408000;
      33503: inst = 32'hc404954;
      33504: inst = 32'h8220000;
      33505: inst = 32'h10408000;
      33506: inst = 32'hc404955;
      33507: inst = 32'h8220000;
      33508: inst = 32'h10408000;
      33509: inst = 32'hc404956;
      33510: inst = 32'h8220000;
      33511: inst = 32'h10408000;
      33512: inst = 32'hc404957;
      33513: inst = 32'h8220000;
      33514: inst = 32'h10408000;
      33515: inst = 32'hc404958;
      33516: inst = 32'h8220000;
      33517: inst = 32'h10408000;
      33518: inst = 32'hc404959;
      33519: inst = 32'h8220000;
      33520: inst = 32'h10408000;
      33521: inst = 32'hc40495a;
      33522: inst = 32'h8220000;
      33523: inst = 32'h10408000;
      33524: inst = 32'hc40495b;
      33525: inst = 32'h8220000;
      33526: inst = 32'h10408000;
      33527: inst = 32'hc40495c;
      33528: inst = 32'h8220000;
      33529: inst = 32'h10408000;
      33530: inst = 32'hc40495d;
      33531: inst = 32'h8220000;
      33532: inst = 32'h10408000;
      33533: inst = 32'hc40495e;
      33534: inst = 32'h8220000;
      33535: inst = 32'h10408000;
      33536: inst = 32'hc40495f;
      33537: inst = 32'h8220000;
      33538: inst = 32'h10408000;
      33539: inst = 32'hc404960;
      33540: inst = 32'h8220000;
      33541: inst = 32'h10408000;
      33542: inst = 32'hc404961;
      33543: inst = 32'h8220000;
      33544: inst = 32'h10408000;
      33545: inst = 32'hc404962;
      33546: inst = 32'h8220000;
      33547: inst = 32'h10408000;
      33548: inst = 32'hc404963;
      33549: inst = 32'h8220000;
      33550: inst = 32'h10408000;
      33551: inst = 32'hc404964;
      33552: inst = 32'h8220000;
      33553: inst = 32'h10408000;
      33554: inst = 32'hc404965;
      33555: inst = 32'h8220000;
      33556: inst = 32'h10408000;
      33557: inst = 32'hc404966;
      33558: inst = 32'h8220000;
      33559: inst = 32'h10408000;
      33560: inst = 32'hc404967;
      33561: inst = 32'h8220000;
      33562: inst = 32'h10408000;
      33563: inst = 32'hc404968;
      33564: inst = 32'h8220000;
      33565: inst = 32'h10408000;
      33566: inst = 32'hc404969;
      33567: inst = 32'h8220000;
      33568: inst = 32'h10408000;
      33569: inst = 32'hc40496a;
      33570: inst = 32'h8220000;
      33571: inst = 32'h10408000;
      33572: inst = 32'hc40496b;
      33573: inst = 32'h8220000;
      33574: inst = 32'h10408000;
      33575: inst = 32'hc40496c;
      33576: inst = 32'h8220000;
      33577: inst = 32'h10408000;
      33578: inst = 32'hc40496d;
      33579: inst = 32'h8220000;
      33580: inst = 32'h10408000;
      33581: inst = 32'hc40496e;
      33582: inst = 32'h8220000;
      33583: inst = 32'h10408000;
      33584: inst = 32'hc40496f;
      33585: inst = 32'h8220000;
      33586: inst = 32'h10408000;
      33587: inst = 32'hc404970;
      33588: inst = 32'h8220000;
      33589: inst = 32'h10408000;
      33590: inst = 32'hc404971;
      33591: inst = 32'h8220000;
      33592: inst = 32'h10408000;
      33593: inst = 32'hc404972;
      33594: inst = 32'h8220000;
      33595: inst = 32'h10408000;
      33596: inst = 32'hc404973;
      33597: inst = 32'h8220000;
      33598: inst = 32'h10408000;
      33599: inst = 32'hc404974;
      33600: inst = 32'h8220000;
      33601: inst = 32'h10408000;
      33602: inst = 32'hc404975;
      33603: inst = 32'h8220000;
      33604: inst = 32'h10408000;
      33605: inst = 32'hc404976;
      33606: inst = 32'h8220000;
      33607: inst = 32'h10408000;
      33608: inst = 32'hc404977;
      33609: inst = 32'h8220000;
      33610: inst = 32'h10408000;
      33611: inst = 32'hc404978;
      33612: inst = 32'h8220000;
      33613: inst = 32'h10408000;
      33614: inst = 32'hc404979;
      33615: inst = 32'h8220000;
      33616: inst = 32'h10408000;
      33617: inst = 32'hc40497a;
      33618: inst = 32'h8220000;
      33619: inst = 32'h10408000;
      33620: inst = 32'hc40497b;
      33621: inst = 32'h8220000;
      33622: inst = 32'h10408000;
      33623: inst = 32'hc40497c;
      33624: inst = 32'h8220000;
      33625: inst = 32'h10408000;
      33626: inst = 32'hc40497d;
      33627: inst = 32'h8220000;
      33628: inst = 32'h10408000;
      33629: inst = 32'hc40497e;
      33630: inst = 32'h8220000;
      33631: inst = 32'h10408000;
      33632: inst = 32'hc40497f;
      33633: inst = 32'h8220000;
      33634: inst = 32'h10408000;
      33635: inst = 32'hc404980;
      33636: inst = 32'h8220000;
      33637: inst = 32'h10408000;
      33638: inst = 32'hc404981;
      33639: inst = 32'h8220000;
      33640: inst = 32'h10408000;
      33641: inst = 32'hc404982;
      33642: inst = 32'h8220000;
      33643: inst = 32'h10408000;
      33644: inst = 32'hc404983;
      33645: inst = 32'h8220000;
      33646: inst = 32'h10408000;
      33647: inst = 32'hc404984;
      33648: inst = 32'h8220000;
      33649: inst = 32'h10408000;
      33650: inst = 32'hc404985;
      33651: inst = 32'h8220000;
      33652: inst = 32'h10408000;
      33653: inst = 32'hc40498f;
      33654: inst = 32'h8220000;
      33655: inst = 32'h10408000;
      33656: inst = 32'hc404990;
      33657: inst = 32'h8220000;
      33658: inst = 32'h10408000;
      33659: inst = 32'hc404991;
      33660: inst = 32'h8220000;
      33661: inst = 32'h10408000;
      33662: inst = 32'hc404992;
      33663: inst = 32'h8220000;
      33664: inst = 32'h10408000;
      33665: inst = 32'hc404993;
      33666: inst = 32'h8220000;
      33667: inst = 32'h10408000;
      33668: inst = 32'hc404994;
      33669: inst = 32'h8220000;
      33670: inst = 32'h10408000;
      33671: inst = 32'hc404995;
      33672: inst = 32'h8220000;
      33673: inst = 32'h10408000;
      33674: inst = 32'hc404996;
      33675: inst = 32'h8220000;
      33676: inst = 32'h10408000;
      33677: inst = 32'hc404997;
      33678: inst = 32'h8220000;
      33679: inst = 32'h10408000;
      33680: inst = 32'hc404998;
      33681: inst = 32'h8220000;
      33682: inst = 32'h10408000;
      33683: inst = 32'hc404999;
      33684: inst = 32'h8220000;
      33685: inst = 32'h10408000;
      33686: inst = 32'hc40499a;
      33687: inst = 32'h8220000;
      33688: inst = 32'h10408000;
      33689: inst = 32'hc40499b;
      33690: inst = 32'h8220000;
      33691: inst = 32'h10408000;
      33692: inst = 32'hc40499c;
      33693: inst = 32'h8220000;
      33694: inst = 32'h10408000;
      33695: inst = 32'hc4049a3;
      33696: inst = 32'h8220000;
      33697: inst = 32'h10408000;
      33698: inst = 32'hc4049a4;
      33699: inst = 32'h8220000;
      33700: inst = 32'h10408000;
      33701: inst = 32'hc4049a5;
      33702: inst = 32'h8220000;
      33703: inst = 32'h10408000;
      33704: inst = 32'hc4049a6;
      33705: inst = 32'h8220000;
      33706: inst = 32'h10408000;
      33707: inst = 32'hc4049a7;
      33708: inst = 32'h8220000;
      33709: inst = 32'h10408000;
      33710: inst = 32'hc4049a8;
      33711: inst = 32'h8220000;
      33712: inst = 32'h10408000;
      33713: inst = 32'hc4049a9;
      33714: inst = 32'h8220000;
      33715: inst = 32'h10408000;
      33716: inst = 32'hc4049aa;
      33717: inst = 32'h8220000;
      33718: inst = 32'h10408000;
      33719: inst = 32'hc4049ab;
      33720: inst = 32'h8220000;
      33721: inst = 32'h10408000;
      33722: inst = 32'hc4049ac;
      33723: inst = 32'h8220000;
      33724: inst = 32'h10408000;
      33725: inst = 32'hc4049ad;
      33726: inst = 32'h8220000;
      33727: inst = 32'h10408000;
      33728: inst = 32'hc4049b1;
      33729: inst = 32'h8220000;
      33730: inst = 32'h10408000;
      33731: inst = 32'hc4049b2;
      33732: inst = 32'h8220000;
      33733: inst = 32'h10408000;
      33734: inst = 32'hc4049b3;
      33735: inst = 32'h8220000;
      33736: inst = 32'h10408000;
      33737: inst = 32'hc4049b4;
      33738: inst = 32'h8220000;
      33739: inst = 32'h10408000;
      33740: inst = 32'hc4049b5;
      33741: inst = 32'h8220000;
      33742: inst = 32'h10408000;
      33743: inst = 32'hc4049b6;
      33744: inst = 32'h8220000;
      33745: inst = 32'h10408000;
      33746: inst = 32'hc4049b7;
      33747: inst = 32'h8220000;
      33748: inst = 32'h10408000;
      33749: inst = 32'hc4049b8;
      33750: inst = 32'h8220000;
      33751: inst = 32'h10408000;
      33752: inst = 32'hc4049b9;
      33753: inst = 32'h8220000;
      33754: inst = 32'h10408000;
      33755: inst = 32'hc4049ba;
      33756: inst = 32'h8220000;
      33757: inst = 32'h10408000;
      33758: inst = 32'hc4049bb;
      33759: inst = 32'h8220000;
      33760: inst = 32'h10408000;
      33761: inst = 32'hc4049bc;
      33762: inst = 32'h8220000;
      33763: inst = 32'h10408000;
      33764: inst = 32'hc4049bd;
      33765: inst = 32'h8220000;
      33766: inst = 32'h10408000;
      33767: inst = 32'hc4049be;
      33768: inst = 32'h8220000;
      33769: inst = 32'h10408000;
      33770: inst = 32'hc4049bf;
      33771: inst = 32'h8220000;
      33772: inst = 32'h10408000;
      33773: inst = 32'hc4049c0;
      33774: inst = 32'h8220000;
      33775: inst = 32'h10408000;
      33776: inst = 32'hc4049c1;
      33777: inst = 32'h8220000;
      33778: inst = 32'h10408000;
      33779: inst = 32'hc4049c2;
      33780: inst = 32'h8220000;
      33781: inst = 32'h10408000;
      33782: inst = 32'hc4049c3;
      33783: inst = 32'h8220000;
      33784: inst = 32'h10408000;
      33785: inst = 32'hc4049c4;
      33786: inst = 32'h8220000;
      33787: inst = 32'h10408000;
      33788: inst = 32'hc4049c5;
      33789: inst = 32'h8220000;
      33790: inst = 32'h10408000;
      33791: inst = 32'hc4049c6;
      33792: inst = 32'h8220000;
      33793: inst = 32'h10408000;
      33794: inst = 32'hc4049c7;
      33795: inst = 32'h8220000;
      33796: inst = 32'h10408000;
      33797: inst = 32'hc4049c8;
      33798: inst = 32'h8220000;
      33799: inst = 32'h10408000;
      33800: inst = 32'hc4049c9;
      33801: inst = 32'h8220000;
      33802: inst = 32'h10408000;
      33803: inst = 32'hc4049ca;
      33804: inst = 32'h8220000;
      33805: inst = 32'h10408000;
      33806: inst = 32'hc4049cb;
      33807: inst = 32'h8220000;
      33808: inst = 32'h10408000;
      33809: inst = 32'hc4049cc;
      33810: inst = 32'h8220000;
      33811: inst = 32'h10408000;
      33812: inst = 32'hc4049cd;
      33813: inst = 32'h8220000;
      33814: inst = 32'h10408000;
      33815: inst = 32'hc4049ce;
      33816: inst = 32'h8220000;
      33817: inst = 32'h10408000;
      33818: inst = 32'hc4049cf;
      33819: inst = 32'h8220000;
      33820: inst = 32'h10408000;
      33821: inst = 32'hc4049d0;
      33822: inst = 32'h8220000;
      33823: inst = 32'h10408000;
      33824: inst = 32'hc4049d1;
      33825: inst = 32'h8220000;
      33826: inst = 32'h10408000;
      33827: inst = 32'hc4049d2;
      33828: inst = 32'h8220000;
      33829: inst = 32'h10408000;
      33830: inst = 32'hc4049d3;
      33831: inst = 32'h8220000;
      33832: inst = 32'h10408000;
      33833: inst = 32'hc4049d4;
      33834: inst = 32'h8220000;
      33835: inst = 32'h10408000;
      33836: inst = 32'hc4049d5;
      33837: inst = 32'h8220000;
      33838: inst = 32'h10408000;
      33839: inst = 32'hc4049d6;
      33840: inst = 32'h8220000;
      33841: inst = 32'h10408000;
      33842: inst = 32'hc4049d7;
      33843: inst = 32'h8220000;
      33844: inst = 32'h10408000;
      33845: inst = 32'hc4049d8;
      33846: inst = 32'h8220000;
      33847: inst = 32'h10408000;
      33848: inst = 32'hc4049d9;
      33849: inst = 32'h8220000;
      33850: inst = 32'h10408000;
      33851: inst = 32'hc4049da;
      33852: inst = 32'h8220000;
      33853: inst = 32'h10408000;
      33854: inst = 32'hc4049db;
      33855: inst = 32'h8220000;
      33856: inst = 32'h10408000;
      33857: inst = 32'hc4049dc;
      33858: inst = 32'h8220000;
      33859: inst = 32'h10408000;
      33860: inst = 32'hc4049dd;
      33861: inst = 32'h8220000;
      33862: inst = 32'h10408000;
      33863: inst = 32'hc4049de;
      33864: inst = 32'h8220000;
      33865: inst = 32'h10408000;
      33866: inst = 32'hc4049df;
      33867: inst = 32'h8220000;
      33868: inst = 32'h10408000;
      33869: inst = 32'hc4049e0;
      33870: inst = 32'h8220000;
      33871: inst = 32'h10408000;
      33872: inst = 32'hc4049e1;
      33873: inst = 32'h8220000;
      33874: inst = 32'h10408000;
      33875: inst = 32'hc4049e2;
      33876: inst = 32'h8220000;
      33877: inst = 32'h10408000;
      33878: inst = 32'hc4049e3;
      33879: inst = 32'h8220000;
      33880: inst = 32'h10408000;
      33881: inst = 32'hc4049e4;
      33882: inst = 32'h8220000;
      33883: inst = 32'h10408000;
      33884: inst = 32'hc4049e5;
      33885: inst = 32'h8220000;
      33886: inst = 32'h10408000;
      33887: inst = 32'hc4049ef;
      33888: inst = 32'h8220000;
      33889: inst = 32'h10408000;
      33890: inst = 32'hc4049f0;
      33891: inst = 32'h8220000;
      33892: inst = 32'h10408000;
      33893: inst = 32'hc4049f1;
      33894: inst = 32'h8220000;
      33895: inst = 32'h10408000;
      33896: inst = 32'hc4049f2;
      33897: inst = 32'h8220000;
      33898: inst = 32'h10408000;
      33899: inst = 32'hc4049f3;
      33900: inst = 32'h8220000;
      33901: inst = 32'h10408000;
      33902: inst = 32'hc4049f4;
      33903: inst = 32'h8220000;
      33904: inst = 32'h10408000;
      33905: inst = 32'hc4049f5;
      33906: inst = 32'h8220000;
      33907: inst = 32'h10408000;
      33908: inst = 32'hc4049f6;
      33909: inst = 32'h8220000;
      33910: inst = 32'h10408000;
      33911: inst = 32'hc4049f7;
      33912: inst = 32'h8220000;
      33913: inst = 32'h10408000;
      33914: inst = 32'hc4049f8;
      33915: inst = 32'h8220000;
      33916: inst = 32'h10408000;
      33917: inst = 32'hc4049f9;
      33918: inst = 32'h8220000;
      33919: inst = 32'h10408000;
      33920: inst = 32'hc4049fa;
      33921: inst = 32'h8220000;
      33922: inst = 32'h10408000;
      33923: inst = 32'hc4049fb;
      33924: inst = 32'h8220000;
      33925: inst = 32'h10408000;
      33926: inst = 32'hc4049fc;
      33927: inst = 32'h8220000;
      33928: inst = 32'h10408000;
      33929: inst = 32'hc404a03;
      33930: inst = 32'h8220000;
      33931: inst = 32'h10408000;
      33932: inst = 32'hc404a04;
      33933: inst = 32'h8220000;
      33934: inst = 32'h10408000;
      33935: inst = 32'hc404a05;
      33936: inst = 32'h8220000;
      33937: inst = 32'h10408000;
      33938: inst = 32'hc404a06;
      33939: inst = 32'h8220000;
      33940: inst = 32'h10408000;
      33941: inst = 32'hc404a07;
      33942: inst = 32'h8220000;
      33943: inst = 32'h10408000;
      33944: inst = 32'hc404a08;
      33945: inst = 32'h8220000;
      33946: inst = 32'h10408000;
      33947: inst = 32'hc404a09;
      33948: inst = 32'h8220000;
      33949: inst = 32'h10408000;
      33950: inst = 32'hc404a0a;
      33951: inst = 32'h8220000;
      33952: inst = 32'h10408000;
      33953: inst = 32'hc404a0b;
      33954: inst = 32'h8220000;
      33955: inst = 32'h10408000;
      33956: inst = 32'hc404a0c;
      33957: inst = 32'h8220000;
      33958: inst = 32'h10408000;
      33959: inst = 32'hc404a0d;
      33960: inst = 32'h8220000;
      33961: inst = 32'h10408000;
      33962: inst = 32'hc404a11;
      33963: inst = 32'h8220000;
      33964: inst = 32'h10408000;
      33965: inst = 32'hc404a12;
      33966: inst = 32'h8220000;
      33967: inst = 32'h10408000;
      33968: inst = 32'hc404a13;
      33969: inst = 32'h8220000;
      33970: inst = 32'h10408000;
      33971: inst = 32'hc404a14;
      33972: inst = 32'h8220000;
      33973: inst = 32'h10408000;
      33974: inst = 32'hc404a15;
      33975: inst = 32'h8220000;
      33976: inst = 32'h10408000;
      33977: inst = 32'hc404a16;
      33978: inst = 32'h8220000;
      33979: inst = 32'h10408000;
      33980: inst = 32'hc404a17;
      33981: inst = 32'h8220000;
      33982: inst = 32'h10408000;
      33983: inst = 32'hc404a18;
      33984: inst = 32'h8220000;
      33985: inst = 32'h10408000;
      33986: inst = 32'hc404a19;
      33987: inst = 32'h8220000;
      33988: inst = 32'h10408000;
      33989: inst = 32'hc404a1a;
      33990: inst = 32'h8220000;
      33991: inst = 32'h10408000;
      33992: inst = 32'hc404a1b;
      33993: inst = 32'h8220000;
      33994: inst = 32'h10408000;
      33995: inst = 32'hc404a1c;
      33996: inst = 32'h8220000;
      33997: inst = 32'h10408000;
      33998: inst = 32'hc404a1d;
      33999: inst = 32'h8220000;
      34000: inst = 32'h10408000;
      34001: inst = 32'hc404a1e;
      34002: inst = 32'h8220000;
      34003: inst = 32'h10408000;
      34004: inst = 32'hc404a1f;
      34005: inst = 32'h8220000;
      34006: inst = 32'h10408000;
      34007: inst = 32'hc404a20;
      34008: inst = 32'h8220000;
      34009: inst = 32'h10408000;
      34010: inst = 32'hc404a21;
      34011: inst = 32'h8220000;
      34012: inst = 32'h10408000;
      34013: inst = 32'hc404a22;
      34014: inst = 32'h8220000;
      34015: inst = 32'h10408000;
      34016: inst = 32'hc404a23;
      34017: inst = 32'h8220000;
      34018: inst = 32'h10408000;
      34019: inst = 32'hc404a24;
      34020: inst = 32'h8220000;
      34021: inst = 32'h10408000;
      34022: inst = 32'hc404a25;
      34023: inst = 32'h8220000;
      34024: inst = 32'h10408000;
      34025: inst = 32'hc404a26;
      34026: inst = 32'h8220000;
      34027: inst = 32'h10408000;
      34028: inst = 32'hc404a27;
      34029: inst = 32'h8220000;
      34030: inst = 32'h10408000;
      34031: inst = 32'hc404a28;
      34032: inst = 32'h8220000;
      34033: inst = 32'h10408000;
      34034: inst = 32'hc404a29;
      34035: inst = 32'h8220000;
      34036: inst = 32'h10408000;
      34037: inst = 32'hc404a2a;
      34038: inst = 32'h8220000;
      34039: inst = 32'h10408000;
      34040: inst = 32'hc404a2b;
      34041: inst = 32'h8220000;
      34042: inst = 32'h10408000;
      34043: inst = 32'hc404a2c;
      34044: inst = 32'h8220000;
      34045: inst = 32'h10408000;
      34046: inst = 32'hc404a2d;
      34047: inst = 32'h8220000;
      34048: inst = 32'h10408000;
      34049: inst = 32'hc404a2e;
      34050: inst = 32'h8220000;
      34051: inst = 32'h10408000;
      34052: inst = 32'hc404a2f;
      34053: inst = 32'h8220000;
      34054: inst = 32'h10408000;
      34055: inst = 32'hc404a30;
      34056: inst = 32'h8220000;
      34057: inst = 32'h10408000;
      34058: inst = 32'hc404a31;
      34059: inst = 32'h8220000;
      34060: inst = 32'h10408000;
      34061: inst = 32'hc404a32;
      34062: inst = 32'h8220000;
      34063: inst = 32'h10408000;
      34064: inst = 32'hc404a33;
      34065: inst = 32'h8220000;
      34066: inst = 32'h10408000;
      34067: inst = 32'hc404a34;
      34068: inst = 32'h8220000;
      34069: inst = 32'h10408000;
      34070: inst = 32'hc404a35;
      34071: inst = 32'h8220000;
      34072: inst = 32'h10408000;
      34073: inst = 32'hc404a36;
      34074: inst = 32'h8220000;
      34075: inst = 32'h10408000;
      34076: inst = 32'hc404a37;
      34077: inst = 32'h8220000;
      34078: inst = 32'h10408000;
      34079: inst = 32'hc404a38;
      34080: inst = 32'h8220000;
      34081: inst = 32'h10408000;
      34082: inst = 32'hc404a39;
      34083: inst = 32'h8220000;
      34084: inst = 32'h10408000;
      34085: inst = 32'hc404a3a;
      34086: inst = 32'h8220000;
      34087: inst = 32'h10408000;
      34088: inst = 32'hc404a3b;
      34089: inst = 32'h8220000;
      34090: inst = 32'h10408000;
      34091: inst = 32'hc404a3c;
      34092: inst = 32'h8220000;
      34093: inst = 32'h10408000;
      34094: inst = 32'hc404a3d;
      34095: inst = 32'h8220000;
      34096: inst = 32'h10408000;
      34097: inst = 32'hc404a3e;
      34098: inst = 32'h8220000;
      34099: inst = 32'h10408000;
      34100: inst = 32'hc404a3f;
      34101: inst = 32'h8220000;
      34102: inst = 32'h10408000;
      34103: inst = 32'hc404a40;
      34104: inst = 32'h8220000;
      34105: inst = 32'h10408000;
      34106: inst = 32'hc404a41;
      34107: inst = 32'h8220000;
      34108: inst = 32'h10408000;
      34109: inst = 32'hc404a42;
      34110: inst = 32'h8220000;
      34111: inst = 32'h10408000;
      34112: inst = 32'hc404a43;
      34113: inst = 32'h8220000;
      34114: inst = 32'h10408000;
      34115: inst = 32'hc404a44;
      34116: inst = 32'h8220000;
      34117: inst = 32'h10408000;
      34118: inst = 32'hc404a45;
      34119: inst = 32'h8220000;
      34120: inst = 32'h10408000;
      34121: inst = 32'hc404a4f;
      34122: inst = 32'h8220000;
      34123: inst = 32'h10408000;
      34124: inst = 32'hc404a50;
      34125: inst = 32'h8220000;
      34126: inst = 32'h10408000;
      34127: inst = 32'hc404a51;
      34128: inst = 32'h8220000;
      34129: inst = 32'h10408000;
      34130: inst = 32'hc404a52;
      34131: inst = 32'h8220000;
      34132: inst = 32'h10408000;
      34133: inst = 32'hc404a53;
      34134: inst = 32'h8220000;
      34135: inst = 32'h10408000;
      34136: inst = 32'hc404a54;
      34137: inst = 32'h8220000;
      34138: inst = 32'h10408000;
      34139: inst = 32'hc404a55;
      34140: inst = 32'h8220000;
      34141: inst = 32'h10408000;
      34142: inst = 32'hc404a56;
      34143: inst = 32'h8220000;
      34144: inst = 32'h10408000;
      34145: inst = 32'hc404a57;
      34146: inst = 32'h8220000;
      34147: inst = 32'h10408000;
      34148: inst = 32'hc404a58;
      34149: inst = 32'h8220000;
      34150: inst = 32'h10408000;
      34151: inst = 32'hc404a59;
      34152: inst = 32'h8220000;
      34153: inst = 32'h10408000;
      34154: inst = 32'hc404a5a;
      34155: inst = 32'h8220000;
      34156: inst = 32'h10408000;
      34157: inst = 32'hc404a5b;
      34158: inst = 32'h8220000;
      34159: inst = 32'h10408000;
      34160: inst = 32'hc404a5c;
      34161: inst = 32'h8220000;
      34162: inst = 32'h10408000;
      34163: inst = 32'hc404a63;
      34164: inst = 32'h8220000;
      34165: inst = 32'h10408000;
      34166: inst = 32'hc404a64;
      34167: inst = 32'h8220000;
      34168: inst = 32'h10408000;
      34169: inst = 32'hc404a65;
      34170: inst = 32'h8220000;
      34171: inst = 32'h10408000;
      34172: inst = 32'hc404a66;
      34173: inst = 32'h8220000;
      34174: inst = 32'h10408000;
      34175: inst = 32'hc404a67;
      34176: inst = 32'h8220000;
      34177: inst = 32'h10408000;
      34178: inst = 32'hc404a68;
      34179: inst = 32'h8220000;
      34180: inst = 32'h10408000;
      34181: inst = 32'hc404a69;
      34182: inst = 32'h8220000;
      34183: inst = 32'h10408000;
      34184: inst = 32'hc404a6a;
      34185: inst = 32'h8220000;
      34186: inst = 32'h10408000;
      34187: inst = 32'hc404a6b;
      34188: inst = 32'h8220000;
      34189: inst = 32'h10408000;
      34190: inst = 32'hc404a6c;
      34191: inst = 32'h8220000;
      34192: inst = 32'h10408000;
      34193: inst = 32'hc404a6d;
      34194: inst = 32'h8220000;
      34195: inst = 32'h10408000;
      34196: inst = 32'hc404a71;
      34197: inst = 32'h8220000;
      34198: inst = 32'h10408000;
      34199: inst = 32'hc404a72;
      34200: inst = 32'h8220000;
      34201: inst = 32'h10408000;
      34202: inst = 32'hc404a73;
      34203: inst = 32'h8220000;
      34204: inst = 32'h10408000;
      34205: inst = 32'hc404a74;
      34206: inst = 32'h8220000;
      34207: inst = 32'h10408000;
      34208: inst = 32'hc404a75;
      34209: inst = 32'h8220000;
      34210: inst = 32'h10408000;
      34211: inst = 32'hc404a76;
      34212: inst = 32'h8220000;
      34213: inst = 32'h10408000;
      34214: inst = 32'hc404a77;
      34215: inst = 32'h8220000;
      34216: inst = 32'h10408000;
      34217: inst = 32'hc404a78;
      34218: inst = 32'h8220000;
      34219: inst = 32'h10408000;
      34220: inst = 32'hc404a79;
      34221: inst = 32'h8220000;
      34222: inst = 32'h10408000;
      34223: inst = 32'hc404a7a;
      34224: inst = 32'h8220000;
      34225: inst = 32'h10408000;
      34226: inst = 32'hc404a7b;
      34227: inst = 32'h8220000;
      34228: inst = 32'h10408000;
      34229: inst = 32'hc404a7c;
      34230: inst = 32'h8220000;
      34231: inst = 32'h10408000;
      34232: inst = 32'hc404a7d;
      34233: inst = 32'h8220000;
      34234: inst = 32'h10408000;
      34235: inst = 32'hc404a7e;
      34236: inst = 32'h8220000;
      34237: inst = 32'h10408000;
      34238: inst = 32'hc404a7f;
      34239: inst = 32'h8220000;
      34240: inst = 32'h10408000;
      34241: inst = 32'hc404a80;
      34242: inst = 32'h8220000;
      34243: inst = 32'h10408000;
      34244: inst = 32'hc404a81;
      34245: inst = 32'h8220000;
      34246: inst = 32'h10408000;
      34247: inst = 32'hc404a82;
      34248: inst = 32'h8220000;
      34249: inst = 32'h10408000;
      34250: inst = 32'hc404a83;
      34251: inst = 32'h8220000;
      34252: inst = 32'h10408000;
      34253: inst = 32'hc404a84;
      34254: inst = 32'h8220000;
      34255: inst = 32'h10408000;
      34256: inst = 32'hc404a85;
      34257: inst = 32'h8220000;
      34258: inst = 32'h10408000;
      34259: inst = 32'hc404a86;
      34260: inst = 32'h8220000;
      34261: inst = 32'h10408000;
      34262: inst = 32'hc404a87;
      34263: inst = 32'h8220000;
      34264: inst = 32'h10408000;
      34265: inst = 32'hc404a88;
      34266: inst = 32'h8220000;
      34267: inst = 32'h10408000;
      34268: inst = 32'hc404a89;
      34269: inst = 32'h8220000;
      34270: inst = 32'h10408000;
      34271: inst = 32'hc404a8a;
      34272: inst = 32'h8220000;
      34273: inst = 32'h10408000;
      34274: inst = 32'hc404a8b;
      34275: inst = 32'h8220000;
      34276: inst = 32'h10408000;
      34277: inst = 32'hc404a8c;
      34278: inst = 32'h8220000;
      34279: inst = 32'h10408000;
      34280: inst = 32'hc404a8d;
      34281: inst = 32'h8220000;
      34282: inst = 32'h10408000;
      34283: inst = 32'hc404a8e;
      34284: inst = 32'h8220000;
      34285: inst = 32'h10408000;
      34286: inst = 32'hc404a8f;
      34287: inst = 32'h8220000;
      34288: inst = 32'h10408000;
      34289: inst = 32'hc404a90;
      34290: inst = 32'h8220000;
      34291: inst = 32'h10408000;
      34292: inst = 32'hc404a91;
      34293: inst = 32'h8220000;
      34294: inst = 32'h10408000;
      34295: inst = 32'hc404a92;
      34296: inst = 32'h8220000;
      34297: inst = 32'h10408000;
      34298: inst = 32'hc404a93;
      34299: inst = 32'h8220000;
      34300: inst = 32'h10408000;
      34301: inst = 32'hc404a94;
      34302: inst = 32'h8220000;
      34303: inst = 32'h10408000;
      34304: inst = 32'hc404a95;
      34305: inst = 32'h8220000;
      34306: inst = 32'h10408000;
      34307: inst = 32'hc404a96;
      34308: inst = 32'h8220000;
      34309: inst = 32'h10408000;
      34310: inst = 32'hc404a97;
      34311: inst = 32'h8220000;
      34312: inst = 32'h10408000;
      34313: inst = 32'hc404a98;
      34314: inst = 32'h8220000;
      34315: inst = 32'h10408000;
      34316: inst = 32'hc404a99;
      34317: inst = 32'h8220000;
      34318: inst = 32'h10408000;
      34319: inst = 32'hc404a9a;
      34320: inst = 32'h8220000;
      34321: inst = 32'h10408000;
      34322: inst = 32'hc404a9b;
      34323: inst = 32'h8220000;
      34324: inst = 32'h10408000;
      34325: inst = 32'hc404a9c;
      34326: inst = 32'h8220000;
      34327: inst = 32'h10408000;
      34328: inst = 32'hc404a9d;
      34329: inst = 32'h8220000;
      34330: inst = 32'h10408000;
      34331: inst = 32'hc404a9e;
      34332: inst = 32'h8220000;
      34333: inst = 32'h10408000;
      34334: inst = 32'hc404a9f;
      34335: inst = 32'h8220000;
      34336: inst = 32'h10408000;
      34337: inst = 32'hc404aa0;
      34338: inst = 32'h8220000;
      34339: inst = 32'h10408000;
      34340: inst = 32'hc404aa1;
      34341: inst = 32'h8220000;
      34342: inst = 32'h10408000;
      34343: inst = 32'hc404aa2;
      34344: inst = 32'h8220000;
      34345: inst = 32'h10408000;
      34346: inst = 32'hc404aa3;
      34347: inst = 32'h8220000;
      34348: inst = 32'h10408000;
      34349: inst = 32'hc404aa4;
      34350: inst = 32'h8220000;
      34351: inst = 32'h10408000;
      34352: inst = 32'hc404aa5;
      34353: inst = 32'h8220000;
      34354: inst = 32'h10408000;
      34355: inst = 32'hc404aa6;
      34356: inst = 32'h8220000;
      34357: inst = 32'h10408000;
      34358: inst = 32'hc404aa7;
      34359: inst = 32'h8220000;
      34360: inst = 32'h10408000;
      34361: inst = 32'hc404aa8;
      34362: inst = 32'h8220000;
      34363: inst = 32'h10408000;
      34364: inst = 32'hc404aa9;
      34365: inst = 32'h8220000;
      34366: inst = 32'h10408000;
      34367: inst = 32'hc404aaa;
      34368: inst = 32'h8220000;
      34369: inst = 32'h10408000;
      34370: inst = 32'hc404aab;
      34371: inst = 32'h8220000;
      34372: inst = 32'h10408000;
      34373: inst = 32'hc404aac;
      34374: inst = 32'h8220000;
      34375: inst = 32'h10408000;
      34376: inst = 32'hc404aad;
      34377: inst = 32'h8220000;
      34378: inst = 32'h10408000;
      34379: inst = 32'hc404aae;
      34380: inst = 32'h8220000;
      34381: inst = 32'h10408000;
      34382: inst = 32'hc404aaf;
      34383: inst = 32'h8220000;
      34384: inst = 32'h10408000;
      34385: inst = 32'hc404ab0;
      34386: inst = 32'h8220000;
      34387: inst = 32'h10408000;
      34388: inst = 32'hc404ab1;
      34389: inst = 32'h8220000;
      34390: inst = 32'h10408000;
      34391: inst = 32'hc404ab2;
      34392: inst = 32'h8220000;
      34393: inst = 32'h10408000;
      34394: inst = 32'hc404ab3;
      34395: inst = 32'h8220000;
      34396: inst = 32'h10408000;
      34397: inst = 32'hc404ab4;
      34398: inst = 32'h8220000;
      34399: inst = 32'h10408000;
      34400: inst = 32'hc404ab5;
      34401: inst = 32'h8220000;
      34402: inst = 32'h10408000;
      34403: inst = 32'hc404ab6;
      34404: inst = 32'h8220000;
      34405: inst = 32'h10408000;
      34406: inst = 32'hc404ab7;
      34407: inst = 32'h8220000;
      34408: inst = 32'h10408000;
      34409: inst = 32'hc404ab8;
      34410: inst = 32'h8220000;
      34411: inst = 32'h10408000;
      34412: inst = 32'hc404ab9;
      34413: inst = 32'h8220000;
      34414: inst = 32'h10408000;
      34415: inst = 32'hc404aba;
      34416: inst = 32'h8220000;
      34417: inst = 32'h10408000;
      34418: inst = 32'hc404abb;
      34419: inst = 32'h8220000;
      34420: inst = 32'h10408000;
      34421: inst = 32'hc404abc;
      34422: inst = 32'h8220000;
      34423: inst = 32'h10408000;
      34424: inst = 32'hc404ac3;
      34425: inst = 32'h8220000;
      34426: inst = 32'h10408000;
      34427: inst = 32'hc404ac4;
      34428: inst = 32'h8220000;
      34429: inst = 32'h10408000;
      34430: inst = 32'hc404ac5;
      34431: inst = 32'h8220000;
      34432: inst = 32'h10408000;
      34433: inst = 32'hc404ac6;
      34434: inst = 32'h8220000;
      34435: inst = 32'h10408000;
      34436: inst = 32'hc404ac7;
      34437: inst = 32'h8220000;
      34438: inst = 32'h10408000;
      34439: inst = 32'hc404ac8;
      34440: inst = 32'h8220000;
      34441: inst = 32'h10408000;
      34442: inst = 32'hc404ac9;
      34443: inst = 32'h8220000;
      34444: inst = 32'h10408000;
      34445: inst = 32'hc404aca;
      34446: inst = 32'h8220000;
      34447: inst = 32'h10408000;
      34448: inst = 32'hc404acb;
      34449: inst = 32'h8220000;
      34450: inst = 32'h10408000;
      34451: inst = 32'hc404acc;
      34452: inst = 32'h8220000;
      34453: inst = 32'h10408000;
      34454: inst = 32'hc404acd;
      34455: inst = 32'h8220000;
      34456: inst = 32'h10408000;
      34457: inst = 32'hc404ad1;
      34458: inst = 32'h8220000;
      34459: inst = 32'h10408000;
      34460: inst = 32'hc404ad2;
      34461: inst = 32'h8220000;
      34462: inst = 32'h10408000;
      34463: inst = 32'hc404ad3;
      34464: inst = 32'h8220000;
      34465: inst = 32'h10408000;
      34466: inst = 32'hc404ad4;
      34467: inst = 32'h8220000;
      34468: inst = 32'h10408000;
      34469: inst = 32'hc404ad5;
      34470: inst = 32'h8220000;
      34471: inst = 32'h10408000;
      34472: inst = 32'hc404ad6;
      34473: inst = 32'h8220000;
      34474: inst = 32'h10408000;
      34475: inst = 32'hc404ad7;
      34476: inst = 32'h8220000;
      34477: inst = 32'h10408000;
      34478: inst = 32'hc404ad8;
      34479: inst = 32'h8220000;
      34480: inst = 32'h10408000;
      34481: inst = 32'hc404ad9;
      34482: inst = 32'h8220000;
      34483: inst = 32'h10408000;
      34484: inst = 32'hc404ada;
      34485: inst = 32'h8220000;
      34486: inst = 32'h10408000;
      34487: inst = 32'hc404adb;
      34488: inst = 32'h8220000;
      34489: inst = 32'h10408000;
      34490: inst = 32'hc404adc;
      34491: inst = 32'h8220000;
      34492: inst = 32'h10408000;
      34493: inst = 32'hc404add;
      34494: inst = 32'h8220000;
      34495: inst = 32'h10408000;
      34496: inst = 32'hc404ade;
      34497: inst = 32'h8220000;
      34498: inst = 32'h10408000;
      34499: inst = 32'hc404adf;
      34500: inst = 32'h8220000;
      34501: inst = 32'h10408000;
      34502: inst = 32'hc404ae0;
      34503: inst = 32'h8220000;
      34504: inst = 32'h10408000;
      34505: inst = 32'hc404ae1;
      34506: inst = 32'h8220000;
      34507: inst = 32'h10408000;
      34508: inst = 32'hc404ae2;
      34509: inst = 32'h8220000;
      34510: inst = 32'h10408000;
      34511: inst = 32'hc404ae3;
      34512: inst = 32'h8220000;
      34513: inst = 32'h10408000;
      34514: inst = 32'hc404ae4;
      34515: inst = 32'h8220000;
      34516: inst = 32'h10408000;
      34517: inst = 32'hc404ae5;
      34518: inst = 32'h8220000;
      34519: inst = 32'h10408000;
      34520: inst = 32'hc404ae6;
      34521: inst = 32'h8220000;
      34522: inst = 32'h10408000;
      34523: inst = 32'hc404ae7;
      34524: inst = 32'h8220000;
      34525: inst = 32'h10408000;
      34526: inst = 32'hc404ae8;
      34527: inst = 32'h8220000;
      34528: inst = 32'h10408000;
      34529: inst = 32'hc404ae9;
      34530: inst = 32'h8220000;
      34531: inst = 32'h10408000;
      34532: inst = 32'hc404aea;
      34533: inst = 32'h8220000;
      34534: inst = 32'h10408000;
      34535: inst = 32'hc404aeb;
      34536: inst = 32'h8220000;
      34537: inst = 32'h10408000;
      34538: inst = 32'hc404aec;
      34539: inst = 32'h8220000;
      34540: inst = 32'h10408000;
      34541: inst = 32'hc404aed;
      34542: inst = 32'h8220000;
      34543: inst = 32'h10408000;
      34544: inst = 32'hc404aee;
      34545: inst = 32'h8220000;
      34546: inst = 32'h10408000;
      34547: inst = 32'hc404aef;
      34548: inst = 32'h8220000;
      34549: inst = 32'h10408000;
      34550: inst = 32'hc404af0;
      34551: inst = 32'h8220000;
      34552: inst = 32'h10408000;
      34553: inst = 32'hc404af1;
      34554: inst = 32'h8220000;
      34555: inst = 32'h10408000;
      34556: inst = 32'hc404af2;
      34557: inst = 32'h8220000;
      34558: inst = 32'h10408000;
      34559: inst = 32'hc404af3;
      34560: inst = 32'h8220000;
      34561: inst = 32'h10408000;
      34562: inst = 32'hc404af4;
      34563: inst = 32'h8220000;
      34564: inst = 32'h10408000;
      34565: inst = 32'hc404af5;
      34566: inst = 32'h8220000;
      34567: inst = 32'h10408000;
      34568: inst = 32'hc404af6;
      34569: inst = 32'h8220000;
      34570: inst = 32'h10408000;
      34571: inst = 32'hc404af7;
      34572: inst = 32'h8220000;
      34573: inst = 32'h10408000;
      34574: inst = 32'hc404af8;
      34575: inst = 32'h8220000;
      34576: inst = 32'h10408000;
      34577: inst = 32'hc404af9;
      34578: inst = 32'h8220000;
      34579: inst = 32'h10408000;
      34580: inst = 32'hc404afa;
      34581: inst = 32'h8220000;
      34582: inst = 32'h10408000;
      34583: inst = 32'hc404afb;
      34584: inst = 32'h8220000;
      34585: inst = 32'h10408000;
      34586: inst = 32'hc404afc;
      34587: inst = 32'h8220000;
      34588: inst = 32'h10408000;
      34589: inst = 32'hc404afd;
      34590: inst = 32'h8220000;
      34591: inst = 32'h10408000;
      34592: inst = 32'hc404afe;
      34593: inst = 32'h8220000;
      34594: inst = 32'h10408000;
      34595: inst = 32'hc404aff;
      34596: inst = 32'h8220000;
      34597: inst = 32'h10408000;
      34598: inst = 32'hc404b00;
      34599: inst = 32'h8220000;
      34600: inst = 32'h10408000;
      34601: inst = 32'hc404b01;
      34602: inst = 32'h8220000;
      34603: inst = 32'h10408000;
      34604: inst = 32'hc404b02;
      34605: inst = 32'h8220000;
      34606: inst = 32'h10408000;
      34607: inst = 32'hc404b03;
      34608: inst = 32'h8220000;
      34609: inst = 32'h10408000;
      34610: inst = 32'hc404b04;
      34611: inst = 32'h8220000;
      34612: inst = 32'h10408000;
      34613: inst = 32'hc404b05;
      34614: inst = 32'h8220000;
      34615: inst = 32'h10408000;
      34616: inst = 32'hc404b06;
      34617: inst = 32'h8220000;
      34618: inst = 32'h10408000;
      34619: inst = 32'hc404b07;
      34620: inst = 32'h8220000;
      34621: inst = 32'h10408000;
      34622: inst = 32'hc404b08;
      34623: inst = 32'h8220000;
      34624: inst = 32'h10408000;
      34625: inst = 32'hc404b09;
      34626: inst = 32'h8220000;
      34627: inst = 32'h10408000;
      34628: inst = 32'hc404b0a;
      34629: inst = 32'h8220000;
      34630: inst = 32'h10408000;
      34631: inst = 32'hc404b0b;
      34632: inst = 32'h8220000;
      34633: inst = 32'h10408000;
      34634: inst = 32'hc404b0c;
      34635: inst = 32'h8220000;
      34636: inst = 32'h10408000;
      34637: inst = 32'hc404b0d;
      34638: inst = 32'h8220000;
      34639: inst = 32'h10408000;
      34640: inst = 32'hc404b0e;
      34641: inst = 32'h8220000;
      34642: inst = 32'h10408000;
      34643: inst = 32'hc404b0f;
      34644: inst = 32'h8220000;
      34645: inst = 32'h10408000;
      34646: inst = 32'hc404b10;
      34647: inst = 32'h8220000;
      34648: inst = 32'h10408000;
      34649: inst = 32'hc404b11;
      34650: inst = 32'h8220000;
      34651: inst = 32'h10408000;
      34652: inst = 32'hc404b12;
      34653: inst = 32'h8220000;
      34654: inst = 32'h10408000;
      34655: inst = 32'hc404b13;
      34656: inst = 32'h8220000;
      34657: inst = 32'h10408000;
      34658: inst = 32'hc404b14;
      34659: inst = 32'h8220000;
      34660: inst = 32'h10408000;
      34661: inst = 32'hc404b15;
      34662: inst = 32'h8220000;
      34663: inst = 32'h10408000;
      34664: inst = 32'hc404b16;
      34665: inst = 32'h8220000;
      34666: inst = 32'h10408000;
      34667: inst = 32'hc404b17;
      34668: inst = 32'h8220000;
      34669: inst = 32'h10408000;
      34670: inst = 32'hc404b18;
      34671: inst = 32'h8220000;
      34672: inst = 32'h10408000;
      34673: inst = 32'hc404b19;
      34674: inst = 32'h8220000;
      34675: inst = 32'h10408000;
      34676: inst = 32'hc404b1a;
      34677: inst = 32'h8220000;
      34678: inst = 32'h10408000;
      34679: inst = 32'hc404b1b;
      34680: inst = 32'h8220000;
      34681: inst = 32'h10408000;
      34682: inst = 32'hc404b1c;
      34683: inst = 32'h8220000;
      34684: inst = 32'h10408000;
      34685: inst = 32'hc404b31;
      34686: inst = 32'h8220000;
      34687: inst = 32'h10408000;
      34688: inst = 32'hc404b32;
      34689: inst = 32'h8220000;
      34690: inst = 32'h10408000;
      34691: inst = 32'hc404b33;
      34692: inst = 32'h8220000;
      34693: inst = 32'h10408000;
      34694: inst = 32'hc404b34;
      34695: inst = 32'h8220000;
      34696: inst = 32'h10408000;
      34697: inst = 32'hc404b35;
      34698: inst = 32'h8220000;
      34699: inst = 32'h10408000;
      34700: inst = 32'hc404b36;
      34701: inst = 32'h8220000;
      34702: inst = 32'h10408000;
      34703: inst = 32'hc404b37;
      34704: inst = 32'h8220000;
      34705: inst = 32'h10408000;
      34706: inst = 32'hc404b38;
      34707: inst = 32'h8220000;
      34708: inst = 32'h10408000;
      34709: inst = 32'hc404b39;
      34710: inst = 32'h8220000;
      34711: inst = 32'h10408000;
      34712: inst = 32'hc404b3a;
      34713: inst = 32'h8220000;
      34714: inst = 32'h10408000;
      34715: inst = 32'hc404b3b;
      34716: inst = 32'h8220000;
      34717: inst = 32'h10408000;
      34718: inst = 32'hc404b3c;
      34719: inst = 32'h8220000;
      34720: inst = 32'h10408000;
      34721: inst = 32'hc404b3d;
      34722: inst = 32'h8220000;
      34723: inst = 32'h10408000;
      34724: inst = 32'hc404b3e;
      34725: inst = 32'h8220000;
      34726: inst = 32'h10408000;
      34727: inst = 32'hc404b3f;
      34728: inst = 32'h8220000;
      34729: inst = 32'h10408000;
      34730: inst = 32'hc404b40;
      34731: inst = 32'h8220000;
      34732: inst = 32'h10408000;
      34733: inst = 32'hc404b41;
      34734: inst = 32'h8220000;
      34735: inst = 32'h10408000;
      34736: inst = 32'hc404b42;
      34737: inst = 32'h8220000;
      34738: inst = 32'h10408000;
      34739: inst = 32'hc404b43;
      34740: inst = 32'h8220000;
      34741: inst = 32'h10408000;
      34742: inst = 32'hc404b44;
      34743: inst = 32'h8220000;
      34744: inst = 32'h10408000;
      34745: inst = 32'hc404b45;
      34746: inst = 32'h8220000;
      34747: inst = 32'h10408000;
      34748: inst = 32'hc404b46;
      34749: inst = 32'h8220000;
      34750: inst = 32'h10408000;
      34751: inst = 32'hc404b47;
      34752: inst = 32'h8220000;
      34753: inst = 32'h10408000;
      34754: inst = 32'hc404b48;
      34755: inst = 32'h8220000;
      34756: inst = 32'h10408000;
      34757: inst = 32'hc404b49;
      34758: inst = 32'h8220000;
      34759: inst = 32'h10408000;
      34760: inst = 32'hc404b4a;
      34761: inst = 32'h8220000;
      34762: inst = 32'h10408000;
      34763: inst = 32'hc404b4b;
      34764: inst = 32'h8220000;
      34765: inst = 32'h10408000;
      34766: inst = 32'hc404b4c;
      34767: inst = 32'h8220000;
      34768: inst = 32'h10408000;
      34769: inst = 32'hc404b4d;
      34770: inst = 32'h8220000;
      34771: inst = 32'h10408000;
      34772: inst = 32'hc404b4e;
      34773: inst = 32'h8220000;
      34774: inst = 32'h10408000;
      34775: inst = 32'hc404b4f;
      34776: inst = 32'h8220000;
      34777: inst = 32'h10408000;
      34778: inst = 32'hc404b50;
      34779: inst = 32'h8220000;
      34780: inst = 32'h10408000;
      34781: inst = 32'hc404b51;
      34782: inst = 32'h8220000;
      34783: inst = 32'h10408000;
      34784: inst = 32'hc404b52;
      34785: inst = 32'h8220000;
      34786: inst = 32'h10408000;
      34787: inst = 32'hc404b53;
      34788: inst = 32'h8220000;
      34789: inst = 32'h10408000;
      34790: inst = 32'hc404b54;
      34791: inst = 32'h8220000;
      34792: inst = 32'h10408000;
      34793: inst = 32'hc404b55;
      34794: inst = 32'h8220000;
      34795: inst = 32'h10408000;
      34796: inst = 32'hc404b56;
      34797: inst = 32'h8220000;
      34798: inst = 32'h10408000;
      34799: inst = 32'hc404b57;
      34800: inst = 32'h8220000;
      34801: inst = 32'h10408000;
      34802: inst = 32'hc404b58;
      34803: inst = 32'h8220000;
      34804: inst = 32'h10408000;
      34805: inst = 32'hc404b59;
      34806: inst = 32'h8220000;
      34807: inst = 32'h10408000;
      34808: inst = 32'hc404b5a;
      34809: inst = 32'h8220000;
      34810: inst = 32'h10408000;
      34811: inst = 32'hc404b5b;
      34812: inst = 32'h8220000;
      34813: inst = 32'h10408000;
      34814: inst = 32'hc404b5c;
      34815: inst = 32'h8220000;
      34816: inst = 32'h10408000;
      34817: inst = 32'hc404b5d;
      34818: inst = 32'h8220000;
      34819: inst = 32'h10408000;
      34820: inst = 32'hc404b5e;
      34821: inst = 32'h8220000;
      34822: inst = 32'h10408000;
      34823: inst = 32'hc404b5f;
      34824: inst = 32'h8220000;
      34825: inst = 32'h10408000;
      34826: inst = 32'hc404b60;
      34827: inst = 32'h8220000;
      34828: inst = 32'h10408000;
      34829: inst = 32'hc404b61;
      34830: inst = 32'h8220000;
      34831: inst = 32'h10408000;
      34832: inst = 32'hc404b62;
      34833: inst = 32'h8220000;
      34834: inst = 32'h10408000;
      34835: inst = 32'hc404b63;
      34836: inst = 32'h8220000;
      34837: inst = 32'h10408000;
      34838: inst = 32'hc404b64;
      34839: inst = 32'h8220000;
      34840: inst = 32'h10408000;
      34841: inst = 32'hc404b65;
      34842: inst = 32'h8220000;
      34843: inst = 32'h10408000;
      34844: inst = 32'hc404b66;
      34845: inst = 32'h8220000;
      34846: inst = 32'h10408000;
      34847: inst = 32'hc404b67;
      34848: inst = 32'h8220000;
      34849: inst = 32'h10408000;
      34850: inst = 32'hc404b68;
      34851: inst = 32'h8220000;
      34852: inst = 32'h10408000;
      34853: inst = 32'hc404b69;
      34854: inst = 32'h8220000;
      34855: inst = 32'h10408000;
      34856: inst = 32'hc404b6a;
      34857: inst = 32'h8220000;
      34858: inst = 32'h10408000;
      34859: inst = 32'hc404b6b;
      34860: inst = 32'h8220000;
      34861: inst = 32'h10408000;
      34862: inst = 32'hc404b6c;
      34863: inst = 32'h8220000;
      34864: inst = 32'h10408000;
      34865: inst = 32'hc404b6d;
      34866: inst = 32'h8220000;
      34867: inst = 32'h10408000;
      34868: inst = 32'hc404b6e;
      34869: inst = 32'h8220000;
      34870: inst = 32'h10408000;
      34871: inst = 32'hc404b6f;
      34872: inst = 32'h8220000;
      34873: inst = 32'h10408000;
      34874: inst = 32'hc404b70;
      34875: inst = 32'h8220000;
      34876: inst = 32'h10408000;
      34877: inst = 32'hc404b71;
      34878: inst = 32'h8220000;
      34879: inst = 32'h10408000;
      34880: inst = 32'hc404b72;
      34881: inst = 32'h8220000;
      34882: inst = 32'h10408000;
      34883: inst = 32'hc404b73;
      34884: inst = 32'h8220000;
      34885: inst = 32'h10408000;
      34886: inst = 32'hc404b74;
      34887: inst = 32'h8220000;
      34888: inst = 32'h10408000;
      34889: inst = 32'hc404b75;
      34890: inst = 32'h8220000;
      34891: inst = 32'h10408000;
      34892: inst = 32'hc404b76;
      34893: inst = 32'h8220000;
      34894: inst = 32'h10408000;
      34895: inst = 32'hc404b77;
      34896: inst = 32'h8220000;
      34897: inst = 32'h10408000;
      34898: inst = 32'hc404b78;
      34899: inst = 32'h8220000;
      34900: inst = 32'h10408000;
      34901: inst = 32'hc404b79;
      34902: inst = 32'h8220000;
      34903: inst = 32'h10408000;
      34904: inst = 32'hc404b7a;
      34905: inst = 32'h8220000;
      34906: inst = 32'h10408000;
      34907: inst = 32'hc404b7b;
      34908: inst = 32'h8220000;
      34909: inst = 32'h10408000;
      34910: inst = 32'hc404b7c;
      34911: inst = 32'h8220000;
      34912: inst = 32'h10408000;
      34913: inst = 32'hc404b91;
      34914: inst = 32'h8220000;
      34915: inst = 32'h10408000;
      34916: inst = 32'hc404b92;
      34917: inst = 32'h8220000;
      34918: inst = 32'h10408000;
      34919: inst = 32'hc404b93;
      34920: inst = 32'h8220000;
      34921: inst = 32'h10408000;
      34922: inst = 32'hc404b94;
      34923: inst = 32'h8220000;
      34924: inst = 32'h10408000;
      34925: inst = 32'hc404b95;
      34926: inst = 32'h8220000;
      34927: inst = 32'h10408000;
      34928: inst = 32'hc404b96;
      34929: inst = 32'h8220000;
      34930: inst = 32'h10408000;
      34931: inst = 32'hc404b97;
      34932: inst = 32'h8220000;
      34933: inst = 32'h10408000;
      34934: inst = 32'hc404b98;
      34935: inst = 32'h8220000;
      34936: inst = 32'h10408000;
      34937: inst = 32'hc404b99;
      34938: inst = 32'h8220000;
      34939: inst = 32'h10408000;
      34940: inst = 32'hc404b9a;
      34941: inst = 32'h8220000;
      34942: inst = 32'h10408000;
      34943: inst = 32'hc404b9b;
      34944: inst = 32'h8220000;
      34945: inst = 32'h10408000;
      34946: inst = 32'hc404b9c;
      34947: inst = 32'h8220000;
      34948: inst = 32'h10408000;
      34949: inst = 32'hc404b9d;
      34950: inst = 32'h8220000;
      34951: inst = 32'h10408000;
      34952: inst = 32'hc404b9e;
      34953: inst = 32'h8220000;
      34954: inst = 32'h10408000;
      34955: inst = 32'hc404b9f;
      34956: inst = 32'h8220000;
      34957: inst = 32'h10408000;
      34958: inst = 32'hc404ba0;
      34959: inst = 32'h8220000;
      34960: inst = 32'h10408000;
      34961: inst = 32'hc404ba1;
      34962: inst = 32'h8220000;
      34963: inst = 32'h10408000;
      34964: inst = 32'hc404ba2;
      34965: inst = 32'h8220000;
      34966: inst = 32'h10408000;
      34967: inst = 32'hc404ba3;
      34968: inst = 32'h8220000;
      34969: inst = 32'h10408000;
      34970: inst = 32'hc404ba4;
      34971: inst = 32'h8220000;
      34972: inst = 32'h10408000;
      34973: inst = 32'hc404ba5;
      34974: inst = 32'h8220000;
      34975: inst = 32'h10408000;
      34976: inst = 32'hc404ba6;
      34977: inst = 32'h8220000;
      34978: inst = 32'h10408000;
      34979: inst = 32'hc404ba7;
      34980: inst = 32'h8220000;
      34981: inst = 32'h10408000;
      34982: inst = 32'hc404ba8;
      34983: inst = 32'h8220000;
      34984: inst = 32'h10408000;
      34985: inst = 32'hc404ba9;
      34986: inst = 32'h8220000;
      34987: inst = 32'h10408000;
      34988: inst = 32'hc404baa;
      34989: inst = 32'h8220000;
      34990: inst = 32'h10408000;
      34991: inst = 32'hc404bab;
      34992: inst = 32'h8220000;
      34993: inst = 32'h10408000;
      34994: inst = 32'hc404bac;
      34995: inst = 32'h8220000;
      34996: inst = 32'h10408000;
      34997: inst = 32'hc404bad;
      34998: inst = 32'h8220000;
      34999: inst = 32'h10408000;
      35000: inst = 32'hc404bae;
      35001: inst = 32'h8220000;
      35002: inst = 32'h10408000;
      35003: inst = 32'hc404baf;
      35004: inst = 32'h8220000;
      35005: inst = 32'h10408000;
      35006: inst = 32'hc404bb0;
      35007: inst = 32'h8220000;
      35008: inst = 32'h10408000;
      35009: inst = 32'hc404bb1;
      35010: inst = 32'h8220000;
      35011: inst = 32'h10408000;
      35012: inst = 32'hc404bb2;
      35013: inst = 32'h8220000;
      35014: inst = 32'h10408000;
      35015: inst = 32'hc404bb3;
      35016: inst = 32'h8220000;
      35017: inst = 32'h10408000;
      35018: inst = 32'hc404bb4;
      35019: inst = 32'h8220000;
      35020: inst = 32'h10408000;
      35021: inst = 32'hc404bb5;
      35022: inst = 32'h8220000;
      35023: inst = 32'h10408000;
      35024: inst = 32'hc404bb6;
      35025: inst = 32'h8220000;
      35026: inst = 32'h10408000;
      35027: inst = 32'hc404bb7;
      35028: inst = 32'h8220000;
      35029: inst = 32'h10408000;
      35030: inst = 32'hc404bb8;
      35031: inst = 32'h8220000;
      35032: inst = 32'h10408000;
      35033: inst = 32'hc404bb9;
      35034: inst = 32'h8220000;
      35035: inst = 32'h10408000;
      35036: inst = 32'hc404bba;
      35037: inst = 32'h8220000;
      35038: inst = 32'h10408000;
      35039: inst = 32'hc404bbb;
      35040: inst = 32'h8220000;
      35041: inst = 32'h10408000;
      35042: inst = 32'hc404bbc;
      35043: inst = 32'h8220000;
      35044: inst = 32'h10408000;
      35045: inst = 32'hc404bbd;
      35046: inst = 32'h8220000;
      35047: inst = 32'h10408000;
      35048: inst = 32'hc404bbe;
      35049: inst = 32'h8220000;
      35050: inst = 32'h10408000;
      35051: inst = 32'hc404bbf;
      35052: inst = 32'h8220000;
      35053: inst = 32'h10408000;
      35054: inst = 32'hc404bc0;
      35055: inst = 32'h8220000;
      35056: inst = 32'h10408000;
      35057: inst = 32'hc404bc1;
      35058: inst = 32'h8220000;
      35059: inst = 32'h10408000;
      35060: inst = 32'hc404bc2;
      35061: inst = 32'h8220000;
      35062: inst = 32'h10408000;
      35063: inst = 32'hc404bc3;
      35064: inst = 32'h8220000;
      35065: inst = 32'h10408000;
      35066: inst = 32'hc404bc4;
      35067: inst = 32'h8220000;
      35068: inst = 32'h10408000;
      35069: inst = 32'hc404bc5;
      35070: inst = 32'h8220000;
      35071: inst = 32'h10408000;
      35072: inst = 32'hc404bc6;
      35073: inst = 32'h8220000;
      35074: inst = 32'h10408000;
      35075: inst = 32'hc404bc7;
      35076: inst = 32'h8220000;
      35077: inst = 32'h10408000;
      35078: inst = 32'hc404bc8;
      35079: inst = 32'h8220000;
      35080: inst = 32'h10408000;
      35081: inst = 32'hc404bc9;
      35082: inst = 32'h8220000;
      35083: inst = 32'h10408000;
      35084: inst = 32'hc404bca;
      35085: inst = 32'h8220000;
      35086: inst = 32'h10408000;
      35087: inst = 32'hc404bcb;
      35088: inst = 32'h8220000;
      35089: inst = 32'h10408000;
      35090: inst = 32'hc404bcc;
      35091: inst = 32'h8220000;
      35092: inst = 32'h10408000;
      35093: inst = 32'hc404bcd;
      35094: inst = 32'h8220000;
      35095: inst = 32'h10408000;
      35096: inst = 32'hc404bce;
      35097: inst = 32'h8220000;
      35098: inst = 32'h10408000;
      35099: inst = 32'hc404bcf;
      35100: inst = 32'h8220000;
      35101: inst = 32'h10408000;
      35102: inst = 32'hc404bd0;
      35103: inst = 32'h8220000;
      35104: inst = 32'h10408000;
      35105: inst = 32'hc404bd1;
      35106: inst = 32'h8220000;
      35107: inst = 32'h10408000;
      35108: inst = 32'hc404bd2;
      35109: inst = 32'h8220000;
      35110: inst = 32'h10408000;
      35111: inst = 32'hc404bd3;
      35112: inst = 32'h8220000;
      35113: inst = 32'h10408000;
      35114: inst = 32'hc404bd4;
      35115: inst = 32'h8220000;
      35116: inst = 32'h10408000;
      35117: inst = 32'hc404bd5;
      35118: inst = 32'h8220000;
      35119: inst = 32'h10408000;
      35120: inst = 32'hc404bd6;
      35121: inst = 32'h8220000;
      35122: inst = 32'h10408000;
      35123: inst = 32'hc404bd7;
      35124: inst = 32'h8220000;
      35125: inst = 32'h10408000;
      35126: inst = 32'hc404bd8;
      35127: inst = 32'h8220000;
      35128: inst = 32'h10408000;
      35129: inst = 32'hc404bd9;
      35130: inst = 32'h8220000;
      35131: inst = 32'h10408000;
      35132: inst = 32'hc404bda;
      35133: inst = 32'h8220000;
      35134: inst = 32'h10408000;
      35135: inst = 32'hc404bdb;
      35136: inst = 32'h8220000;
      35137: inst = 32'h10408000;
      35138: inst = 32'hc404bdc;
      35139: inst = 32'h8220000;
      35140: inst = 32'h10408000;
      35141: inst = 32'hc404bf1;
      35142: inst = 32'h8220000;
      35143: inst = 32'h10408000;
      35144: inst = 32'hc404bf2;
      35145: inst = 32'h8220000;
      35146: inst = 32'h10408000;
      35147: inst = 32'hc404bf3;
      35148: inst = 32'h8220000;
      35149: inst = 32'h10408000;
      35150: inst = 32'hc404bf4;
      35151: inst = 32'h8220000;
      35152: inst = 32'h10408000;
      35153: inst = 32'hc404bf5;
      35154: inst = 32'h8220000;
      35155: inst = 32'h10408000;
      35156: inst = 32'hc404bf6;
      35157: inst = 32'h8220000;
      35158: inst = 32'h10408000;
      35159: inst = 32'hc404bf7;
      35160: inst = 32'h8220000;
      35161: inst = 32'h10408000;
      35162: inst = 32'hc404bf8;
      35163: inst = 32'h8220000;
      35164: inst = 32'h10408000;
      35165: inst = 32'hc404bf9;
      35166: inst = 32'h8220000;
      35167: inst = 32'h10408000;
      35168: inst = 32'hc404bfa;
      35169: inst = 32'h8220000;
      35170: inst = 32'h10408000;
      35171: inst = 32'hc404bfb;
      35172: inst = 32'h8220000;
      35173: inst = 32'h10408000;
      35174: inst = 32'hc404bfc;
      35175: inst = 32'h8220000;
      35176: inst = 32'h10408000;
      35177: inst = 32'hc404bfd;
      35178: inst = 32'h8220000;
      35179: inst = 32'h10408000;
      35180: inst = 32'hc404bfe;
      35181: inst = 32'h8220000;
      35182: inst = 32'h10408000;
      35183: inst = 32'hc404bff;
      35184: inst = 32'h8220000;
      35185: inst = 32'h10408000;
      35186: inst = 32'hc404c00;
      35187: inst = 32'h8220000;
      35188: inst = 32'h10408000;
      35189: inst = 32'hc404c01;
      35190: inst = 32'h8220000;
      35191: inst = 32'h10408000;
      35192: inst = 32'hc404c02;
      35193: inst = 32'h8220000;
      35194: inst = 32'h10408000;
      35195: inst = 32'hc404c03;
      35196: inst = 32'h8220000;
      35197: inst = 32'h10408000;
      35198: inst = 32'hc404c04;
      35199: inst = 32'h8220000;
      35200: inst = 32'h10408000;
      35201: inst = 32'hc404c05;
      35202: inst = 32'h8220000;
      35203: inst = 32'h10408000;
      35204: inst = 32'hc404c06;
      35205: inst = 32'h8220000;
      35206: inst = 32'h10408000;
      35207: inst = 32'hc404c07;
      35208: inst = 32'h8220000;
      35209: inst = 32'h10408000;
      35210: inst = 32'hc404c08;
      35211: inst = 32'h8220000;
      35212: inst = 32'h10408000;
      35213: inst = 32'hc404c09;
      35214: inst = 32'h8220000;
      35215: inst = 32'h10408000;
      35216: inst = 32'hc404c0a;
      35217: inst = 32'h8220000;
      35218: inst = 32'h10408000;
      35219: inst = 32'hc404c0b;
      35220: inst = 32'h8220000;
      35221: inst = 32'h10408000;
      35222: inst = 32'hc404c0c;
      35223: inst = 32'h8220000;
      35224: inst = 32'h10408000;
      35225: inst = 32'hc404c0d;
      35226: inst = 32'h8220000;
      35227: inst = 32'h10408000;
      35228: inst = 32'hc404c0e;
      35229: inst = 32'h8220000;
      35230: inst = 32'h10408000;
      35231: inst = 32'hc404c0f;
      35232: inst = 32'h8220000;
      35233: inst = 32'h10408000;
      35234: inst = 32'hc404c10;
      35235: inst = 32'h8220000;
      35236: inst = 32'h10408000;
      35237: inst = 32'hc404c11;
      35238: inst = 32'h8220000;
      35239: inst = 32'h10408000;
      35240: inst = 32'hc404c12;
      35241: inst = 32'h8220000;
      35242: inst = 32'h10408000;
      35243: inst = 32'hc404c13;
      35244: inst = 32'h8220000;
      35245: inst = 32'h10408000;
      35246: inst = 32'hc404c14;
      35247: inst = 32'h8220000;
      35248: inst = 32'h10408000;
      35249: inst = 32'hc404c15;
      35250: inst = 32'h8220000;
      35251: inst = 32'h10408000;
      35252: inst = 32'hc404c16;
      35253: inst = 32'h8220000;
      35254: inst = 32'h10408000;
      35255: inst = 32'hc404c17;
      35256: inst = 32'h8220000;
      35257: inst = 32'h10408000;
      35258: inst = 32'hc404c18;
      35259: inst = 32'h8220000;
      35260: inst = 32'h10408000;
      35261: inst = 32'hc404c19;
      35262: inst = 32'h8220000;
      35263: inst = 32'h10408000;
      35264: inst = 32'hc404c1a;
      35265: inst = 32'h8220000;
      35266: inst = 32'h10408000;
      35267: inst = 32'hc404c1b;
      35268: inst = 32'h8220000;
      35269: inst = 32'h10408000;
      35270: inst = 32'hc404c1c;
      35271: inst = 32'h8220000;
      35272: inst = 32'h10408000;
      35273: inst = 32'hc404c1d;
      35274: inst = 32'h8220000;
      35275: inst = 32'h10408000;
      35276: inst = 32'hc404c1e;
      35277: inst = 32'h8220000;
      35278: inst = 32'h10408000;
      35279: inst = 32'hc404c1f;
      35280: inst = 32'h8220000;
      35281: inst = 32'h10408000;
      35282: inst = 32'hc404c20;
      35283: inst = 32'h8220000;
      35284: inst = 32'h10408000;
      35285: inst = 32'hc404c21;
      35286: inst = 32'h8220000;
      35287: inst = 32'h10408000;
      35288: inst = 32'hc404c22;
      35289: inst = 32'h8220000;
      35290: inst = 32'h10408000;
      35291: inst = 32'hc404c23;
      35292: inst = 32'h8220000;
      35293: inst = 32'h10408000;
      35294: inst = 32'hc404c24;
      35295: inst = 32'h8220000;
      35296: inst = 32'h10408000;
      35297: inst = 32'hc404c25;
      35298: inst = 32'h8220000;
      35299: inst = 32'h10408000;
      35300: inst = 32'hc404c26;
      35301: inst = 32'h8220000;
      35302: inst = 32'h10408000;
      35303: inst = 32'hc404c27;
      35304: inst = 32'h8220000;
      35305: inst = 32'h10408000;
      35306: inst = 32'hc404c28;
      35307: inst = 32'h8220000;
      35308: inst = 32'h10408000;
      35309: inst = 32'hc404c29;
      35310: inst = 32'h8220000;
      35311: inst = 32'h10408000;
      35312: inst = 32'hc404c2a;
      35313: inst = 32'h8220000;
      35314: inst = 32'h10408000;
      35315: inst = 32'hc404c2b;
      35316: inst = 32'h8220000;
      35317: inst = 32'h10408000;
      35318: inst = 32'hc404c2c;
      35319: inst = 32'h8220000;
      35320: inst = 32'h10408000;
      35321: inst = 32'hc404c2d;
      35322: inst = 32'h8220000;
      35323: inst = 32'h10408000;
      35324: inst = 32'hc404c2e;
      35325: inst = 32'h8220000;
      35326: inst = 32'h10408000;
      35327: inst = 32'hc404c2f;
      35328: inst = 32'h8220000;
      35329: inst = 32'h10408000;
      35330: inst = 32'hc404c30;
      35331: inst = 32'h8220000;
      35332: inst = 32'h10408000;
      35333: inst = 32'hc404c31;
      35334: inst = 32'h8220000;
      35335: inst = 32'h10408000;
      35336: inst = 32'hc404c32;
      35337: inst = 32'h8220000;
      35338: inst = 32'h10408000;
      35339: inst = 32'hc404c33;
      35340: inst = 32'h8220000;
      35341: inst = 32'h10408000;
      35342: inst = 32'hc404c34;
      35343: inst = 32'h8220000;
      35344: inst = 32'h10408000;
      35345: inst = 32'hc404c35;
      35346: inst = 32'h8220000;
      35347: inst = 32'h10408000;
      35348: inst = 32'hc404c36;
      35349: inst = 32'h8220000;
      35350: inst = 32'h10408000;
      35351: inst = 32'hc404c37;
      35352: inst = 32'h8220000;
      35353: inst = 32'h10408000;
      35354: inst = 32'hc404c38;
      35355: inst = 32'h8220000;
      35356: inst = 32'h10408000;
      35357: inst = 32'hc404c39;
      35358: inst = 32'h8220000;
      35359: inst = 32'h10408000;
      35360: inst = 32'hc404c3a;
      35361: inst = 32'h8220000;
      35362: inst = 32'h10408000;
      35363: inst = 32'hc404c3b;
      35364: inst = 32'h8220000;
      35365: inst = 32'h10408000;
      35366: inst = 32'hc404c3c;
      35367: inst = 32'h8220000;
      35368: inst = 32'h10408000;
      35369: inst = 32'hc404c43;
      35370: inst = 32'h8220000;
      35371: inst = 32'h10408000;
      35372: inst = 32'hc404c44;
      35373: inst = 32'h8220000;
      35374: inst = 32'h10408000;
      35375: inst = 32'hc404c45;
      35376: inst = 32'h8220000;
      35377: inst = 32'h10408000;
      35378: inst = 32'hc404c46;
      35379: inst = 32'h8220000;
      35380: inst = 32'h10408000;
      35381: inst = 32'hc404c47;
      35382: inst = 32'h8220000;
      35383: inst = 32'h10408000;
      35384: inst = 32'hc404c48;
      35385: inst = 32'h8220000;
      35386: inst = 32'h10408000;
      35387: inst = 32'hc404c49;
      35388: inst = 32'h8220000;
      35389: inst = 32'h10408000;
      35390: inst = 32'hc404c4a;
      35391: inst = 32'h8220000;
      35392: inst = 32'h10408000;
      35393: inst = 32'hc404c4b;
      35394: inst = 32'h8220000;
      35395: inst = 32'h10408000;
      35396: inst = 32'hc404c4c;
      35397: inst = 32'h8220000;
      35398: inst = 32'h10408000;
      35399: inst = 32'hc404c4d;
      35400: inst = 32'h8220000;
      35401: inst = 32'h10408000;
      35402: inst = 32'hc404c4e;
      35403: inst = 32'h8220000;
      35404: inst = 32'h10408000;
      35405: inst = 32'hc404c4f;
      35406: inst = 32'h8220000;
      35407: inst = 32'h10408000;
      35408: inst = 32'hc404c50;
      35409: inst = 32'h8220000;
      35410: inst = 32'h10408000;
      35411: inst = 32'hc404c51;
      35412: inst = 32'h8220000;
      35413: inst = 32'h10408000;
      35414: inst = 32'hc404c52;
      35415: inst = 32'h8220000;
      35416: inst = 32'h10408000;
      35417: inst = 32'hc404c53;
      35418: inst = 32'h8220000;
      35419: inst = 32'h10408000;
      35420: inst = 32'hc404c54;
      35421: inst = 32'h8220000;
      35422: inst = 32'h10408000;
      35423: inst = 32'hc404c55;
      35424: inst = 32'h8220000;
      35425: inst = 32'h10408000;
      35426: inst = 32'hc404c56;
      35427: inst = 32'h8220000;
      35428: inst = 32'h10408000;
      35429: inst = 32'hc404c57;
      35430: inst = 32'h8220000;
      35431: inst = 32'h10408000;
      35432: inst = 32'hc404c58;
      35433: inst = 32'h8220000;
      35434: inst = 32'h10408000;
      35435: inst = 32'hc404c59;
      35436: inst = 32'h8220000;
      35437: inst = 32'h10408000;
      35438: inst = 32'hc404c5a;
      35439: inst = 32'h8220000;
      35440: inst = 32'h10408000;
      35441: inst = 32'hc404c5b;
      35442: inst = 32'h8220000;
      35443: inst = 32'h10408000;
      35444: inst = 32'hc404c5c;
      35445: inst = 32'h8220000;
      35446: inst = 32'h10408000;
      35447: inst = 32'hc404c5d;
      35448: inst = 32'h8220000;
      35449: inst = 32'h10408000;
      35450: inst = 32'hc404c5e;
      35451: inst = 32'h8220000;
      35452: inst = 32'h10408000;
      35453: inst = 32'hc404c5f;
      35454: inst = 32'h8220000;
      35455: inst = 32'h10408000;
      35456: inst = 32'hc404c60;
      35457: inst = 32'h8220000;
      35458: inst = 32'h10408000;
      35459: inst = 32'hc404c61;
      35460: inst = 32'h8220000;
      35461: inst = 32'h10408000;
      35462: inst = 32'hc404c62;
      35463: inst = 32'h8220000;
      35464: inst = 32'h10408000;
      35465: inst = 32'hc404c63;
      35466: inst = 32'h8220000;
      35467: inst = 32'h10408000;
      35468: inst = 32'hc404c64;
      35469: inst = 32'h8220000;
      35470: inst = 32'h10408000;
      35471: inst = 32'hc404c65;
      35472: inst = 32'h8220000;
      35473: inst = 32'h10408000;
      35474: inst = 32'hc404c66;
      35475: inst = 32'h8220000;
      35476: inst = 32'h10408000;
      35477: inst = 32'hc404c67;
      35478: inst = 32'h8220000;
      35479: inst = 32'h10408000;
      35480: inst = 32'hc404c68;
      35481: inst = 32'h8220000;
      35482: inst = 32'h10408000;
      35483: inst = 32'hc404c69;
      35484: inst = 32'h8220000;
      35485: inst = 32'h10408000;
      35486: inst = 32'hc404c6a;
      35487: inst = 32'h8220000;
      35488: inst = 32'h10408000;
      35489: inst = 32'hc404c6b;
      35490: inst = 32'h8220000;
      35491: inst = 32'h10408000;
      35492: inst = 32'hc404c6c;
      35493: inst = 32'h8220000;
      35494: inst = 32'h10408000;
      35495: inst = 32'hc404c6d;
      35496: inst = 32'h8220000;
      35497: inst = 32'h10408000;
      35498: inst = 32'hc404c6e;
      35499: inst = 32'h8220000;
      35500: inst = 32'h10408000;
      35501: inst = 32'hc404c6f;
      35502: inst = 32'h8220000;
      35503: inst = 32'h10408000;
      35504: inst = 32'hc404c70;
      35505: inst = 32'h8220000;
      35506: inst = 32'h10408000;
      35507: inst = 32'hc404c71;
      35508: inst = 32'h8220000;
      35509: inst = 32'h10408000;
      35510: inst = 32'hc404c72;
      35511: inst = 32'h8220000;
      35512: inst = 32'h10408000;
      35513: inst = 32'hc404c73;
      35514: inst = 32'h8220000;
      35515: inst = 32'h10408000;
      35516: inst = 32'hc404c74;
      35517: inst = 32'h8220000;
      35518: inst = 32'h10408000;
      35519: inst = 32'hc404c75;
      35520: inst = 32'h8220000;
      35521: inst = 32'h10408000;
      35522: inst = 32'hc404c76;
      35523: inst = 32'h8220000;
      35524: inst = 32'h10408000;
      35525: inst = 32'hc404c77;
      35526: inst = 32'h8220000;
      35527: inst = 32'h10408000;
      35528: inst = 32'hc404c78;
      35529: inst = 32'h8220000;
      35530: inst = 32'h10408000;
      35531: inst = 32'hc404c79;
      35532: inst = 32'h8220000;
      35533: inst = 32'h10408000;
      35534: inst = 32'hc404c7a;
      35535: inst = 32'h8220000;
      35536: inst = 32'h10408000;
      35537: inst = 32'hc404c7b;
      35538: inst = 32'h8220000;
      35539: inst = 32'h10408000;
      35540: inst = 32'hc404c7c;
      35541: inst = 32'h8220000;
      35542: inst = 32'h10408000;
      35543: inst = 32'hc404c7d;
      35544: inst = 32'h8220000;
      35545: inst = 32'h10408000;
      35546: inst = 32'hc404c7e;
      35547: inst = 32'h8220000;
      35548: inst = 32'h10408000;
      35549: inst = 32'hc404c7f;
      35550: inst = 32'h8220000;
      35551: inst = 32'h10408000;
      35552: inst = 32'hc404c80;
      35553: inst = 32'h8220000;
      35554: inst = 32'h10408000;
      35555: inst = 32'hc404c81;
      35556: inst = 32'h8220000;
      35557: inst = 32'h10408000;
      35558: inst = 32'hc404c82;
      35559: inst = 32'h8220000;
      35560: inst = 32'h10408000;
      35561: inst = 32'hc404c83;
      35562: inst = 32'h8220000;
      35563: inst = 32'h10408000;
      35564: inst = 32'hc404c84;
      35565: inst = 32'h8220000;
      35566: inst = 32'h10408000;
      35567: inst = 32'hc404c85;
      35568: inst = 32'h8220000;
      35569: inst = 32'h10408000;
      35570: inst = 32'hc404c86;
      35571: inst = 32'h8220000;
      35572: inst = 32'h10408000;
      35573: inst = 32'hc404c87;
      35574: inst = 32'h8220000;
      35575: inst = 32'h10408000;
      35576: inst = 32'hc404c88;
      35577: inst = 32'h8220000;
      35578: inst = 32'h10408000;
      35579: inst = 32'hc404c89;
      35580: inst = 32'h8220000;
      35581: inst = 32'h10408000;
      35582: inst = 32'hc404c8a;
      35583: inst = 32'h8220000;
      35584: inst = 32'h10408000;
      35585: inst = 32'hc404c8b;
      35586: inst = 32'h8220000;
      35587: inst = 32'h10408000;
      35588: inst = 32'hc404c8c;
      35589: inst = 32'h8220000;
      35590: inst = 32'h10408000;
      35591: inst = 32'hc404c8d;
      35592: inst = 32'h8220000;
      35593: inst = 32'h10408000;
      35594: inst = 32'hc404c8e;
      35595: inst = 32'h8220000;
      35596: inst = 32'h10408000;
      35597: inst = 32'hc404c8f;
      35598: inst = 32'h8220000;
      35599: inst = 32'h10408000;
      35600: inst = 32'hc404c90;
      35601: inst = 32'h8220000;
      35602: inst = 32'h10408000;
      35603: inst = 32'hc404c91;
      35604: inst = 32'h8220000;
      35605: inst = 32'h10408000;
      35606: inst = 32'hc404c92;
      35607: inst = 32'h8220000;
      35608: inst = 32'h10408000;
      35609: inst = 32'hc404c93;
      35610: inst = 32'h8220000;
      35611: inst = 32'h10408000;
      35612: inst = 32'hc404c94;
      35613: inst = 32'h8220000;
      35614: inst = 32'h10408000;
      35615: inst = 32'hc404c95;
      35616: inst = 32'h8220000;
      35617: inst = 32'h10408000;
      35618: inst = 32'hc404c96;
      35619: inst = 32'h8220000;
      35620: inst = 32'h10408000;
      35621: inst = 32'hc404c97;
      35622: inst = 32'h8220000;
      35623: inst = 32'h10408000;
      35624: inst = 32'hc404c98;
      35625: inst = 32'h8220000;
      35626: inst = 32'h10408000;
      35627: inst = 32'hc404c99;
      35628: inst = 32'h8220000;
      35629: inst = 32'h10408000;
      35630: inst = 32'hc404c9a;
      35631: inst = 32'h8220000;
      35632: inst = 32'h10408000;
      35633: inst = 32'hc404c9b;
      35634: inst = 32'h8220000;
      35635: inst = 32'h10408000;
      35636: inst = 32'hc404c9c;
      35637: inst = 32'h8220000;
      35638: inst = 32'h10408000;
      35639: inst = 32'hc404ca3;
      35640: inst = 32'h8220000;
      35641: inst = 32'h10408000;
      35642: inst = 32'hc404ca4;
      35643: inst = 32'h8220000;
      35644: inst = 32'h10408000;
      35645: inst = 32'hc404ca5;
      35646: inst = 32'h8220000;
      35647: inst = 32'h10408000;
      35648: inst = 32'hc404ca6;
      35649: inst = 32'h8220000;
      35650: inst = 32'h10408000;
      35651: inst = 32'hc404ca7;
      35652: inst = 32'h8220000;
      35653: inst = 32'h10408000;
      35654: inst = 32'hc404ca8;
      35655: inst = 32'h8220000;
      35656: inst = 32'h10408000;
      35657: inst = 32'hc404ca9;
      35658: inst = 32'h8220000;
      35659: inst = 32'h10408000;
      35660: inst = 32'hc404caa;
      35661: inst = 32'h8220000;
      35662: inst = 32'h10408000;
      35663: inst = 32'hc404cab;
      35664: inst = 32'h8220000;
      35665: inst = 32'h10408000;
      35666: inst = 32'hc404cac;
      35667: inst = 32'h8220000;
      35668: inst = 32'h10408000;
      35669: inst = 32'hc404cad;
      35670: inst = 32'h8220000;
      35671: inst = 32'h10408000;
      35672: inst = 32'hc404cae;
      35673: inst = 32'h8220000;
      35674: inst = 32'h10408000;
      35675: inst = 32'hc404caf;
      35676: inst = 32'h8220000;
      35677: inst = 32'h10408000;
      35678: inst = 32'hc404cb0;
      35679: inst = 32'h8220000;
      35680: inst = 32'h10408000;
      35681: inst = 32'hc404cb1;
      35682: inst = 32'h8220000;
      35683: inst = 32'h10408000;
      35684: inst = 32'hc404cb2;
      35685: inst = 32'h8220000;
      35686: inst = 32'h10408000;
      35687: inst = 32'hc404cb3;
      35688: inst = 32'h8220000;
      35689: inst = 32'h10408000;
      35690: inst = 32'hc404cb4;
      35691: inst = 32'h8220000;
      35692: inst = 32'h10408000;
      35693: inst = 32'hc404cb5;
      35694: inst = 32'h8220000;
      35695: inst = 32'h10408000;
      35696: inst = 32'hc404cb6;
      35697: inst = 32'h8220000;
      35698: inst = 32'h10408000;
      35699: inst = 32'hc404cb7;
      35700: inst = 32'h8220000;
      35701: inst = 32'h10408000;
      35702: inst = 32'hc404cb8;
      35703: inst = 32'h8220000;
      35704: inst = 32'h10408000;
      35705: inst = 32'hc404cb9;
      35706: inst = 32'h8220000;
      35707: inst = 32'h10408000;
      35708: inst = 32'hc404cba;
      35709: inst = 32'h8220000;
      35710: inst = 32'h10408000;
      35711: inst = 32'hc404cbb;
      35712: inst = 32'h8220000;
      35713: inst = 32'h10408000;
      35714: inst = 32'hc404cbc;
      35715: inst = 32'h8220000;
      35716: inst = 32'h10408000;
      35717: inst = 32'hc404cbd;
      35718: inst = 32'h8220000;
      35719: inst = 32'h10408000;
      35720: inst = 32'hc404cbe;
      35721: inst = 32'h8220000;
      35722: inst = 32'h10408000;
      35723: inst = 32'hc404cbf;
      35724: inst = 32'h8220000;
      35725: inst = 32'h10408000;
      35726: inst = 32'hc404cc0;
      35727: inst = 32'h8220000;
      35728: inst = 32'h10408000;
      35729: inst = 32'hc404cc1;
      35730: inst = 32'h8220000;
      35731: inst = 32'h10408000;
      35732: inst = 32'hc404cc2;
      35733: inst = 32'h8220000;
      35734: inst = 32'h10408000;
      35735: inst = 32'hc404cc3;
      35736: inst = 32'h8220000;
      35737: inst = 32'h10408000;
      35738: inst = 32'hc404cc4;
      35739: inst = 32'h8220000;
      35740: inst = 32'h10408000;
      35741: inst = 32'hc404cc5;
      35742: inst = 32'h8220000;
      35743: inst = 32'h10408000;
      35744: inst = 32'hc404cc6;
      35745: inst = 32'h8220000;
      35746: inst = 32'h10408000;
      35747: inst = 32'hc404cc7;
      35748: inst = 32'h8220000;
      35749: inst = 32'h10408000;
      35750: inst = 32'hc404cc8;
      35751: inst = 32'h8220000;
      35752: inst = 32'h10408000;
      35753: inst = 32'hc404cc9;
      35754: inst = 32'h8220000;
      35755: inst = 32'h10408000;
      35756: inst = 32'hc404cca;
      35757: inst = 32'h8220000;
      35758: inst = 32'h10408000;
      35759: inst = 32'hc404ccb;
      35760: inst = 32'h8220000;
      35761: inst = 32'h10408000;
      35762: inst = 32'hc404ccc;
      35763: inst = 32'h8220000;
      35764: inst = 32'h10408000;
      35765: inst = 32'hc404ccd;
      35766: inst = 32'h8220000;
      35767: inst = 32'h10408000;
      35768: inst = 32'hc404cce;
      35769: inst = 32'h8220000;
      35770: inst = 32'h10408000;
      35771: inst = 32'hc404ccf;
      35772: inst = 32'h8220000;
      35773: inst = 32'h10408000;
      35774: inst = 32'hc404cd0;
      35775: inst = 32'h8220000;
      35776: inst = 32'h10408000;
      35777: inst = 32'hc404cd1;
      35778: inst = 32'h8220000;
      35779: inst = 32'h10408000;
      35780: inst = 32'hc404cd2;
      35781: inst = 32'h8220000;
      35782: inst = 32'h10408000;
      35783: inst = 32'hc404cd3;
      35784: inst = 32'h8220000;
      35785: inst = 32'h10408000;
      35786: inst = 32'hc404cd4;
      35787: inst = 32'h8220000;
      35788: inst = 32'h10408000;
      35789: inst = 32'hc404cd5;
      35790: inst = 32'h8220000;
      35791: inst = 32'h10408000;
      35792: inst = 32'hc404cd6;
      35793: inst = 32'h8220000;
      35794: inst = 32'h10408000;
      35795: inst = 32'hc404cd7;
      35796: inst = 32'h8220000;
      35797: inst = 32'h10408000;
      35798: inst = 32'hc404cd8;
      35799: inst = 32'h8220000;
      35800: inst = 32'h10408000;
      35801: inst = 32'hc404cd9;
      35802: inst = 32'h8220000;
      35803: inst = 32'h10408000;
      35804: inst = 32'hc404cda;
      35805: inst = 32'h8220000;
      35806: inst = 32'h10408000;
      35807: inst = 32'hc404cdb;
      35808: inst = 32'h8220000;
      35809: inst = 32'h10408000;
      35810: inst = 32'hc404cdc;
      35811: inst = 32'h8220000;
      35812: inst = 32'h10408000;
      35813: inst = 32'hc404cdd;
      35814: inst = 32'h8220000;
      35815: inst = 32'h10408000;
      35816: inst = 32'hc404cde;
      35817: inst = 32'h8220000;
      35818: inst = 32'h10408000;
      35819: inst = 32'hc404cdf;
      35820: inst = 32'h8220000;
      35821: inst = 32'h10408000;
      35822: inst = 32'hc404ce0;
      35823: inst = 32'h8220000;
      35824: inst = 32'h10408000;
      35825: inst = 32'hc404ce1;
      35826: inst = 32'h8220000;
      35827: inst = 32'h10408000;
      35828: inst = 32'hc404ce2;
      35829: inst = 32'h8220000;
      35830: inst = 32'h10408000;
      35831: inst = 32'hc404ce3;
      35832: inst = 32'h8220000;
      35833: inst = 32'h10408000;
      35834: inst = 32'hc404ce4;
      35835: inst = 32'h8220000;
      35836: inst = 32'h10408000;
      35837: inst = 32'hc404ce5;
      35838: inst = 32'h8220000;
      35839: inst = 32'h10408000;
      35840: inst = 32'hc404ce6;
      35841: inst = 32'h8220000;
      35842: inst = 32'h10408000;
      35843: inst = 32'hc404ce7;
      35844: inst = 32'h8220000;
      35845: inst = 32'h10408000;
      35846: inst = 32'hc404ce8;
      35847: inst = 32'h8220000;
      35848: inst = 32'h10408000;
      35849: inst = 32'hc404ce9;
      35850: inst = 32'h8220000;
      35851: inst = 32'h10408000;
      35852: inst = 32'hc404cea;
      35853: inst = 32'h8220000;
      35854: inst = 32'h10408000;
      35855: inst = 32'hc404ceb;
      35856: inst = 32'h8220000;
      35857: inst = 32'h10408000;
      35858: inst = 32'hc404cec;
      35859: inst = 32'h8220000;
      35860: inst = 32'h10408000;
      35861: inst = 32'hc404ced;
      35862: inst = 32'h8220000;
      35863: inst = 32'h10408000;
      35864: inst = 32'hc404cee;
      35865: inst = 32'h8220000;
      35866: inst = 32'h10408000;
      35867: inst = 32'hc404cef;
      35868: inst = 32'h8220000;
      35869: inst = 32'h10408000;
      35870: inst = 32'hc404cf0;
      35871: inst = 32'h8220000;
      35872: inst = 32'h10408000;
      35873: inst = 32'hc404cf1;
      35874: inst = 32'h8220000;
      35875: inst = 32'h10408000;
      35876: inst = 32'hc404cf2;
      35877: inst = 32'h8220000;
      35878: inst = 32'h10408000;
      35879: inst = 32'hc404cf3;
      35880: inst = 32'h8220000;
      35881: inst = 32'h10408000;
      35882: inst = 32'hc404cf4;
      35883: inst = 32'h8220000;
      35884: inst = 32'h10408000;
      35885: inst = 32'hc404cf5;
      35886: inst = 32'h8220000;
      35887: inst = 32'h10408000;
      35888: inst = 32'hc404cf6;
      35889: inst = 32'h8220000;
      35890: inst = 32'h10408000;
      35891: inst = 32'hc404cf7;
      35892: inst = 32'h8220000;
      35893: inst = 32'h10408000;
      35894: inst = 32'hc404cf8;
      35895: inst = 32'h8220000;
      35896: inst = 32'h10408000;
      35897: inst = 32'hc404cf9;
      35898: inst = 32'h8220000;
      35899: inst = 32'h10408000;
      35900: inst = 32'hc404cfa;
      35901: inst = 32'h8220000;
      35902: inst = 32'h10408000;
      35903: inst = 32'hc404cfb;
      35904: inst = 32'h8220000;
      35905: inst = 32'h10408000;
      35906: inst = 32'hc404cfc;
      35907: inst = 32'h8220000;
      35908: inst = 32'h10408000;
      35909: inst = 32'hc404d03;
      35910: inst = 32'h8220000;
      35911: inst = 32'h10408000;
      35912: inst = 32'hc404d04;
      35913: inst = 32'h8220000;
      35914: inst = 32'h10408000;
      35915: inst = 32'hc404d05;
      35916: inst = 32'h8220000;
      35917: inst = 32'h10408000;
      35918: inst = 32'hc404d06;
      35919: inst = 32'h8220000;
      35920: inst = 32'h10408000;
      35921: inst = 32'hc404d07;
      35922: inst = 32'h8220000;
      35923: inst = 32'h10408000;
      35924: inst = 32'hc404d08;
      35925: inst = 32'h8220000;
      35926: inst = 32'h10408000;
      35927: inst = 32'hc404d09;
      35928: inst = 32'h8220000;
      35929: inst = 32'h10408000;
      35930: inst = 32'hc404d0a;
      35931: inst = 32'h8220000;
      35932: inst = 32'h10408000;
      35933: inst = 32'hc404d0b;
      35934: inst = 32'h8220000;
      35935: inst = 32'h10408000;
      35936: inst = 32'hc404d0c;
      35937: inst = 32'h8220000;
      35938: inst = 32'h10408000;
      35939: inst = 32'hc404d0d;
      35940: inst = 32'h8220000;
      35941: inst = 32'h10408000;
      35942: inst = 32'hc404d0e;
      35943: inst = 32'h8220000;
      35944: inst = 32'h10408000;
      35945: inst = 32'hc404d0f;
      35946: inst = 32'h8220000;
      35947: inst = 32'h10408000;
      35948: inst = 32'hc404d10;
      35949: inst = 32'h8220000;
      35950: inst = 32'h10408000;
      35951: inst = 32'hc404d11;
      35952: inst = 32'h8220000;
      35953: inst = 32'h10408000;
      35954: inst = 32'hc404d12;
      35955: inst = 32'h8220000;
      35956: inst = 32'h10408000;
      35957: inst = 32'hc404d13;
      35958: inst = 32'h8220000;
      35959: inst = 32'h10408000;
      35960: inst = 32'hc404d14;
      35961: inst = 32'h8220000;
      35962: inst = 32'h10408000;
      35963: inst = 32'hc404d15;
      35964: inst = 32'h8220000;
      35965: inst = 32'h10408000;
      35966: inst = 32'hc404d16;
      35967: inst = 32'h8220000;
      35968: inst = 32'h10408000;
      35969: inst = 32'hc404d17;
      35970: inst = 32'h8220000;
      35971: inst = 32'h10408000;
      35972: inst = 32'hc404d18;
      35973: inst = 32'h8220000;
      35974: inst = 32'h10408000;
      35975: inst = 32'hc404d19;
      35976: inst = 32'h8220000;
      35977: inst = 32'h10408000;
      35978: inst = 32'hc404d1a;
      35979: inst = 32'h8220000;
      35980: inst = 32'h10408000;
      35981: inst = 32'hc404d1b;
      35982: inst = 32'h8220000;
      35983: inst = 32'h10408000;
      35984: inst = 32'hc404d1c;
      35985: inst = 32'h8220000;
      35986: inst = 32'h10408000;
      35987: inst = 32'hc404d1d;
      35988: inst = 32'h8220000;
      35989: inst = 32'h10408000;
      35990: inst = 32'hc404d1e;
      35991: inst = 32'h8220000;
      35992: inst = 32'h10408000;
      35993: inst = 32'hc404d1f;
      35994: inst = 32'h8220000;
      35995: inst = 32'h10408000;
      35996: inst = 32'hc404d20;
      35997: inst = 32'h8220000;
      35998: inst = 32'h10408000;
      35999: inst = 32'hc404d21;
      36000: inst = 32'h8220000;
      36001: inst = 32'h10408000;
      36002: inst = 32'hc404d22;
      36003: inst = 32'h8220000;
      36004: inst = 32'h10408000;
      36005: inst = 32'hc404d23;
      36006: inst = 32'h8220000;
      36007: inst = 32'h10408000;
      36008: inst = 32'hc404d24;
      36009: inst = 32'h8220000;
      36010: inst = 32'h10408000;
      36011: inst = 32'hc404d3b;
      36012: inst = 32'h8220000;
      36013: inst = 32'h10408000;
      36014: inst = 32'hc404d3c;
      36015: inst = 32'h8220000;
      36016: inst = 32'h10408000;
      36017: inst = 32'hc404d3d;
      36018: inst = 32'h8220000;
      36019: inst = 32'h10408000;
      36020: inst = 32'hc404d3e;
      36021: inst = 32'h8220000;
      36022: inst = 32'h10408000;
      36023: inst = 32'hc404d3f;
      36024: inst = 32'h8220000;
      36025: inst = 32'h10408000;
      36026: inst = 32'hc404d40;
      36027: inst = 32'h8220000;
      36028: inst = 32'h10408000;
      36029: inst = 32'hc404d41;
      36030: inst = 32'h8220000;
      36031: inst = 32'h10408000;
      36032: inst = 32'hc404d42;
      36033: inst = 32'h8220000;
      36034: inst = 32'h10408000;
      36035: inst = 32'hc404d43;
      36036: inst = 32'h8220000;
      36037: inst = 32'h10408000;
      36038: inst = 32'hc404d44;
      36039: inst = 32'h8220000;
      36040: inst = 32'h10408000;
      36041: inst = 32'hc404d45;
      36042: inst = 32'h8220000;
      36043: inst = 32'h10408000;
      36044: inst = 32'hc404d46;
      36045: inst = 32'h8220000;
      36046: inst = 32'h10408000;
      36047: inst = 32'hc404d47;
      36048: inst = 32'h8220000;
      36049: inst = 32'h10408000;
      36050: inst = 32'hc404d48;
      36051: inst = 32'h8220000;
      36052: inst = 32'h10408000;
      36053: inst = 32'hc404d49;
      36054: inst = 32'h8220000;
      36055: inst = 32'h10408000;
      36056: inst = 32'hc404d4a;
      36057: inst = 32'h8220000;
      36058: inst = 32'h10408000;
      36059: inst = 32'hc404d4b;
      36060: inst = 32'h8220000;
      36061: inst = 32'h10408000;
      36062: inst = 32'hc404d4c;
      36063: inst = 32'h8220000;
      36064: inst = 32'h10408000;
      36065: inst = 32'hc404d4d;
      36066: inst = 32'h8220000;
      36067: inst = 32'h10408000;
      36068: inst = 32'hc404d4e;
      36069: inst = 32'h8220000;
      36070: inst = 32'h10408000;
      36071: inst = 32'hc404d4f;
      36072: inst = 32'h8220000;
      36073: inst = 32'h10408000;
      36074: inst = 32'hc404d50;
      36075: inst = 32'h8220000;
      36076: inst = 32'h10408000;
      36077: inst = 32'hc404d51;
      36078: inst = 32'h8220000;
      36079: inst = 32'h10408000;
      36080: inst = 32'hc404d52;
      36081: inst = 32'h8220000;
      36082: inst = 32'h10408000;
      36083: inst = 32'hc404d53;
      36084: inst = 32'h8220000;
      36085: inst = 32'h10408000;
      36086: inst = 32'hc404d54;
      36087: inst = 32'h8220000;
      36088: inst = 32'h10408000;
      36089: inst = 32'hc404d55;
      36090: inst = 32'h8220000;
      36091: inst = 32'h10408000;
      36092: inst = 32'hc404d56;
      36093: inst = 32'h8220000;
      36094: inst = 32'h10408000;
      36095: inst = 32'hc404d57;
      36096: inst = 32'h8220000;
      36097: inst = 32'h10408000;
      36098: inst = 32'hc404d58;
      36099: inst = 32'h8220000;
      36100: inst = 32'h10408000;
      36101: inst = 32'hc404d59;
      36102: inst = 32'h8220000;
      36103: inst = 32'h10408000;
      36104: inst = 32'hc404d5a;
      36105: inst = 32'h8220000;
      36106: inst = 32'h10408000;
      36107: inst = 32'hc404d5b;
      36108: inst = 32'h8220000;
      36109: inst = 32'h10408000;
      36110: inst = 32'hc404d5c;
      36111: inst = 32'h8220000;
      36112: inst = 32'h10408000;
      36113: inst = 32'hc404d63;
      36114: inst = 32'h8220000;
      36115: inst = 32'h10408000;
      36116: inst = 32'hc404d64;
      36117: inst = 32'h8220000;
      36118: inst = 32'h10408000;
      36119: inst = 32'hc404d65;
      36120: inst = 32'h8220000;
      36121: inst = 32'h10408000;
      36122: inst = 32'hc404d66;
      36123: inst = 32'h8220000;
      36124: inst = 32'h10408000;
      36125: inst = 32'hc404d67;
      36126: inst = 32'h8220000;
      36127: inst = 32'h10408000;
      36128: inst = 32'hc404d68;
      36129: inst = 32'h8220000;
      36130: inst = 32'h10408000;
      36131: inst = 32'hc404d69;
      36132: inst = 32'h8220000;
      36133: inst = 32'h10408000;
      36134: inst = 32'hc404d6a;
      36135: inst = 32'h8220000;
      36136: inst = 32'h10408000;
      36137: inst = 32'hc404d6b;
      36138: inst = 32'h8220000;
      36139: inst = 32'h10408000;
      36140: inst = 32'hc404d6c;
      36141: inst = 32'h8220000;
      36142: inst = 32'h10408000;
      36143: inst = 32'hc404d6d;
      36144: inst = 32'h8220000;
      36145: inst = 32'h10408000;
      36146: inst = 32'hc404d6e;
      36147: inst = 32'h8220000;
      36148: inst = 32'h10408000;
      36149: inst = 32'hc404d6f;
      36150: inst = 32'h8220000;
      36151: inst = 32'h10408000;
      36152: inst = 32'hc404d70;
      36153: inst = 32'h8220000;
      36154: inst = 32'h10408000;
      36155: inst = 32'hc404d71;
      36156: inst = 32'h8220000;
      36157: inst = 32'h10408000;
      36158: inst = 32'hc404d72;
      36159: inst = 32'h8220000;
      36160: inst = 32'h10408000;
      36161: inst = 32'hc404d73;
      36162: inst = 32'h8220000;
      36163: inst = 32'h10408000;
      36164: inst = 32'hc404d74;
      36165: inst = 32'h8220000;
      36166: inst = 32'h10408000;
      36167: inst = 32'hc404d75;
      36168: inst = 32'h8220000;
      36169: inst = 32'h10408000;
      36170: inst = 32'hc404d76;
      36171: inst = 32'h8220000;
      36172: inst = 32'h10408000;
      36173: inst = 32'hc404d77;
      36174: inst = 32'h8220000;
      36175: inst = 32'h10408000;
      36176: inst = 32'hc404d78;
      36177: inst = 32'h8220000;
      36178: inst = 32'h10408000;
      36179: inst = 32'hc404d79;
      36180: inst = 32'h8220000;
      36181: inst = 32'h10408000;
      36182: inst = 32'hc404d7a;
      36183: inst = 32'h8220000;
      36184: inst = 32'h10408000;
      36185: inst = 32'hc404d7b;
      36186: inst = 32'h8220000;
      36187: inst = 32'h10408000;
      36188: inst = 32'hc404d7c;
      36189: inst = 32'h8220000;
      36190: inst = 32'h10408000;
      36191: inst = 32'hc404d7d;
      36192: inst = 32'h8220000;
      36193: inst = 32'h10408000;
      36194: inst = 32'hc404d7e;
      36195: inst = 32'h8220000;
      36196: inst = 32'h10408000;
      36197: inst = 32'hc404d7f;
      36198: inst = 32'h8220000;
      36199: inst = 32'h10408000;
      36200: inst = 32'hc404d80;
      36201: inst = 32'h8220000;
      36202: inst = 32'h10408000;
      36203: inst = 32'hc404d81;
      36204: inst = 32'h8220000;
      36205: inst = 32'h10408000;
      36206: inst = 32'hc404d82;
      36207: inst = 32'h8220000;
      36208: inst = 32'h10408000;
      36209: inst = 32'hc404d83;
      36210: inst = 32'h8220000;
      36211: inst = 32'h10408000;
      36212: inst = 32'hc404d84;
      36213: inst = 32'h8220000;
      36214: inst = 32'h10408000;
      36215: inst = 32'hc404d9b;
      36216: inst = 32'h8220000;
      36217: inst = 32'h10408000;
      36218: inst = 32'hc404d9c;
      36219: inst = 32'h8220000;
      36220: inst = 32'h10408000;
      36221: inst = 32'hc404d9d;
      36222: inst = 32'h8220000;
      36223: inst = 32'h10408000;
      36224: inst = 32'hc404d9e;
      36225: inst = 32'h8220000;
      36226: inst = 32'h10408000;
      36227: inst = 32'hc404d9f;
      36228: inst = 32'h8220000;
      36229: inst = 32'h10408000;
      36230: inst = 32'hc404da0;
      36231: inst = 32'h8220000;
      36232: inst = 32'h10408000;
      36233: inst = 32'hc404da1;
      36234: inst = 32'h8220000;
      36235: inst = 32'h10408000;
      36236: inst = 32'hc404da2;
      36237: inst = 32'h8220000;
      36238: inst = 32'h10408000;
      36239: inst = 32'hc404da3;
      36240: inst = 32'h8220000;
      36241: inst = 32'h10408000;
      36242: inst = 32'hc404da4;
      36243: inst = 32'h8220000;
      36244: inst = 32'h10408000;
      36245: inst = 32'hc404da5;
      36246: inst = 32'h8220000;
      36247: inst = 32'h10408000;
      36248: inst = 32'hc404da6;
      36249: inst = 32'h8220000;
      36250: inst = 32'h10408000;
      36251: inst = 32'hc404da7;
      36252: inst = 32'h8220000;
      36253: inst = 32'h10408000;
      36254: inst = 32'hc404da8;
      36255: inst = 32'h8220000;
      36256: inst = 32'h10408000;
      36257: inst = 32'hc404da9;
      36258: inst = 32'h8220000;
      36259: inst = 32'h10408000;
      36260: inst = 32'hc404daa;
      36261: inst = 32'h8220000;
      36262: inst = 32'h10408000;
      36263: inst = 32'hc404dab;
      36264: inst = 32'h8220000;
      36265: inst = 32'h10408000;
      36266: inst = 32'hc404dac;
      36267: inst = 32'h8220000;
      36268: inst = 32'h10408000;
      36269: inst = 32'hc404dad;
      36270: inst = 32'h8220000;
      36271: inst = 32'h10408000;
      36272: inst = 32'hc404dae;
      36273: inst = 32'h8220000;
      36274: inst = 32'h10408000;
      36275: inst = 32'hc404daf;
      36276: inst = 32'h8220000;
      36277: inst = 32'h10408000;
      36278: inst = 32'hc404db0;
      36279: inst = 32'h8220000;
      36280: inst = 32'h10408000;
      36281: inst = 32'hc404db1;
      36282: inst = 32'h8220000;
      36283: inst = 32'h10408000;
      36284: inst = 32'hc404db2;
      36285: inst = 32'h8220000;
      36286: inst = 32'h10408000;
      36287: inst = 32'hc404db3;
      36288: inst = 32'h8220000;
      36289: inst = 32'h10408000;
      36290: inst = 32'hc404db4;
      36291: inst = 32'h8220000;
      36292: inst = 32'h10408000;
      36293: inst = 32'hc404db5;
      36294: inst = 32'h8220000;
      36295: inst = 32'h10408000;
      36296: inst = 32'hc404db6;
      36297: inst = 32'h8220000;
      36298: inst = 32'h10408000;
      36299: inst = 32'hc404db7;
      36300: inst = 32'h8220000;
      36301: inst = 32'h10408000;
      36302: inst = 32'hc404db8;
      36303: inst = 32'h8220000;
      36304: inst = 32'h10408000;
      36305: inst = 32'hc404db9;
      36306: inst = 32'h8220000;
      36307: inst = 32'h10408000;
      36308: inst = 32'hc404dba;
      36309: inst = 32'h8220000;
      36310: inst = 32'h10408000;
      36311: inst = 32'hc404dbb;
      36312: inst = 32'h8220000;
      36313: inst = 32'h10408000;
      36314: inst = 32'hc404dbc;
      36315: inst = 32'h8220000;
      36316: inst = 32'h10408000;
      36317: inst = 32'hc404dc3;
      36318: inst = 32'h8220000;
      36319: inst = 32'h10408000;
      36320: inst = 32'hc404dc4;
      36321: inst = 32'h8220000;
      36322: inst = 32'h10408000;
      36323: inst = 32'hc404dc5;
      36324: inst = 32'h8220000;
      36325: inst = 32'h10408000;
      36326: inst = 32'hc404dc6;
      36327: inst = 32'h8220000;
      36328: inst = 32'h10408000;
      36329: inst = 32'hc404dc7;
      36330: inst = 32'h8220000;
      36331: inst = 32'h10408000;
      36332: inst = 32'hc404dc8;
      36333: inst = 32'h8220000;
      36334: inst = 32'h10408000;
      36335: inst = 32'hc404dc9;
      36336: inst = 32'h8220000;
      36337: inst = 32'h10408000;
      36338: inst = 32'hc404dca;
      36339: inst = 32'h8220000;
      36340: inst = 32'h10408000;
      36341: inst = 32'hc404dcb;
      36342: inst = 32'h8220000;
      36343: inst = 32'h10408000;
      36344: inst = 32'hc404dcc;
      36345: inst = 32'h8220000;
      36346: inst = 32'h10408000;
      36347: inst = 32'hc404dcd;
      36348: inst = 32'h8220000;
      36349: inst = 32'h10408000;
      36350: inst = 32'hc404dce;
      36351: inst = 32'h8220000;
      36352: inst = 32'h10408000;
      36353: inst = 32'hc404dcf;
      36354: inst = 32'h8220000;
      36355: inst = 32'h10408000;
      36356: inst = 32'hc404dd0;
      36357: inst = 32'h8220000;
      36358: inst = 32'h10408000;
      36359: inst = 32'hc404dd1;
      36360: inst = 32'h8220000;
      36361: inst = 32'h10408000;
      36362: inst = 32'hc404dd2;
      36363: inst = 32'h8220000;
      36364: inst = 32'h10408000;
      36365: inst = 32'hc404dd3;
      36366: inst = 32'h8220000;
      36367: inst = 32'h10408000;
      36368: inst = 32'hc404dd4;
      36369: inst = 32'h8220000;
      36370: inst = 32'h10408000;
      36371: inst = 32'hc404dd5;
      36372: inst = 32'h8220000;
      36373: inst = 32'h10408000;
      36374: inst = 32'hc404dd6;
      36375: inst = 32'h8220000;
      36376: inst = 32'h10408000;
      36377: inst = 32'hc404dd7;
      36378: inst = 32'h8220000;
      36379: inst = 32'h10408000;
      36380: inst = 32'hc404dd8;
      36381: inst = 32'h8220000;
      36382: inst = 32'h10408000;
      36383: inst = 32'hc404dd9;
      36384: inst = 32'h8220000;
      36385: inst = 32'h10408000;
      36386: inst = 32'hc404dda;
      36387: inst = 32'h8220000;
      36388: inst = 32'h10408000;
      36389: inst = 32'hc404ddb;
      36390: inst = 32'h8220000;
      36391: inst = 32'h10408000;
      36392: inst = 32'hc404ddc;
      36393: inst = 32'h8220000;
      36394: inst = 32'h10408000;
      36395: inst = 32'hc404ddd;
      36396: inst = 32'h8220000;
      36397: inst = 32'h10408000;
      36398: inst = 32'hc404dde;
      36399: inst = 32'h8220000;
      36400: inst = 32'h10408000;
      36401: inst = 32'hc404ddf;
      36402: inst = 32'h8220000;
      36403: inst = 32'h10408000;
      36404: inst = 32'hc404de0;
      36405: inst = 32'h8220000;
      36406: inst = 32'h10408000;
      36407: inst = 32'hc404de1;
      36408: inst = 32'h8220000;
      36409: inst = 32'h10408000;
      36410: inst = 32'hc404de2;
      36411: inst = 32'h8220000;
      36412: inst = 32'h10408000;
      36413: inst = 32'hc404de3;
      36414: inst = 32'h8220000;
      36415: inst = 32'h10408000;
      36416: inst = 32'hc404de4;
      36417: inst = 32'h8220000;
      36418: inst = 32'h10408000;
      36419: inst = 32'hc404dfb;
      36420: inst = 32'h8220000;
      36421: inst = 32'h10408000;
      36422: inst = 32'hc404dfc;
      36423: inst = 32'h8220000;
      36424: inst = 32'h10408000;
      36425: inst = 32'hc404dfd;
      36426: inst = 32'h8220000;
      36427: inst = 32'h10408000;
      36428: inst = 32'hc404dfe;
      36429: inst = 32'h8220000;
      36430: inst = 32'h10408000;
      36431: inst = 32'hc404dff;
      36432: inst = 32'h8220000;
      36433: inst = 32'h10408000;
      36434: inst = 32'hc404e00;
      36435: inst = 32'h8220000;
      36436: inst = 32'h10408000;
      36437: inst = 32'hc404e01;
      36438: inst = 32'h8220000;
      36439: inst = 32'h10408000;
      36440: inst = 32'hc404e02;
      36441: inst = 32'h8220000;
      36442: inst = 32'h10408000;
      36443: inst = 32'hc404e03;
      36444: inst = 32'h8220000;
      36445: inst = 32'h10408000;
      36446: inst = 32'hc404e04;
      36447: inst = 32'h8220000;
      36448: inst = 32'h10408000;
      36449: inst = 32'hc404e05;
      36450: inst = 32'h8220000;
      36451: inst = 32'h10408000;
      36452: inst = 32'hc404e06;
      36453: inst = 32'h8220000;
      36454: inst = 32'h10408000;
      36455: inst = 32'hc404e07;
      36456: inst = 32'h8220000;
      36457: inst = 32'h10408000;
      36458: inst = 32'hc404e08;
      36459: inst = 32'h8220000;
      36460: inst = 32'h10408000;
      36461: inst = 32'hc404e09;
      36462: inst = 32'h8220000;
      36463: inst = 32'h10408000;
      36464: inst = 32'hc404e0a;
      36465: inst = 32'h8220000;
      36466: inst = 32'h10408000;
      36467: inst = 32'hc404e0b;
      36468: inst = 32'h8220000;
      36469: inst = 32'h10408000;
      36470: inst = 32'hc404e0c;
      36471: inst = 32'h8220000;
      36472: inst = 32'h10408000;
      36473: inst = 32'hc404e0d;
      36474: inst = 32'h8220000;
      36475: inst = 32'h10408000;
      36476: inst = 32'hc404e0e;
      36477: inst = 32'h8220000;
      36478: inst = 32'h10408000;
      36479: inst = 32'hc404e0f;
      36480: inst = 32'h8220000;
      36481: inst = 32'h10408000;
      36482: inst = 32'hc404e10;
      36483: inst = 32'h8220000;
      36484: inst = 32'h10408000;
      36485: inst = 32'hc404e11;
      36486: inst = 32'h8220000;
      36487: inst = 32'h10408000;
      36488: inst = 32'hc404e12;
      36489: inst = 32'h8220000;
      36490: inst = 32'h10408000;
      36491: inst = 32'hc404e13;
      36492: inst = 32'h8220000;
      36493: inst = 32'h10408000;
      36494: inst = 32'hc404e14;
      36495: inst = 32'h8220000;
      36496: inst = 32'h10408000;
      36497: inst = 32'hc404e15;
      36498: inst = 32'h8220000;
      36499: inst = 32'h10408000;
      36500: inst = 32'hc404e16;
      36501: inst = 32'h8220000;
      36502: inst = 32'h10408000;
      36503: inst = 32'hc404e17;
      36504: inst = 32'h8220000;
      36505: inst = 32'h10408000;
      36506: inst = 32'hc404e18;
      36507: inst = 32'h8220000;
      36508: inst = 32'h10408000;
      36509: inst = 32'hc404e19;
      36510: inst = 32'h8220000;
      36511: inst = 32'h10408000;
      36512: inst = 32'hc404e1a;
      36513: inst = 32'h8220000;
      36514: inst = 32'h10408000;
      36515: inst = 32'hc404e1b;
      36516: inst = 32'h8220000;
      36517: inst = 32'h10408000;
      36518: inst = 32'hc404e1c;
      36519: inst = 32'h8220000;
      36520: inst = 32'h10408000;
      36521: inst = 32'hc404e23;
      36522: inst = 32'h8220000;
      36523: inst = 32'h10408000;
      36524: inst = 32'hc404e24;
      36525: inst = 32'h8220000;
      36526: inst = 32'h10408000;
      36527: inst = 32'hc404e25;
      36528: inst = 32'h8220000;
      36529: inst = 32'h10408000;
      36530: inst = 32'hc404e26;
      36531: inst = 32'h8220000;
      36532: inst = 32'h10408000;
      36533: inst = 32'hc404e27;
      36534: inst = 32'h8220000;
      36535: inst = 32'h10408000;
      36536: inst = 32'hc404e28;
      36537: inst = 32'h8220000;
      36538: inst = 32'h10408000;
      36539: inst = 32'hc404e29;
      36540: inst = 32'h8220000;
      36541: inst = 32'h10408000;
      36542: inst = 32'hc404e2a;
      36543: inst = 32'h8220000;
      36544: inst = 32'h10408000;
      36545: inst = 32'hc404e2b;
      36546: inst = 32'h8220000;
      36547: inst = 32'h10408000;
      36548: inst = 32'hc404e2c;
      36549: inst = 32'h8220000;
      36550: inst = 32'h10408000;
      36551: inst = 32'hc404e2d;
      36552: inst = 32'h8220000;
      36553: inst = 32'h10408000;
      36554: inst = 32'hc404e2e;
      36555: inst = 32'h8220000;
      36556: inst = 32'h10408000;
      36557: inst = 32'hc404e2f;
      36558: inst = 32'h8220000;
      36559: inst = 32'h10408000;
      36560: inst = 32'hc404e30;
      36561: inst = 32'h8220000;
      36562: inst = 32'h10408000;
      36563: inst = 32'hc404e31;
      36564: inst = 32'h8220000;
      36565: inst = 32'h10408000;
      36566: inst = 32'hc404e32;
      36567: inst = 32'h8220000;
      36568: inst = 32'h10408000;
      36569: inst = 32'hc404e33;
      36570: inst = 32'h8220000;
      36571: inst = 32'h10408000;
      36572: inst = 32'hc404e34;
      36573: inst = 32'h8220000;
      36574: inst = 32'h10408000;
      36575: inst = 32'hc404e35;
      36576: inst = 32'h8220000;
      36577: inst = 32'h10408000;
      36578: inst = 32'hc404e36;
      36579: inst = 32'h8220000;
      36580: inst = 32'h10408000;
      36581: inst = 32'hc404e37;
      36582: inst = 32'h8220000;
      36583: inst = 32'h10408000;
      36584: inst = 32'hc404e38;
      36585: inst = 32'h8220000;
      36586: inst = 32'h10408000;
      36587: inst = 32'hc404e39;
      36588: inst = 32'h8220000;
      36589: inst = 32'h10408000;
      36590: inst = 32'hc404e3a;
      36591: inst = 32'h8220000;
      36592: inst = 32'h10408000;
      36593: inst = 32'hc404e3b;
      36594: inst = 32'h8220000;
      36595: inst = 32'h10408000;
      36596: inst = 32'hc404e3c;
      36597: inst = 32'h8220000;
      36598: inst = 32'h10408000;
      36599: inst = 32'hc404e3d;
      36600: inst = 32'h8220000;
      36601: inst = 32'h10408000;
      36602: inst = 32'hc404e3e;
      36603: inst = 32'h8220000;
      36604: inst = 32'h10408000;
      36605: inst = 32'hc404e3f;
      36606: inst = 32'h8220000;
      36607: inst = 32'h10408000;
      36608: inst = 32'hc404e40;
      36609: inst = 32'h8220000;
      36610: inst = 32'h10408000;
      36611: inst = 32'hc404e41;
      36612: inst = 32'h8220000;
      36613: inst = 32'h10408000;
      36614: inst = 32'hc404e42;
      36615: inst = 32'h8220000;
      36616: inst = 32'h10408000;
      36617: inst = 32'hc404e43;
      36618: inst = 32'h8220000;
      36619: inst = 32'h10408000;
      36620: inst = 32'hc404e44;
      36621: inst = 32'h8220000;
      36622: inst = 32'h10408000;
      36623: inst = 32'hc404e45;
      36624: inst = 32'h8220000;
      36625: inst = 32'h10408000;
      36626: inst = 32'hc404e46;
      36627: inst = 32'h8220000;
      36628: inst = 32'h10408000;
      36629: inst = 32'hc404e47;
      36630: inst = 32'h8220000;
      36631: inst = 32'h10408000;
      36632: inst = 32'hc404e48;
      36633: inst = 32'h8220000;
      36634: inst = 32'h10408000;
      36635: inst = 32'hc404e49;
      36636: inst = 32'h8220000;
      36637: inst = 32'h10408000;
      36638: inst = 32'hc404e4a;
      36639: inst = 32'h8220000;
      36640: inst = 32'h10408000;
      36641: inst = 32'hc404e4b;
      36642: inst = 32'h8220000;
      36643: inst = 32'h10408000;
      36644: inst = 32'hc404e4c;
      36645: inst = 32'h8220000;
      36646: inst = 32'h10408000;
      36647: inst = 32'hc404e4d;
      36648: inst = 32'h8220000;
      36649: inst = 32'h10408000;
      36650: inst = 32'hc404e4e;
      36651: inst = 32'h8220000;
      36652: inst = 32'h10408000;
      36653: inst = 32'hc404e4f;
      36654: inst = 32'h8220000;
      36655: inst = 32'h10408000;
      36656: inst = 32'hc404e50;
      36657: inst = 32'h8220000;
      36658: inst = 32'h10408000;
      36659: inst = 32'hc404e51;
      36660: inst = 32'h8220000;
      36661: inst = 32'h10408000;
      36662: inst = 32'hc404e52;
      36663: inst = 32'h8220000;
      36664: inst = 32'h10408000;
      36665: inst = 32'hc404e53;
      36666: inst = 32'h8220000;
      36667: inst = 32'h10408000;
      36668: inst = 32'hc404e54;
      36669: inst = 32'h8220000;
      36670: inst = 32'h10408000;
      36671: inst = 32'hc404e55;
      36672: inst = 32'h8220000;
      36673: inst = 32'h10408000;
      36674: inst = 32'hc404e56;
      36675: inst = 32'h8220000;
      36676: inst = 32'h10408000;
      36677: inst = 32'hc404e57;
      36678: inst = 32'h8220000;
      36679: inst = 32'h10408000;
      36680: inst = 32'hc404e5b;
      36681: inst = 32'h8220000;
      36682: inst = 32'h10408000;
      36683: inst = 32'hc404e5c;
      36684: inst = 32'h8220000;
      36685: inst = 32'h10408000;
      36686: inst = 32'hc404e5d;
      36687: inst = 32'h8220000;
      36688: inst = 32'h10408000;
      36689: inst = 32'hc404e5e;
      36690: inst = 32'h8220000;
      36691: inst = 32'h10408000;
      36692: inst = 32'hc404e5f;
      36693: inst = 32'h8220000;
      36694: inst = 32'h10408000;
      36695: inst = 32'hc404e60;
      36696: inst = 32'h8220000;
      36697: inst = 32'h10408000;
      36698: inst = 32'hc404e61;
      36699: inst = 32'h8220000;
      36700: inst = 32'h10408000;
      36701: inst = 32'hc404e62;
      36702: inst = 32'h8220000;
      36703: inst = 32'h10408000;
      36704: inst = 32'hc404e63;
      36705: inst = 32'h8220000;
      36706: inst = 32'h10408000;
      36707: inst = 32'hc404e64;
      36708: inst = 32'h8220000;
      36709: inst = 32'h10408000;
      36710: inst = 32'hc404e65;
      36711: inst = 32'h8220000;
      36712: inst = 32'h10408000;
      36713: inst = 32'hc404e66;
      36714: inst = 32'h8220000;
      36715: inst = 32'h10408000;
      36716: inst = 32'hc404e67;
      36717: inst = 32'h8220000;
      36718: inst = 32'h10408000;
      36719: inst = 32'hc404e68;
      36720: inst = 32'h8220000;
      36721: inst = 32'h10408000;
      36722: inst = 32'hc404e69;
      36723: inst = 32'h8220000;
      36724: inst = 32'h10408000;
      36725: inst = 32'hc404e6a;
      36726: inst = 32'h8220000;
      36727: inst = 32'h10408000;
      36728: inst = 32'hc404e6b;
      36729: inst = 32'h8220000;
      36730: inst = 32'h10408000;
      36731: inst = 32'hc404e6c;
      36732: inst = 32'h8220000;
      36733: inst = 32'h10408000;
      36734: inst = 32'hc404e6d;
      36735: inst = 32'h8220000;
      36736: inst = 32'h10408000;
      36737: inst = 32'hc404e6e;
      36738: inst = 32'h8220000;
      36739: inst = 32'h10408000;
      36740: inst = 32'hc404e6f;
      36741: inst = 32'h8220000;
      36742: inst = 32'h10408000;
      36743: inst = 32'hc404e70;
      36744: inst = 32'h8220000;
      36745: inst = 32'h10408000;
      36746: inst = 32'hc404e71;
      36747: inst = 32'h8220000;
      36748: inst = 32'h10408000;
      36749: inst = 32'hc404e72;
      36750: inst = 32'h8220000;
      36751: inst = 32'h10408000;
      36752: inst = 32'hc404e73;
      36753: inst = 32'h8220000;
      36754: inst = 32'h10408000;
      36755: inst = 32'hc404e74;
      36756: inst = 32'h8220000;
      36757: inst = 32'h10408000;
      36758: inst = 32'hc404e75;
      36759: inst = 32'h8220000;
      36760: inst = 32'h10408000;
      36761: inst = 32'hc404e76;
      36762: inst = 32'h8220000;
      36763: inst = 32'h10408000;
      36764: inst = 32'hc404e77;
      36765: inst = 32'h8220000;
      36766: inst = 32'h10408000;
      36767: inst = 32'hc404e78;
      36768: inst = 32'h8220000;
      36769: inst = 32'h10408000;
      36770: inst = 32'hc404e79;
      36771: inst = 32'h8220000;
      36772: inst = 32'h10408000;
      36773: inst = 32'hc404e7a;
      36774: inst = 32'h8220000;
      36775: inst = 32'h10408000;
      36776: inst = 32'hc404e7b;
      36777: inst = 32'h8220000;
      36778: inst = 32'h10408000;
      36779: inst = 32'hc404e7c;
      36780: inst = 32'h8220000;
      36781: inst = 32'h10408000;
      36782: inst = 32'hc404e83;
      36783: inst = 32'h8220000;
      36784: inst = 32'h10408000;
      36785: inst = 32'hc404e84;
      36786: inst = 32'h8220000;
      36787: inst = 32'h10408000;
      36788: inst = 32'hc404e85;
      36789: inst = 32'h8220000;
      36790: inst = 32'h10408000;
      36791: inst = 32'hc404e86;
      36792: inst = 32'h8220000;
      36793: inst = 32'h10408000;
      36794: inst = 32'hc404e87;
      36795: inst = 32'h8220000;
      36796: inst = 32'h10408000;
      36797: inst = 32'hc404e88;
      36798: inst = 32'h8220000;
      36799: inst = 32'h10408000;
      36800: inst = 32'hc404e89;
      36801: inst = 32'h8220000;
      36802: inst = 32'h10408000;
      36803: inst = 32'hc404e8a;
      36804: inst = 32'h8220000;
      36805: inst = 32'h10408000;
      36806: inst = 32'hc404e8b;
      36807: inst = 32'h8220000;
      36808: inst = 32'h10408000;
      36809: inst = 32'hc404e8c;
      36810: inst = 32'h8220000;
      36811: inst = 32'h10408000;
      36812: inst = 32'hc404e8d;
      36813: inst = 32'h8220000;
      36814: inst = 32'h10408000;
      36815: inst = 32'hc404e8e;
      36816: inst = 32'h8220000;
      36817: inst = 32'h10408000;
      36818: inst = 32'hc404e8f;
      36819: inst = 32'h8220000;
      36820: inst = 32'h10408000;
      36821: inst = 32'hc404e90;
      36822: inst = 32'h8220000;
      36823: inst = 32'h10408000;
      36824: inst = 32'hc404e91;
      36825: inst = 32'h8220000;
      36826: inst = 32'h10408000;
      36827: inst = 32'hc404e92;
      36828: inst = 32'h8220000;
      36829: inst = 32'h10408000;
      36830: inst = 32'hc404e93;
      36831: inst = 32'h8220000;
      36832: inst = 32'h10408000;
      36833: inst = 32'hc404e94;
      36834: inst = 32'h8220000;
      36835: inst = 32'h10408000;
      36836: inst = 32'hc404e95;
      36837: inst = 32'h8220000;
      36838: inst = 32'h10408000;
      36839: inst = 32'hc404e96;
      36840: inst = 32'h8220000;
      36841: inst = 32'h10408000;
      36842: inst = 32'hc404e97;
      36843: inst = 32'h8220000;
      36844: inst = 32'h10408000;
      36845: inst = 32'hc404e98;
      36846: inst = 32'h8220000;
      36847: inst = 32'h10408000;
      36848: inst = 32'hc404e99;
      36849: inst = 32'h8220000;
      36850: inst = 32'h10408000;
      36851: inst = 32'hc404e9a;
      36852: inst = 32'h8220000;
      36853: inst = 32'h10408000;
      36854: inst = 32'hc404e9b;
      36855: inst = 32'h8220000;
      36856: inst = 32'h10408000;
      36857: inst = 32'hc404e9c;
      36858: inst = 32'h8220000;
      36859: inst = 32'h10408000;
      36860: inst = 32'hc404e9d;
      36861: inst = 32'h8220000;
      36862: inst = 32'h10408000;
      36863: inst = 32'hc404e9e;
      36864: inst = 32'h8220000;
      36865: inst = 32'h10408000;
      36866: inst = 32'hc404e9f;
      36867: inst = 32'h8220000;
      36868: inst = 32'h10408000;
      36869: inst = 32'hc404ea0;
      36870: inst = 32'h8220000;
      36871: inst = 32'h10408000;
      36872: inst = 32'hc404ea1;
      36873: inst = 32'h8220000;
      36874: inst = 32'h10408000;
      36875: inst = 32'hc404ea2;
      36876: inst = 32'h8220000;
      36877: inst = 32'h10408000;
      36878: inst = 32'hc404ea3;
      36879: inst = 32'h8220000;
      36880: inst = 32'h10408000;
      36881: inst = 32'hc404ea4;
      36882: inst = 32'h8220000;
      36883: inst = 32'h10408000;
      36884: inst = 32'hc404ea5;
      36885: inst = 32'h8220000;
      36886: inst = 32'h10408000;
      36887: inst = 32'hc404ea6;
      36888: inst = 32'h8220000;
      36889: inst = 32'h10408000;
      36890: inst = 32'hc404ea7;
      36891: inst = 32'h8220000;
      36892: inst = 32'h10408000;
      36893: inst = 32'hc404ea8;
      36894: inst = 32'h8220000;
      36895: inst = 32'h10408000;
      36896: inst = 32'hc404ea9;
      36897: inst = 32'h8220000;
      36898: inst = 32'h10408000;
      36899: inst = 32'hc404eaa;
      36900: inst = 32'h8220000;
      36901: inst = 32'h10408000;
      36902: inst = 32'hc404eab;
      36903: inst = 32'h8220000;
      36904: inst = 32'h10408000;
      36905: inst = 32'hc404eac;
      36906: inst = 32'h8220000;
      36907: inst = 32'h10408000;
      36908: inst = 32'hc404ead;
      36909: inst = 32'h8220000;
      36910: inst = 32'h10408000;
      36911: inst = 32'hc404eae;
      36912: inst = 32'h8220000;
      36913: inst = 32'h10408000;
      36914: inst = 32'hc404eaf;
      36915: inst = 32'h8220000;
      36916: inst = 32'h10408000;
      36917: inst = 32'hc404eb0;
      36918: inst = 32'h8220000;
      36919: inst = 32'h10408000;
      36920: inst = 32'hc404eb1;
      36921: inst = 32'h8220000;
      36922: inst = 32'h10408000;
      36923: inst = 32'hc404eb2;
      36924: inst = 32'h8220000;
      36925: inst = 32'h10408000;
      36926: inst = 32'hc404eb3;
      36927: inst = 32'h8220000;
      36928: inst = 32'h10408000;
      36929: inst = 32'hc404eb4;
      36930: inst = 32'h8220000;
      36931: inst = 32'h10408000;
      36932: inst = 32'hc404eb5;
      36933: inst = 32'h8220000;
      36934: inst = 32'h10408000;
      36935: inst = 32'hc404eb6;
      36936: inst = 32'h8220000;
      36937: inst = 32'h10408000;
      36938: inst = 32'hc404eb7;
      36939: inst = 32'h8220000;
      36940: inst = 32'h10408000;
      36941: inst = 32'hc404ebb;
      36942: inst = 32'h8220000;
      36943: inst = 32'h10408000;
      36944: inst = 32'hc404ebc;
      36945: inst = 32'h8220000;
      36946: inst = 32'h10408000;
      36947: inst = 32'hc404ebd;
      36948: inst = 32'h8220000;
      36949: inst = 32'h10408000;
      36950: inst = 32'hc404ebe;
      36951: inst = 32'h8220000;
      36952: inst = 32'h10408000;
      36953: inst = 32'hc404ebf;
      36954: inst = 32'h8220000;
      36955: inst = 32'h10408000;
      36956: inst = 32'hc404ec0;
      36957: inst = 32'h8220000;
      36958: inst = 32'h10408000;
      36959: inst = 32'hc404ec1;
      36960: inst = 32'h8220000;
      36961: inst = 32'h10408000;
      36962: inst = 32'hc404ec2;
      36963: inst = 32'h8220000;
      36964: inst = 32'h10408000;
      36965: inst = 32'hc404ec3;
      36966: inst = 32'h8220000;
      36967: inst = 32'h10408000;
      36968: inst = 32'hc404ec4;
      36969: inst = 32'h8220000;
      36970: inst = 32'h10408000;
      36971: inst = 32'hc404ec5;
      36972: inst = 32'h8220000;
      36973: inst = 32'h10408000;
      36974: inst = 32'hc404ec6;
      36975: inst = 32'h8220000;
      36976: inst = 32'h10408000;
      36977: inst = 32'hc404ec7;
      36978: inst = 32'h8220000;
      36979: inst = 32'h10408000;
      36980: inst = 32'hc404ec8;
      36981: inst = 32'h8220000;
      36982: inst = 32'h10408000;
      36983: inst = 32'hc404ec9;
      36984: inst = 32'h8220000;
      36985: inst = 32'h10408000;
      36986: inst = 32'hc404eca;
      36987: inst = 32'h8220000;
      36988: inst = 32'h10408000;
      36989: inst = 32'hc404ecb;
      36990: inst = 32'h8220000;
      36991: inst = 32'h10408000;
      36992: inst = 32'hc404ecc;
      36993: inst = 32'h8220000;
      36994: inst = 32'h10408000;
      36995: inst = 32'hc404ecd;
      36996: inst = 32'h8220000;
      36997: inst = 32'h10408000;
      36998: inst = 32'hc404ece;
      36999: inst = 32'h8220000;
      37000: inst = 32'h10408000;
      37001: inst = 32'hc404ecf;
      37002: inst = 32'h8220000;
      37003: inst = 32'h10408000;
      37004: inst = 32'hc404ed0;
      37005: inst = 32'h8220000;
      37006: inst = 32'h10408000;
      37007: inst = 32'hc404ed1;
      37008: inst = 32'h8220000;
      37009: inst = 32'h10408000;
      37010: inst = 32'hc404ed2;
      37011: inst = 32'h8220000;
      37012: inst = 32'h10408000;
      37013: inst = 32'hc404ed3;
      37014: inst = 32'h8220000;
      37015: inst = 32'h10408000;
      37016: inst = 32'hc404ed4;
      37017: inst = 32'h8220000;
      37018: inst = 32'h10408000;
      37019: inst = 32'hc404ed5;
      37020: inst = 32'h8220000;
      37021: inst = 32'h10408000;
      37022: inst = 32'hc404ed6;
      37023: inst = 32'h8220000;
      37024: inst = 32'h10408000;
      37025: inst = 32'hc404ed7;
      37026: inst = 32'h8220000;
      37027: inst = 32'h10408000;
      37028: inst = 32'hc404ed8;
      37029: inst = 32'h8220000;
      37030: inst = 32'h10408000;
      37031: inst = 32'hc404ed9;
      37032: inst = 32'h8220000;
      37033: inst = 32'h10408000;
      37034: inst = 32'hc404eda;
      37035: inst = 32'h8220000;
      37036: inst = 32'h10408000;
      37037: inst = 32'hc404edb;
      37038: inst = 32'h8220000;
      37039: inst = 32'h10408000;
      37040: inst = 32'hc404edc;
      37041: inst = 32'h8220000;
      37042: inst = 32'h10408000;
      37043: inst = 32'hc404ee3;
      37044: inst = 32'h8220000;
      37045: inst = 32'h10408000;
      37046: inst = 32'hc404ee4;
      37047: inst = 32'h8220000;
      37048: inst = 32'h10408000;
      37049: inst = 32'hc404ee5;
      37050: inst = 32'h8220000;
      37051: inst = 32'h10408000;
      37052: inst = 32'hc404ee6;
      37053: inst = 32'h8220000;
      37054: inst = 32'h10408000;
      37055: inst = 32'hc404ee7;
      37056: inst = 32'h8220000;
      37057: inst = 32'h10408000;
      37058: inst = 32'hc404ee8;
      37059: inst = 32'h8220000;
      37060: inst = 32'h10408000;
      37061: inst = 32'hc404ee9;
      37062: inst = 32'h8220000;
      37063: inst = 32'h10408000;
      37064: inst = 32'hc404eea;
      37065: inst = 32'h8220000;
      37066: inst = 32'h10408000;
      37067: inst = 32'hc404eeb;
      37068: inst = 32'h8220000;
      37069: inst = 32'h10408000;
      37070: inst = 32'hc404eec;
      37071: inst = 32'h8220000;
      37072: inst = 32'h10408000;
      37073: inst = 32'hc404eed;
      37074: inst = 32'h8220000;
      37075: inst = 32'h10408000;
      37076: inst = 32'hc404eee;
      37077: inst = 32'h8220000;
      37078: inst = 32'h10408000;
      37079: inst = 32'hc404eef;
      37080: inst = 32'h8220000;
      37081: inst = 32'h10408000;
      37082: inst = 32'hc404ef0;
      37083: inst = 32'h8220000;
      37084: inst = 32'h10408000;
      37085: inst = 32'hc404ef1;
      37086: inst = 32'h8220000;
      37087: inst = 32'h10408000;
      37088: inst = 32'hc404ef2;
      37089: inst = 32'h8220000;
      37090: inst = 32'h10408000;
      37091: inst = 32'hc404ef3;
      37092: inst = 32'h8220000;
      37093: inst = 32'h10408000;
      37094: inst = 32'hc404ef4;
      37095: inst = 32'h8220000;
      37096: inst = 32'h10408000;
      37097: inst = 32'hc404ef5;
      37098: inst = 32'h8220000;
      37099: inst = 32'h10408000;
      37100: inst = 32'hc404ef6;
      37101: inst = 32'h8220000;
      37102: inst = 32'h10408000;
      37103: inst = 32'hc404ef7;
      37104: inst = 32'h8220000;
      37105: inst = 32'h10408000;
      37106: inst = 32'hc404ef8;
      37107: inst = 32'h8220000;
      37108: inst = 32'h10408000;
      37109: inst = 32'hc404ef9;
      37110: inst = 32'h8220000;
      37111: inst = 32'h10408000;
      37112: inst = 32'hc404efa;
      37113: inst = 32'h8220000;
      37114: inst = 32'h10408000;
      37115: inst = 32'hc404efb;
      37116: inst = 32'h8220000;
      37117: inst = 32'h10408000;
      37118: inst = 32'hc404efc;
      37119: inst = 32'h8220000;
      37120: inst = 32'h10408000;
      37121: inst = 32'hc404efd;
      37122: inst = 32'h8220000;
      37123: inst = 32'h10408000;
      37124: inst = 32'hc404efe;
      37125: inst = 32'h8220000;
      37126: inst = 32'h10408000;
      37127: inst = 32'hc404eff;
      37128: inst = 32'h8220000;
      37129: inst = 32'h10408000;
      37130: inst = 32'hc404f00;
      37131: inst = 32'h8220000;
      37132: inst = 32'h10408000;
      37133: inst = 32'hc404f01;
      37134: inst = 32'h8220000;
      37135: inst = 32'h10408000;
      37136: inst = 32'hc404f02;
      37137: inst = 32'h8220000;
      37138: inst = 32'h10408000;
      37139: inst = 32'hc404f03;
      37140: inst = 32'h8220000;
      37141: inst = 32'h10408000;
      37142: inst = 32'hc404f04;
      37143: inst = 32'h8220000;
      37144: inst = 32'h10408000;
      37145: inst = 32'hc404f05;
      37146: inst = 32'h8220000;
      37147: inst = 32'h10408000;
      37148: inst = 32'hc404f06;
      37149: inst = 32'h8220000;
      37150: inst = 32'h10408000;
      37151: inst = 32'hc404f07;
      37152: inst = 32'h8220000;
      37153: inst = 32'h10408000;
      37154: inst = 32'hc404f08;
      37155: inst = 32'h8220000;
      37156: inst = 32'h10408000;
      37157: inst = 32'hc404f09;
      37158: inst = 32'h8220000;
      37159: inst = 32'h10408000;
      37160: inst = 32'hc404f0a;
      37161: inst = 32'h8220000;
      37162: inst = 32'h10408000;
      37163: inst = 32'hc404f0b;
      37164: inst = 32'h8220000;
      37165: inst = 32'h10408000;
      37166: inst = 32'hc404f0c;
      37167: inst = 32'h8220000;
      37168: inst = 32'h10408000;
      37169: inst = 32'hc404f0d;
      37170: inst = 32'h8220000;
      37171: inst = 32'h10408000;
      37172: inst = 32'hc404f0e;
      37173: inst = 32'h8220000;
      37174: inst = 32'h10408000;
      37175: inst = 32'hc404f0f;
      37176: inst = 32'h8220000;
      37177: inst = 32'h10408000;
      37178: inst = 32'hc404f10;
      37179: inst = 32'h8220000;
      37180: inst = 32'h10408000;
      37181: inst = 32'hc404f11;
      37182: inst = 32'h8220000;
      37183: inst = 32'h10408000;
      37184: inst = 32'hc404f12;
      37185: inst = 32'h8220000;
      37186: inst = 32'h10408000;
      37187: inst = 32'hc404f13;
      37188: inst = 32'h8220000;
      37189: inst = 32'h10408000;
      37190: inst = 32'hc404f14;
      37191: inst = 32'h8220000;
      37192: inst = 32'h10408000;
      37193: inst = 32'hc404f15;
      37194: inst = 32'h8220000;
      37195: inst = 32'h10408000;
      37196: inst = 32'hc404f16;
      37197: inst = 32'h8220000;
      37198: inst = 32'h10408000;
      37199: inst = 32'hc404f17;
      37200: inst = 32'h8220000;
      37201: inst = 32'h10408000;
      37202: inst = 32'hc404f1b;
      37203: inst = 32'h8220000;
      37204: inst = 32'h10408000;
      37205: inst = 32'hc404f1c;
      37206: inst = 32'h8220000;
      37207: inst = 32'h10408000;
      37208: inst = 32'hc404f1d;
      37209: inst = 32'h8220000;
      37210: inst = 32'h10408000;
      37211: inst = 32'hc404f1e;
      37212: inst = 32'h8220000;
      37213: inst = 32'h10408000;
      37214: inst = 32'hc404f1f;
      37215: inst = 32'h8220000;
      37216: inst = 32'h10408000;
      37217: inst = 32'hc404f20;
      37218: inst = 32'h8220000;
      37219: inst = 32'h10408000;
      37220: inst = 32'hc404f21;
      37221: inst = 32'h8220000;
      37222: inst = 32'h10408000;
      37223: inst = 32'hc404f22;
      37224: inst = 32'h8220000;
      37225: inst = 32'h10408000;
      37226: inst = 32'hc404f23;
      37227: inst = 32'h8220000;
      37228: inst = 32'h10408000;
      37229: inst = 32'hc404f24;
      37230: inst = 32'h8220000;
      37231: inst = 32'h10408000;
      37232: inst = 32'hc404f25;
      37233: inst = 32'h8220000;
      37234: inst = 32'h10408000;
      37235: inst = 32'hc404f26;
      37236: inst = 32'h8220000;
      37237: inst = 32'h10408000;
      37238: inst = 32'hc404f27;
      37239: inst = 32'h8220000;
      37240: inst = 32'h10408000;
      37241: inst = 32'hc404f28;
      37242: inst = 32'h8220000;
      37243: inst = 32'h10408000;
      37244: inst = 32'hc404f29;
      37245: inst = 32'h8220000;
      37246: inst = 32'h10408000;
      37247: inst = 32'hc404f2a;
      37248: inst = 32'h8220000;
      37249: inst = 32'h10408000;
      37250: inst = 32'hc404f2b;
      37251: inst = 32'h8220000;
      37252: inst = 32'h10408000;
      37253: inst = 32'hc404f2c;
      37254: inst = 32'h8220000;
      37255: inst = 32'h10408000;
      37256: inst = 32'hc404f2d;
      37257: inst = 32'h8220000;
      37258: inst = 32'h10408000;
      37259: inst = 32'hc404f2e;
      37260: inst = 32'h8220000;
      37261: inst = 32'h10408000;
      37262: inst = 32'hc404f2f;
      37263: inst = 32'h8220000;
      37264: inst = 32'h10408000;
      37265: inst = 32'hc404f30;
      37266: inst = 32'h8220000;
      37267: inst = 32'h10408000;
      37268: inst = 32'hc404f31;
      37269: inst = 32'h8220000;
      37270: inst = 32'h10408000;
      37271: inst = 32'hc404f32;
      37272: inst = 32'h8220000;
      37273: inst = 32'h10408000;
      37274: inst = 32'hc404f33;
      37275: inst = 32'h8220000;
      37276: inst = 32'h10408000;
      37277: inst = 32'hc404f34;
      37278: inst = 32'h8220000;
      37279: inst = 32'h10408000;
      37280: inst = 32'hc404f35;
      37281: inst = 32'h8220000;
      37282: inst = 32'h10408000;
      37283: inst = 32'hc404f36;
      37284: inst = 32'h8220000;
      37285: inst = 32'h10408000;
      37286: inst = 32'hc404f37;
      37287: inst = 32'h8220000;
      37288: inst = 32'h10408000;
      37289: inst = 32'hc404f38;
      37290: inst = 32'h8220000;
      37291: inst = 32'h10408000;
      37292: inst = 32'hc404f39;
      37293: inst = 32'h8220000;
      37294: inst = 32'h10408000;
      37295: inst = 32'hc404f3a;
      37296: inst = 32'h8220000;
      37297: inst = 32'h10408000;
      37298: inst = 32'hc404f3b;
      37299: inst = 32'h8220000;
      37300: inst = 32'h10408000;
      37301: inst = 32'hc404f3c;
      37302: inst = 32'h8220000;
      37303: inst = 32'h10408000;
      37304: inst = 32'hc404f43;
      37305: inst = 32'h8220000;
      37306: inst = 32'h10408000;
      37307: inst = 32'hc404f44;
      37308: inst = 32'h8220000;
      37309: inst = 32'h10408000;
      37310: inst = 32'hc404f45;
      37311: inst = 32'h8220000;
      37312: inst = 32'h10408000;
      37313: inst = 32'hc404f46;
      37314: inst = 32'h8220000;
      37315: inst = 32'h10408000;
      37316: inst = 32'hc404f47;
      37317: inst = 32'h8220000;
      37318: inst = 32'h10408000;
      37319: inst = 32'hc404f48;
      37320: inst = 32'h8220000;
      37321: inst = 32'h10408000;
      37322: inst = 32'hc404f49;
      37323: inst = 32'h8220000;
      37324: inst = 32'h10408000;
      37325: inst = 32'hc404f4a;
      37326: inst = 32'h8220000;
      37327: inst = 32'h10408000;
      37328: inst = 32'hc404f4b;
      37329: inst = 32'h8220000;
      37330: inst = 32'h10408000;
      37331: inst = 32'hc404f4c;
      37332: inst = 32'h8220000;
      37333: inst = 32'h10408000;
      37334: inst = 32'hc404f4d;
      37335: inst = 32'h8220000;
      37336: inst = 32'h10408000;
      37337: inst = 32'hc404f4e;
      37338: inst = 32'h8220000;
      37339: inst = 32'h10408000;
      37340: inst = 32'hc404f4f;
      37341: inst = 32'h8220000;
      37342: inst = 32'h10408000;
      37343: inst = 32'hc404f50;
      37344: inst = 32'h8220000;
      37345: inst = 32'h10408000;
      37346: inst = 32'hc404f51;
      37347: inst = 32'h8220000;
      37348: inst = 32'h10408000;
      37349: inst = 32'hc404f52;
      37350: inst = 32'h8220000;
      37351: inst = 32'h10408000;
      37352: inst = 32'hc404f53;
      37353: inst = 32'h8220000;
      37354: inst = 32'h10408000;
      37355: inst = 32'hc404f54;
      37356: inst = 32'h8220000;
      37357: inst = 32'h10408000;
      37358: inst = 32'hc404f55;
      37359: inst = 32'h8220000;
      37360: inst = 32'h10408000;
      37361: inst = 32'hc404f56;
      37362: inst = 32'h8220000;
      37363: inst = 32'h10408000;
      37364: inst = 32'hc404f57;
      37365: inst = 32'h8220000;
      37366: inst = 32'h10408000;
      37367: inst = 32'hc404f58;
      37368: inst = 32'h8220000;
      37369: inst = 32'h10408000;
      37370: inst = 32'hc404f59;
      37371: inst = 32'h8220000;
      37372: inst = 32'h10408000;
      37373: inst = 32'hc404f5a;
      37374: inst = 32'h8220000;
      37375: inst = 32'h10408000;
      37376: inst = 32'hc404f5b;
      37377: inst = 32'h8220000;
      37378: inst = 32'h10408000;
      37379: inst = 32'hc404f5c;
      37380: inst = 32'h8220000;
      37381: inst = 32'h10408000;
      37382: inst = 32'hc404f5d;
      37383: inst = 32'h8220000;
      37384: inst = 32'h10408000;
      37385: inst = 32'hc404f5e;
      37386: inst = 32'h8220000;
      37387: inst = 32'h10408000;
      37388: inst = 32'hc404f5f;
      37389: inst = 32'h8220000;
      37390: inst = 32'h10408000;
      37391: inst = 32'hc404f60;
      37392: inst = 32'h8220000;
      37393: inst = 32'h10408000;
      37394: inst = 32'hc404f61;
      37395: inst = 32'h8220000;
      37396: inst = 32'h10408000;
      37397: inst = 32'hc404f62;
      37398: inst = 32'h8220000;
      37399: inst = 32'h10408000;
      37400: inst = 32'hc404f63;
      37401: inst = 32'h8220000;
      37402: inst = 32'h10408000;
      37403: inst = 32'hc404f64;
      37404: inst = 32'h8220000;
      37405: inst = 32'h10408000;
      37406: inst = 32'hc404f65;
      37407: inst = 32'h8220000;
      37408: inst = 32'h10408000;
      37409: inst = 32'hc404f66;
      37410: inst = 32'h8220000;
      37411: inst = 32'h10408000;
      37412: inst = 32'hc404f67;
      37413: inst = 32'h8220000;
      37414: inst = 32'h10408000;
      37415: inst = 32'hc404f68;
      37416: inst = 32'h8220000;
      37417: inst = 32'h10408000;
      37418: inst = 32'hc404f69;
      37419: inst = 32'h8220000;
      37420: inst = 32'h10408000;
      37421: inst = 32'hc404f6a;
      37422: inst = 32'h8220000;
      37423: inst = 32'h10408000;
      37424: inst = 32'hc404f6b;
      37425: inst = 32'h8220000;
      37426: inst = 32'h10408000;
      37427: inst = 32'hc404f6c;
      37428: inst = 32'h8220000;
      37429: inst = 32'h10408000;
      37430: inst = 32'hc404f6d;
      37431: inst = 32'h8220000;
      37432: inst = 32'h10408000;
      37433: inst = 32'hc404f6e;
      37434: inst = 32'h8220000;
      37435: inst = 32'h10408000;
      37436: inst = 32'hc404f6f;
      37437: inst = 32'h8220000;
      37438: inst = 32'h10408000;
      37439: inst = 32'hc404f70;
      37440: inst = 32'h8220000;
      37441: inst = 32'h10408000;
      37442: inst = 32'hc404f71;
      37443: inst = 32'h8220000;
      37444: inst = 32'h10408000;
      37445: inst = 32'hc404f72;
      37446: inst = 32'h8220000;
      37447: inst = 32'h10408000;
      37448: inst = 32'hc404f73;
      37449: inst = 32'h8220000;
      37450: inst = 32'h10408000;
      37451: inst = 32'hc404f74;
      37452: inst = 32'h8220000;
      37453: inst = 32'h10408000;
      37454: inst = 32'hc404f75;
      37455: inst = 32'h8220000;
      37456: inst = 32'h10408000;
      37457: inst = 32'hc404f76;
      37458: inst = 32'h8220000;
      37459: inst = 32'h10408000;
      37460: inst = 32'hc404f77;
      37461: inst = 32'h8220000;
      37462: inst = 32'h10408000;
      37463: inst = 32'hc404f7b;
      37464: inst = 32'h8220000;
      37465: inst = 32'h10408000;
      37466: inst = 32'hc404f7c;
      37467: inst = 32'h8220000;
      37468: inst = 32'h10408000;
      37469: inst = 32'hc404f7d;
      37470: inst = 32'h8220000;
      37471: inst = 32'h10408000;
      37472: inst = 32'hc404f7e;
      37473: inst = 32'h8220000;
      37474: inst = 32'h10408000;
      37475: inst = 32'hc404f7f;
      37476: inst = 32'h8220000;
      37477: inst = 32'h10408000;
      37478: inst = 32'hc404f80;
      37479: inst = 32'h8220000;
      37480: inst = 32'h10408000;
      37481: inst = 32'hc404f81;
      37482: inst = 32'h8220000;
      37483: inst = 32'h10408000;
      37484: inst = 32'hc404f82;
      37485: inst = 32'h8220000;
      37486: inst = 32'h10408000;
      37487: inst = 32'hc404f83;
      37488: inst = 32'h8220000;
      37489: inst = 32'h10408000;
      37490: inst = 32'hc404f84;
      37491: inst = 32'h8220000;
      37492: inst = 32'h10408000;
      37493: inst = 32'hc404f85;
      37494: inst = 32'h8220000;
      37495: inst = 32'h10408000;
      37496: inst = 32'hc404f86;
      37497: inst = 32'h8220000;
      37498: inst = 32'h10408000;
      37499: inst = 32'hc404f87;
      37500: inst = 32'h8220000;
      37501: inst = 32'h10408000;
      37502: inst = 32'hc404f88;
      37503: inst = 32'h8220000;
      37504: inst = 32'h10408000;
      37505: inst = 32'hc404f89;
      37506: inst = 32'h8220000;
      37507: inst = 32'h10408000;
      37508: inst = 32'hc404f8a;
      37509: inst = 32'h8220000;
      37510: inst = 32'h10408000;
      37511: inst = 32'hc404f8b;
      37512: inst = 32'h8220000;
      37513: inst = 32'h10408000;
      37514: inst = 32'hc404f8c;
      37515: inst = 32'h8220000;
      37516: inst = 32'h10408000;
      37517: inst = 32'hc404f8d;
      37518: inst = 32'h8220000;
      37519: inst = 32'h10408000;
      37520: inst = 32'hc404f8e;
      37521: inst = 32'h8220000;
      37522: inst = 32'h10408000;
      37523: inst = 32'hc404f8f;
      37524: inst = 32'h8220000;
      37525: inst = 32'h10408000;
      37526: inst = 32'hc404f90;
      37527: inst = 32'h8220000;
      37528: inst = 32'h10408000;
      37529: inst = 32'hc404f91;
      37530: inst = 32'h8220000;
      37531: inst = 32'h10408000;
      37532: inst = 32'hc404f92;
      37533: inst = 32'h8220000;
      37534: inst = 32'h10408000;
      37535: inst = 32'hc404f93;
      37536: inst = 32'h8220000;
      37537: inst = 32'h10408000;
      37538: inst = 32'hc404f94;
      37539: inst = 32'h8220000;
      37540: inst = 32'h10408000;
      37541: inst = 32'hc404f95;
      37542: inst = 32'h8220000;
      37543: inst = 32'h10408000;
      37544: inst = 32'hc404f96;
      37545: inst = 32'h8220000;
      37546: inst = 32'h10408000;
      37547: inst = 32'hc404f97;
      37548: inst = 32'h8220000;
      37549: inst = 32'h10408000;
      37550: inst = 32'hc404f98;
      37551: inst = 32'h8220000;
      37552: inst = 32'h10408000;
      37553: inst = 32'hc404f99;
      37554: inst = 32'h8220000;
      37555: inst = 32'h10408000;
      37556: inst = 32'hc404f9a;
      37557: inst = 32'h8220000;
      37558: inst = 32'h10408000;
      37559: inst = 32'hc404f9b;
      37560: inst = 32'h8220000;
      37561: inst = 32'h10408000;
      37562: inst = 32'hc404f9c;
      37563: inst = 32'h8220000;
      37564: inst = 32'h10408000;
      37565: inst = 32'hc404fa3;
      37566: inst = 32'h8220000;
      37567: inst = 32'h10408000;
      37568: inst = 32'hc404fa4;
      37569: inst = 32'h8220000;
      37570: inst = 32'h10408000;
      37571: inst = 32'hc404fa5;
      37572: inst = 32'h8220000;
      37573: inst = 32'h10408000;
      37574: inst = 32'hc404fa6;
      37575: inst = 32'h8220000;
      37576: inst = 32'h10408000;
      37577: inst = 32'hc404fa7;
      37578: inst = 32'h8220000;
      37579: inst = 32'h10408000;
      37580: inst = 32'hc404fa8;
      37581: inst = 32'h8220000;
      37582: inst = 32'h10408000;
      37583: inst = 32'hc404fa9;
      37584: inst = 32'h8220000;
      37585: inst = 32'h10408000;
      37586: inst = 32'hc404faa;
      37587: inst = 32'h8220000;
      37588: inst = 32'h10408000;
      37589: inst = 32'hc404fab;
      37590: inst = 32'h8220000;
      37591: inst = 32'h10408000;
      37592: inst = 32'hc404fac;
      37593: inst = 32'h8220000;
      37594: inst = 32'h10408000;
      37595: inst = 32'hc404fad;
      37596: inst = 32'h8220000;
      37597: inst = 32'h10408000;
      37598: inst = 32'hc404fae;
      37599: inst = 32'h8220000;
      37600: inst = 32'h10408000;
      37601: inst = 32'hc404faf;
      37602: inst = 32'h8220000;
      37603: inst = 32'h10408000;
      37604: inst = 32'hc404fb0;
      37605: inst = 32'h8220000;
      37606: inst = 32'h10408000;
      37607: inst = 32'hc404fb1;
      37608: inst = 32'h8220000;
      37609: inst = 32'h10408000;
      37610: inst = 32'hc404fb2;
      37611: inst = 32'h8220000;
      37612: inst = 32'h10408000;
      37613: inst = 32'hc404fb3;
      37614: inst = 32'h8220000;
      37615: inst = 32'h10408000;
      37616: inst = 32'hc404fb4;
      37617: inst = 32'h8220000;
      37618: inst = 32'h10408000;
      37619: inst = 32'hc404fb5;
      37620: inst = 32'h8220000;
      37621: inst = 32'h10408000;
      37622: inst = 32'hc404fb6;
      37623: inst = 32'h8220000;
      37624: inst = 32'h10408000;
      37625: inst = 32'hc404fb7;
      37626: inst = 32'h8220000;
      37627: inst = 32'h10408000;
      37628: inst = 32'hc404fb8;
      37629: inst = 32'h8220000;
      37630: inst = 32'h10408000;
      37631: inst = 32'hc404fb9;
      37632: inst = 32'h8220000;
      37633: inst = 32'h10408000;
      37634: inst = 32'hc404fba;
      37635: inst = 32'h8220000;
      37636: inst = 32'h10408000;
      37637: inst = 32'hc404fbb;
      37638: inst = 32'h8220000;
      37639: inst = 32'h10408000;
      37640: inst = 32'hc404fbc;
      37641: inst = 32'h8220000;
      37642: inst = 32'h10408000;
      37643: inst = 32'hc404fbd;
      37644: inst = 32'h8220000;
      37645: inst = 32'h10408000;
      37646: inst = 32'hc404fbe;
      37647: inst = 32'h8220000;
      37648: inst = 32'h10408000;
      37649: inst = 32'hc404fbf;
      37650: inst = 32'h8220000;
      37651: inst = 32'h10408000;
      37652: inst = 32'hc404fc0;
      37653: inst = 32'h8220000;
      37654: inst = 32'h10408000;
      37655: inst = 32'hc404fc1;
      37656: inst = 32'h8220000;
      37657: inst = 32'h10408000;
      37658: inst = 32'hc404fc2;
      37659: inst = 32'h8220000;
      37660: inst = 32'h10408000;
      37661: inst = 32'hc404fc3;
      37662: inst = 32'h8220000;
      37663: inst = 32'h10408000;
      37664: inst = 32'hc404fc4;
      37665: inst = 32'h8220000;
      37666: inst = 32'h10408000;
      37667: inst = 32'hc404fc5;
      37668: inst = 32'h8220000;
      37669: inst = 32'h10408000;
      37670: inst = 32'hc404fc6;
      37671: inst = 32'h8220000;
      37672: inst = 32'h10408000;
      37673: inst = 32'hc404fc7;
      37674: inst = 32'h8220000;
      37675: inst = 32'h10408000;
      37676: inst = 32'hc404fc8;
      37677: inst = 32'h8220000;
      37678: inst = 32'h10408000;
      37679: inst = 32'hc404fc9;
      37680: inst = 32'h8220000;
      37681: inst = 32'h10408000;
      37682: inst = 32'hc404fca;
      37683: inst = 32'h8220000;
      37684: inst = 32'h10408000;
      37685: inst = 32'hc404fcb;
      37686: inst = 32'h8220000;
      37687: inst = 32'h10408000;
      37688: inst = 32'hc404fcc;
      37689: inst = 32'h8220000;
      37690: inst = 32'h10408000;
      37691: inst = 32'hc404fcd;
      37692: inst = 32'h8220000;
      37693: inst = 32'h10408000;
      37694: inst = 32'hc404fce;
      37695: inst = 32'h8220000;
      37696: inst = 32'h10408000;
      37697: inst = 32'hc404fcf;
      37698: inst = 32'h8220000;
      37699: inst = 32'h10408000;
      37700: inst = 32'hc404fd0;
      37701: inst = 32'h8220000;
      37702: inst = 32'h10408000;
      37703: inst = 32'hc404fd1;
      37704: inst = 32'h8220000;
      37705: inst = 32'h10408000;
      37706: inst = 32'hc404fd2;
      37707: inst = 32'h8220000;
      37708: inst = 32'h10408000;
      37709: inst = 32'hc404fd3;
      37710: inst = 32'h8220000;
      37711: inst = 32'h10408000;
      37712: inst = 32'hc404fd4;
      37713: inst = 32'h8220000;
      37714: inst = 32'h10408000;
      37715: inst = 32'hc404fd5;
      37716: inst = 32'h8220000;
      37717: inst = 32'h10408000;
      37718: inst = 32'hc404fd6;
      37719: inst = 32'h8220000;
      37720: inst = 32'h10408000;
      37721: inst = 32'hc404fd7;
      37722: inst = 32'h8220000;
      37723: inst = 32'h10408000;
      37724: inst = 32'hc404fdb;
      37725: inst = 32'h8220000;
      37726: inst = 32'h10408000;
      37727: inst = 32'hc404fdc;
      37728: inst = 32'h8220000;
      37729: inst = 32'h10408000;
      37730: inst = 32'hc404fdd;
      37731: inst = 32'h8220000;
      37732: inst = 32'h10408000;
      37733: inst = 32'hc404fde;
      37734: inst = 32'h8220000;
      37735: inst = 32'h10408000;
      37736: inst = 32'hc404fdf;
      37737: inst = 32'h8220000;
      37738: inst = 32'h10408000;
      37739: inst = 32'hc404fe0;
      37740: inst = 32'h8220000;
      37741: inst = 32'h10408000;
      37742: inst = 32'hc404fe1;
      37743: inst = 32'h8220000;
      37744: inst = 32'h10408000;
      37745: inst = 32'hc404fe2;
      37746: inst = 32'h8220000;
      37747: inst = 32'h10408000;
      37748: inst = 32'hc404fe3;
      37749: inst = 32'h8220000;
      37750: inst = 32'h10408000;
      37751: inst = 32'hc404fe4;
      37752: inst = 32'h8220000;
      37753: inst = 32'h10408000;
      37754: inst = 32'hc404fe5;
      37755: inst = 32'h8220000;
      37756: inst = 32'h10408000;
      37757: inst = 32'hc404fe6;
      37758: inst = 32'h8220000;
      37759: inst = 32'h10408000;
      37760: inst = 32'hc404fe7;
      37761: inst = 32'h8220000;
      37762: inst = 32'h10408000;
      37763: inst = 32'hc404fe8;
      37764: inst = 32'h8220000;
      37765: inst = 32'h10408000;
      37766: inst = 32'hc404fe9;
      37767: inst = 32'h8220000;
      37768: inst = 32'h10408000;
      37769: inst = 32'hc404fea;
      37770: inst = 32'h8220000;
      37771: inst = 32'h10408000;
      37772: inst = 32'hc404feb;
      37773: inst = 32'h8220000;
      37774: inst = 32'h10408000;
      37775: inst = 32'hc404fec;
      37776: inst = 32'h8220000;
      37777: inst = 32'h10408000;
      37778: inst = 32'hc404fed;
      37779: inst = 32'h8220000;
      37780: inst = 32'h10408000;
      37781: inst = 32'hc404fee;
      37782: inst = 32'h8220000;
      37783: inst = 32'h10408000;
      37784: inst = 32'hc404fef;
      37785: inst = 32'h8220000;
      37786: inst = 32'h10408000;
      37787: inst = 32'hc404ff0;
      37788: inst = 32'h8220000;
      37789: inst = 32'h10408000;
      37790: inst = 32'hc404ff1;
      37791: inst = 32'h8220000;
      37792: inst = 32'h10408000;
      37793: inst = 32'hc404ff2;
      37794: inst = 32'h8220000;
      37795: inst = 32'h10408000;
      37796: inst = 32'hc404ff3;
      37797: inst = 32'h8220000;
      37798: inst = 32'h10408000;
      37799: inst = 32'hc404ff4;
      37800: inst = 32'h8220000;
      37801: inst = 32'h10408000;
      37802: inst = 32'hc404ff5;
      37803: inst = 32'h8220000;
      37804: inst = 32'h10408000;
      37805: inst = 32'hc404ff6;
      37806: inst = 32'h8220000;
      37807: inst = 32'h10408000;
      37808: inst = 32'hc404ff7;
      37809: inst = 32'h8220000;
      37810: inst = 32'h10408000;
      37811: inst = 32'hc404ff8;
      37812: inst = 32'h8220000;
      37813: inst = 32'h10408000;
      37814: inst = 32'hc404ff9;
      37815: inst = 32'h8220000;
      37816: inst = 32'h10408000;
      37817: inst = 32'hc404ffa;
      37818: inst = 32'h8220000;
      37819: inst = 32'h10408000;
      37820: inst = 32'hc404ffb;
      37821: inst = 32'h8220000;
      37822: inst = 32'h10408000;
      37823: inst = 32'hc404ffc;
      37824: inst = 32'h8220000;
      37825: inst = 32'h10408000;
      37826: inst = 32'hc405003;
      37827: inst = 32'h8220000;
      37828: inst = 32'h10408000;
      37829: inst = 32'hc405004;
      37830: inst = 32'h8220000;
      37831: inst = 32'h10408000;
      37832: inst = 32'hc405005;
      37833: inst = 32'h8220000;
      37834: inst = 32'h10408000;
      37835: inst = 32'hc405006;
      37836: inst = 32'h8220000;
      37837: inst = 32'h10408000;
      37838: inst = 32'hc405007;
      37839: inst = 32'h8220000;
      37840: inst = 32'h10408000;
      37841: inst = 32'hc405008;
      37842: inst = 32'h8220000;
      37843: inst = 32'h10408000;
      37844: inst = 32'hc405009;
      37845: inst = 32'h8220000;
      37846: inst = 32'h10408000;
      37847: inst = 32'hc40500a;
      37848: inst = 32'h8220000;
      37849: inst = 32'h10408000;
      37850: inst = 32'hc40500b;
      37851: inst = 32'h8220000;
      37852: inst = 32'h10408000;
      37853: inst = 32'hc40500c;
      37854: inst = 32'h8220000;
      37855: inst = 32'h10408000;
      37856: inst = 32'hc40500d;
      37857: inst = 32'h8220000;
      37858: inst = 32'h10408000;
      37859: inst = 32'hc40500e;
      37860: inst = 32'h8220000;
      37861: inst = 32'h10408000;
      37862: inst = 32'hc40500f;
      37863: inst = 32'h8220000;
      37864: inst = 32'h10408000;
      37865: inst = 32'hc405010;
      37866: inst = 32'h8220000;
      37867: inst = 32'h10408000;
      37868: inst = 32'hc405011;
      37869: inst = 32'h8220000;
      37870: inst = 32'h10408000;
      37871: inst = 32'hc405012;
      37872: inst = 32'h8220000;
      37873: inst = 32'h10408000;
      37874: inst = 32'hc405013;
      37875: inst = 32'h8220000;
      37876: inst = 32'h10408000;
      37877: inst = 32'hc405014;
      37878: inst = 32'h8220000;
      37879: inst = 32'h10408000;
      37880: inst = 32'hc405015;
      37881: inst = 32'h8220000;
      37882: inst = 32'h10408000;
      37883: inst = 32'hc405016;
      37884: inst = 32'h8220000;
      37885: inst = 32'h10408000;
      37886: inst = 32'hc405017;
      37887: inst = 32'h8220000;
      37888: inst = 32'h10408000;
      37889: inst = 32'hc405018;
      37890: inst = 32'h8220000;
      37891: inst = 32'h10408000;
      37892: inst = 32'hc405019;
      37893: inst = 32'h8220000;
      37894: inst = 32'h10408000;
      37895: inst = 32'hc40501a;
      37896: inst = 32'h8220000;
      37897: inst = 32'h10408000;
      37898: inst = 32'hc40501b;
      37899: inst = 32'h8220000;
      37900: inst = 32'h10408000;
      37901: inst = 32'hc40501c;
      37902: inst = 32'h8220000;
      37903: inst = 32'h10408000;
      37904: inst = 32'hc40501d;
      37905: inst = 32'h8220000;
      37906: inst = 32'h10408000;
      37907: inst = 32'hc40501e;
      37908: inst = 32'h8220000;
      37909: inst = 32'h10408000;
      37910: inst = 32'hc40501f;
      37911: inst = 32'h8220000;
      37912: inst = 32'h10408000;
      37913: inst = 32'hc405020;
      37914: inst = 32'h8220000;
      37915: inst = 32'h10408000;
      37916: inst = 32'hc405021;
      37917: inst = 32'h8220000;
      37918: inst = 32'h10408000;
      37919: inst = 32'hc405022;
      37920: inst = 32'h8220000;
      37921: inst = 32'h10408000;
      37922: inst = 32'hc405023;
      37923: inst = 32'h8220000;
      37924: inst = 32'h10408000;
      37925: inst = 32'hc405024;
      37926: inst = 32'h8220000;
      37927: inst = 32'h10408000;
      37928: inst = 32'hc405025;
      37929: inst = 32'h8220000;
      37930: inst = 32'h10408000;
      37931: inst = 32'hc405026;
      37932: inst = 32'h8220000;
      37933: inst = 32'h10408000;
      37934: inst = 32'hc405027;
      37935: inst = 32'h8220000;
      37936: inst = 32'h10408000;
      37937: inst = 32'hc405028;
      37938: inst = 32'h8220000;
      37939: inst = 32'h10408000;
      37940: inst = 32'hc405029;
      37941: inst = 32'h8220000;
      37942: inst = 32'h10408000;
      37943: inst = 32'hc40502a;
      37944: inst = 32'h8220000;
      37945: inst = 32'h10408000;
      37946: inst = 32'hc40502b;
      37947: inst = 32'h8220000;
      37948: inst = 32'h10408000;
      37949: inst = 32'hc40502c;
      37950: inst = 32'h8220000;
      37951: inst = 32'h10408000;
      37952: inst = 32'hc40502d;
      37953: inst = 32'h8220000;
      37954: inst = 32'h10408000;
      37955: inst = 32'hc40502e;
      37956: inst = 32'h8220000;
      37957: inst = 32'h10408000;
      37958: inst = 32'hc40502f;
      37959: inst = 32'h8220000;
      37960: inst = 32'h10408000;
      37961: inst = 32'hc405030;
      37962: inst = 32'h8220000;
      37963: inst = 32'h10408000;
      37964: inst = 32'hc405031;
      37965: inst = 32'h8220000;
      37966: inst = 32'h10408000;
      37967: inst = 32'hc405032;
      37968: inst = 32'h8220000;
      37969: inst = 32'h10408000;
      37970: inst = 32'hc405033;
      37971: inst = 32'h8220000;
      37972: inst = 32'h10408000;
      37973: inst = 32'hc405034;
      37974: inst = 32'h8220000;
      37975: inst = 32'h10408000;
      37976: inst = 32'hc405035;
      37977: inst = 32'h8220000;
      37978: inst = 32'h10408000;
      37979: inst = 32'hc405036;
      37980: inst = 32'h8220000;
      37981: inst = 32'h10408000;
      37982: inst = 32'hc405037;
      37983: inst = 32'h8220000;
      37984: inst = 32'h10408000;
      37985: inst = 32'hc40503b;
      37986: inst = 32'h8220000;
      37987: inst = 32'h10408000;
      37988: inst = 32'hc40503c;
      37989: inst = 32'h8220000;
      37990: inst = 32'h10408000;
      37991: inst = 32'hc40503d;
      37992: inst = 32'h8220000;
      37993: inst = 32'h10408000;
      37994: inst = 32'hc40503e;
      37995: inst = 32'h8220000;
      37996: inst = 32'h10408000;
      37997: inst = 32'hc40503f;
      37998: inst = 32'h8220000;
      37999: inst = 32'h10408000;
      38000: inst = 32'hc405040;
      38001: inst = 32'h8220000;
      38002: inst = 32'h10408000;
      38003: inst = 32'hc405041;
      38004: inst = 32'h8220000;
      38005: inst = 32'h10408000;
      38006: inst = 32'hc405042;
      38007: inst = 32'h8220000;
      38008: inst = 32'h10408000;
      38009: inst = 32'hc405043;
      38010: inst = 32'h8220000;
      38011: inst = 32'h10408000;
      38012: inst = 32'hc405044;
      38013: inst = 32'h8220000;
      38014: inst = 32'h10408000;
      38015: inst = 32'hc405045;
      38016: inst = 32'h8220000;
      38017: inst = 32'h10408000;
      38018: inst = 32'hc405046;
      38019: inst = 32'h8220000;
      38020: inst = 32'h10408000;
      38021: inst = 32'hc405047;
      38022: inst = 32'h8220000;
      38023: inst = 32'h10408000;
      38024: inst = 32'hc405048;
      38025: inst = 32'h8220000;
      38026: inst = 32'h10408000;
      38027: inst = 32'hc405049;
      38028: inst = 32'h8220000;
      38029: inst = 32'h10408000;
      38030: inst = 32'hc40504a;
      38031: inst = 32'h8220000;
      38032: inst = 32'h10408000;
      38033: inst = 32'hc40504b;
      38034: inst = 32'h8220000;
      38035: inst = 32'h10408000;
      38036: inst = 32'hc40504c;
      38037: inst = 32'h8220000;
      38038: inst = 32'h10408000;
      38039: inst = 32'hc40504d;
      38040: inst = 32'h8220000;
      38041: inst = 32'h10408000;
      38042: inst = 32'hc40504e;
      38043: inst = 32'h8220000;
      38044: inst = 32'h10408000;
      38045: inst = 32'hc40504f;
      38046: inst = 32'h8220000;
      38047: inst = 32'h10408000;
      38048: inst = 32'hc405050;
      38049: inst = 32'h8220000;
      38050: inst = 32'h10408000;
      38051: inst = 32'hc405051;
      38052: inst = 32'h8220000;
      38053: inst = 32'h10408000;
      38054: inst = 32'hc405052;
      38055: inst = 32'h8220000;
      38056: inst = 32'h10408000;
      38057: inst = 32'hc405053;
      38058: inst = 32'h8220000;
      38059: inst = 32'h10408000;
      38060: inst = 32'hc405054;
      38061: inst = 32'h8220000;
      38062: inst = 32'h10408000;
      38063: inst = 32'hc405055;
      38064: inst = 32'h8220000;
      38065: inst = 32'h10408000;
      38066: inst = 32'hc405056;
      38067: inst = 32'h8220000;
      38068: inst = 32'h10408000;
      38069: inst = 32'hc405057;
      38070: inst = 32'h8220000;
      38071: inst = 32'h10408000;
      38072: inst = 32'hc405058;
      38073: inst = 32'h8220000;
      38074: inst = 32'h10408000;
      38075: inst = 32'hc405059;
      38076: inst = 32'h8220000;
      38077: inst = 32'h10408000;
      38078: inst = 32'hc40505a;
      38079: inst = 32'h8220000;
      38080: inst = 32'h10408000;
      38081: inst = 32'hc40505b;
      38082: inst = 32'h8220000;
      38083: inst = 32'h10408000;
      38084: inst = 32'hc40505c;
      38085: inst = 32'h8220000;
      38086: inst = 32'h10408000;
      38087: inst = 32'hc405063;
      38088: inst = 32'h8220000;
      38089: inst = 32'h10408000;
      38090: inst = 32'hc405064;
      38091: inst = 32'h8220000;
      38092: inst = 32'h10408000;
      38093: inst = 32'hc405065;
      38094: inst = 32'h8220000;
      38095: inst = 32'h10408000;
      38096: inst = 32'hc405066;
      38097: inst = 32'h8220000;
      38098: inst = 32'h10408000;
      38099: inst = 32'hc405067;
      38100: inst = 32'h8220000;
      38101: inst = 32'h10408000;
      38102: inst = 32'hc405068;
      38103: inst = 32'h8220000;
      38104: inst = 32'h10408000;
      38105: inst = 32'hc405069;
      38106: inst = 32'h8220000;
      38107: inst = 32'h10408000;
      38108: inst = 32'hc40506a;
      38109: inst = 32'h8220000;
      38110: inst = 32'h10408000;
      38111: inst = 32'hc40506b;
      38112: inst = 32'h8220000;
      38113: inst = 32'h10408000;
      38114: inst = 32'hc40506c;
      38115: inst = 32'h8220000;
      38116: inst = 32'h10408000;
      38117: inst = 32'hc40506d;
      38118: inst = 32'h8220000;
      38119: inst = 32'h10408000;
      38120: inst = 32'hc40506e;
      38121: inst = 32'h8220000;
      38122: inst = 32'h10408000;
      38123: inst = 32'hc40506f;
      38124: inst = 32'h8220000;
      38125: inst = 32'h10408000;
      38126: inst = 32'hc405070;
      38127: inst = 32'h8220000;
      38128: inst = 32'h10408000;
      38129: inst = 32'hc405071;
      38130: inst = 32'h8220000;
      38131: inst = 32'h10408000;
      38132: inst = 32'hc405072;
      38133: inst = 32'h8220000;
      38134: inst = 32'h10408000;
      38135: inst = 32'hc405073;
      38136: inst = 32'h8220000;
      38137: inst = 32'h10408000;
      38138: inst = 32'hc405074;
      38139: inst = 32'h8220000;
      38140: inst = 32'h10408000;
      38141: inst = 32'hc405075;
      38142: inst = 32'h8220000;
      38143: inst = 32'h10408000;
      38144: inst = 32'hc405076;
      38145: inst = 32'h8220000;
      38146: inst = 32'h10408000;
      38147: inst = 32'hc405077;
      38148: inst = 32'h8220000;
      38149: inst = 32'h10408000;
      38150: inst = 32'hc405078;
      38151: inst = 32'h8220000;
      38152: inst = 32'h10408000;
      38153: inst = 32'hc405079;
      38154: inst = 32'h8220000;
      38155: inst = 32'h10408000;
      38156: inst = 32'hc40507a;
      38157: inst = 32'h8220000;
      38158: inst = 32'h10408000;
      38159: inst = 32'hc40507b;
      38160: inst = 32'h8220000;
      38161: inst = 32'h10408000;
      38162: inst = 32'hc40507c;
      38163: inst = 32'h8220000;
      38164: inst = 32'h10408000;
      38165: inst = 32'hc40507d;
      38166: inst = 32'h8220000;
      38167: inst = 32'h10408000;
      38168: inst = 32'hc40507e;
      38169: inst = 32'h8220000;
      38170: inst = 32'h10408000;
      38171: inst = 32'hc40507f;
      38172: inst = 32'h8220000;
      38173: inst = 32'h10408000;
      38174: inst = 32'hc405080;
      38175: inst = 32'h8220000;
      38176: inst = 32'h10408000;
      38177: inst = 32'hc405081;
      38178: inst = 32'h8220000;
      38179: inst = 32'h10408000;
      38180: inst = 32'hc405082;
      38181: inst = 32'h8220000;
      38182: inst = 32'h10408000;
      38183: inst = 32'hc405083;
      38184: inst = 32'h8220000;
      38185: inst = 32'h10408000;
      38186: inst = 32'hc405084;
      38187: inst = 32'h8220000;
      38188: inst = 32'h10408000;
      38189: inst = 32'hc405085;
      38190: inst = 32'h8220000;
      38191: inst = 32'h10408000;
      38192: inst = 32'hc405086;
      38193: inst = 32'h8220000;
      38194: inst = 32'h10408000;
      38195: inst = 32'hc405087;
      38196: inst = 32'h8220000;
      38197: inst = 32'h10408000;
      38198: inst = 32'hc405088;
      38199: inst = 32'h8220000;
      38200: inst = 32'h10408000;
      38201: inst = 32'hc405089;
      38202: inst = 32'h8220000;
      38203: inst = 32'h10408000;
      38204: inst = 32'hc40508a;
      38205: inst = 32'h8220000;
      38206: inst = 32'h10408000;
      38207: inst = 32'hc40508b;
      38208: inst = 32'h8220000;
      38209: inst = 32'h10408000;
      38210: inst = 32'hc40508c;
      38211: inst = 32'h8220000;
      38212: inst = 32'h10408000;
      38213: inst = 32'hc40508d;
      38214: inst = 32'h8220000;
      38215: inst = 32'h10408000;
      38216: inst = 32'hc40508e;
      38217: inst = 32'h8220000;
      38218: inst = 32'h10408000;
      38219: inst = 32'hc40508f;
      38220: inst = 32'h8220000;
      38221: inst = 32'h10408000;
      38222: inst = 32'hc405090;
      38223: inst = 32'h8220000;
      38224: inst = 32'h10408000;
      38225: inst = 32'hc405091;
      38226: inst = 32'h8220000;
      38227: inst = 32'h10408000;
      38228: inst = 32'hc405092;
      38229: inst = 32'h8220000;
      38230: inst = 32'h10408000;
      38231: inst = 32'hc405093;
      38232: inst = 32'h8220000;
      38233: inst = 32'h10408000;
      38234: inst = 32'hc405094;
      38235: inst = 32'h8220000;
      38236: inst = 32'h10408000;
      38237: inst = 32'hc405095;
      38238: inst = 32'h8220000;
      38239: inst = 32'h10408000;
      38240: inst = 32'hc405096;
      38241: inst = 32'h8220000;
      38242: inst = 32'h10408000;
      38243: inst = 32'hc405097;
      38244: inst = 32'h8220000;
      38245: inst = 32'h10408000;
      38246: inst = 32'hc4050c3;
      38247: inst = 32'h8220000;
      38248: inst = 32'h10408000;
      38249: inst = 32'hc4050c4;
      38250: inst = 32'h8220000;
      38251: inst = 32'h10408000;
      38252: inst = 32'hc4050c5;
      38253: inst = 32'h8220000;
      38254: inst = 32'h10408000;
      38255: inst = 32'hc4050c6;
      38256: inst = 32'h8220000;
      38257: inst = 32'h10408000;
      38258: inst = 32'hc4050c7;
      38259: inst = 32'h8220000;
      38260: inst = 32'h10408000;
      38261: inst = 32'hc4050c8;
      38262: inst = 32'h8220000;
      38263: inst = 32'h10408000;
      38264: inst = 32'hc4050c9;
      38265: inst = 32'h8220000;
      38266: inst = 32'h10408000;
      38267: inst = 32'hc4050ca;
      38268: inst = 32'h8220000;
      38269: inst = 32'h10408000;
      38270: inst = 32'hc4050cb;
      38271: inst = 32'h8220000;
      38272: inst = 32'h10408000;
      38273: inst = 32'hc4050cc;
      38274: inst = 32'h8220000;
      38275: inst = 32'h10408000;
      38276: inst = 32'hc4050cd;
      38277: inst = 32'h8220000;
      38278: inst = 32'h10408000;
      38279: inst = 32'hc4050ce;
      38280: inst = 32'h8220000;
      38281: inst = 32'h10408000;
      38282: inst = 32'hc4050cf;
      38283: inst = 32'h8220000;
      38284: inst = 32'h10408000;
      38285: inst = 32'hc4050d0;
      38286: inst = 32'h8220000;
      38287: inst = 32'h10408000;
      38288: inst = 32'hc4050d1;
      38289: inst = 32'h8220000;
      38290: inst = 32'h10408000;
      38291: inst = 32'hc4050d2;
      38292: inst = 32'h8220000;
      38293: inst = 32'h10408000;
      38294: inst = 32'hc4050d3;
      38295: inst = 32'h8220000;
      38296: inst = 32'h10408000;
      38297: inst = 32'hc4050d4;
      38298: inst = 32'h8220000;
      38299: inst = 32'h10408000;
      38300: inst = 32'hc4050d5;
      38301: inst = 32'h8220000;
      38302: inst = 32'h10408000;
      38303: inst = 32'hc4050d6;
      38304: inst = 32'h8220000;
      38305: inst = 32'h10408000;
      38306: inst = 32'hc4050d7;
      38307: inst = 32'h8220000;
      38308: inst = 32'h10408000;
      38309: inst = 32'hc4050d8;
      38310: inst = 32'h8220000;
      38311: inst = 32'h10408000;
      38312: inst = 32'hc4050d9;
      38313: inst = 32'h8220000;
      38314: inst = 32'h10408000;
      38315: inst = 32'hc4050da;
      38316: inst = 32'h8220000;
      38317: inst = 32'h10408000;
      38318: inst = 32'hc4050db;
      38319: inst = 32'h8220000;
      38320: inst = 32'h10408000;
      38321: inst = 32'hc4050dc;
      38322: inst = 32'h8220000;
      38323: inst = 32'h10408000;
      38324: inst = 32'hc4050dd;
      38325: inst = 32'h8220000;
      38326: inst = 32'h10408000;
      38327: inst = 32'hc4050de;
      38328: inst = 32'h8220000;
      38329: inst = 32'h10408000;
      38330: inst = 32'hc4050df;
      38331: inst = 32'h8220000;
      38332: inst = 32'h10408000;
      38333: inst = 32'hc4050e0;
      38334: inst = 32'h8220000;
      38335: inst = 32'h10408000;
      38336: inst = 32'hc4050e1;
      38337: inst = 32'h8220000;
      38338: inst = 32'h10408000;
      38339: inst = 32'hc4050e2;
      38340: inst = 32'h8220000;
      38341: inst = 32'h10408000;
      38342: inst = 32'hc4050e3;
      38343: inst = 32'h8220000;
      38344: inst = 32'h10408000;
      38345: inst = 32'hc4050e4;
      38346: inst = 32'h8220000;
      38347: inst = 32'h10408000;
      38348: inst = 32'hc4050e5;
      38349: inst = 32'h8220000;
      38350: inst = 32'h10408000;
      38351: inst = 32'hc4050e6;
      38352: inst = 32'h8220000;
      38353: inst = 32'h10408000;
      38354: inst = 32'hc4050e7;
      38355: inst = 32'h8220000;
      38356: inst = 32'h10408000;
      38357: inst = 32'hc4050e8;
      38358: inst = 32'h8220000;
      38359: inst = 32'h10408000;
      38360: inst = 32'hc4050e9;
      38361: inst = 32'h8220000;
      38362: inst = 32'h10408000;
      38363: inst = 32'hc4050ea;
      38364: inst = 32'h8220000;
      38365: inst = 32'h10408000;
      38366: inst = 32'hc4050eb;
      38367: inst = 32'h8220000;
      38368: inst = 32'h10408000;
      38369: inst = 32'hc4050ec;
      38370: inst = 32'h8220000;
      38371: inst = 32'h10408000;
      38372: inst = 32'hc4050ed;
      38373: inst = 32'h8220000;
      38374: inst = 32'h10408000;
      38375: inst = 32'hc4050ee;
      38376: inst = 32'h8220000;
      38377: inst = 32'h10408000;
      38378: inst = 32'hc4050ef;
      38379: inst = 32'h8220000;
      38380: inst = 32'h10408000;
      38381: inst = 32'hc4050f0;
      38382: inst = 32'h8220000;
      38383: inst = 32'h10408000;
      38384: inst = 32'hc4050f1;
      38385: inst = 32'h8220000;
      38386: inst = 32'h10408000;
      38387: inst = 32'hc4050f2;
      38388: inst = 32'h8220000;
      38389: inst = 32'h10408000;
      38390: inst = 32'hc4050f3;
      38391: inst = 32'h8220000;
      38392: inst = 32'h10408000;
      38393: inst = 32'hc4050f4;
      38394: inst = 32'h8220000;
      38395: inst = 32'h10408000;
      38396: inst = 32'hc4050f5;
      38397: inst = 32'h8220000;
      38398: inst = 32'h10408000;
      38399: inst = 32'hc4050f6;
      38400: inst = 32'h8220000;
      38401: inst = 32'h10408000;
      38402: inst = 32'hc4050f7;
      38403: inst = 32'h8220000;
      38404: inst = 32'h10408000;
      38405: inst = 32'hc405123;
      38406: inst = 32'h8220000;
      38407: inst = 32'h10408000;
      38408: inst = 32'hc405124;
      38409: inst = 32'h8220000;
      38410: inst = 32'h10408000;
      38411: inst = 32'hc405125;
      38412: inst = 32'h8220000;
      38413: inst = 32'h10408000;
      38414: inst = 32'hc405126;
      38415: inst = 32'h8220000;
      38416: inst = 32'h10408000;
      38417: inst = 32'hc405127;
      38418: inst = 32'h8220000;
      38419: inst = 32'h10408000;
      38420: inst = 32'hc405128;
      38421: inst = 32'h8220000;
      38422: inst = 32'h10408000;
      38423: inst = 32'hc405129;
      38424: inst = 32'h8220000;
      38425: inst = 32'h10408000;
      38426: inst = 32'hc40512a;
      38427: inst = 32'h8220000;
      38428: inst = 32'h10408000;
      38429: inst = 32'hc40512b;
      38430: inst = 32'h8220000;
      38431: inst = 32'h10408000;
      38432: inst = 32'hc40512c;
      38433: inst = 32'h8220000;
      38434: inst = 32'h10408000;
      38435: inst = 32'hc40512d;
      38436: inst = 32'h8220000;
      38437: inst = 32'h10408000;
      38438: inst = 32'hc40512e;
      38439: inst = 32'h8220000;
      38440: inst = 32'h10408000;
      38441: inst = 32'hc40512f;
      38442: inst = 32'h8220000;
      38443: inst = 32'h10408000;
      38444: inst = 32'hc405130;
      38445: inst = 32'h8220000;
      38446: inst = 32'h10408000;
      38447: inst = 32'hc405131;
      38448: inst = 32'h8220000;
      38449: inst = 32'h10408000;
      38450: inst = 32'hc405132;
      38451: inst = 32'h8220000;
      38452: inst = 32'h10408000;
      38453: inst = 32'hc405133;
      38454: inst = 32'h8220000;
      38455: inst = 32'h10408000;
      38456: inst = 32'hc405134;
      38457: inst = 32'h8220000;
      38458: inst = 32'h10408000;
      38459: inst = 32'hc405135;
      38460: inst = 32'h8220000;
      38461: inst = 32'h10408000;
      38462: inst = 32'hc405139;
      38463: inst = 32'h8220000;
      38464: inst = 32'h10408000;
      38465: inst = 32'hc40513a;
      38466: inst = 32'h8220000;
      38467: inst = 32'h10408000;
      38468: inst = 32'hc40513b;
      38469: inst = 32'h8220000;
      38470: inst = 32'h10408000;
      38471: inst = 32'hc40513c;
      38472: inst = 32'h8220000;
      38473: inst = 32'h10408000;
      38474: inst = 32'hc40513d;
      38475: inst = 32'h8220000;
      38476: inst = 32'h10408000;
      38477: inst = 32'hc40513e;
      38478: inst = 32'h8220000;
      38479: inst = 32'h10408000;
      38480: inst = 32'hc40513f;
      38481: inst = 32'h8220000;
      38482: inst = 32'h10408000;
      38483: inst = 32'hc405140;
      38484: inst = 32'h8220000;
      38485: inst = 32'h10408000;
      38486: inst = 32'hc405141;
      38487: inst = 32'h8220000;
      38488: inst = 32'h10408000;
      38489: inst = 32'hc405142;
      38490: inst = 32'h8220000;
      38491: inst = 32'h10408000;
      38492: inst = 32'hc405143;
      38493: inst = 32'h8220000;
      38494: inst = 32'h10408000;
      38495: inst = 32'hc405144;
      38496: inst = 32'h8220000;
      38497: inst = 32'h10408000;
      38498: inst = 32'hc405145;
      38499: inst = 32'h8220000;
      38500: inst = 32'h10408000;
      38501: inst = 32'hc405146;
      38502: inst = 32'h8220000;
      38503: inst = 32'h10408000;
      38504: inst = 32'hc405147;
      38505: inst = 32'h8220000;
      38506: inst = 32'h10408000;
      38507: inst = 32'hc405148;
      38508: inst = 32'h8220000;
      38509: inst = 32'h10408000;
      38510: inst = 32'hc405149;
      38511: inst = 32'h8220000;
      38512: inst = 32'h10408000;
      38513: inst = 32'hc40514a;
      38514: inst = 32'h8220000;
      38515: inst = 32'h10408000;
      38516: inst = 32'hc40514b;
      38517: inst = 32'h8220000;
      38518: inst = 32'h10408000;
      38519: inst = 32'hc40514c;
      38520: inst = 32'h8220000;
      38521: inst = 32'h10408000;
      38522: inst = 32'hc40514d;
      38523: inst = 32'h8220000;
      38524: inst = 32'h10408000;
      38525: inst = 32'hc40514e;
      38526: inst = 32'h8220000;
      38527: inst = 32'h10408000;
      38528: inst = 32'hc40514f;
      38529: inst = 32'h8220000;
      38530: inst = 32'h10408000;
      38531: inst = 32'hc405150;
      38532: inst = 32'h8220000;
      38533: inst = 32'h10408000;
      38534: inst = 32'hc405151;
      38535: inst = 32'h8220000;
      38536: inst = 32'h10408000;
      38537: inst = 32'hc405152;
      38538: inst = 32'h8220000;
      38539: inst = 32'h10408000;
      38540: inst = 32'hc405153;
      38541: inst = 32'h8220000;
      38542: inst = 32'h10408000;
      38543: inst = 32'hc405154;
      38544: inst = 32'h8220000;
      38545: inst = 32'h10408000;
      38546: inst = 32'hc405155;
      38547: inst = 32'h8220000;
      38548: inst = 32'h10408000;
      38549: inst = 32'hc405156;
      38550: inst = 32'h8220000;
      38551: inst = 32'h10408000;
      38552: inst = 32'hc405157;
      38553: inst = 32'h8220000;
      38554: inst = 32'h10408000;
      38555: inst = 32'hc405183;
      38556: inst = 32'h8220000;
      38557: inst = 32'h10408000;
      38558: inst = 32'hc405184;
      38559: inst = 32'h8220000;
      38560: inst = 32'h10408000;
      38561: inst = 32'hc405185;
      38562: inst = 32'h8220000;
      38563: inst = 32'h10408000;
      38564: inst = 32'hc405186;
      38565: inst = 32'h8220000;
      38566: inst = 32'h10408000;
      38567: inst = 32'hc405187;
      38568: inst = 32'h8220000;
      38569: inst = 32'h10408000;
      38570: inst = 32'hc405188;
      38571: inst = 32'h8220000;
      38572: inst = 32'h10408000;
      38573: inst = 32'hc405189;
      38574: inst = 32'h8220000;
      38575: inst = 32'h10408000;
      38576: inst = 32'hc40518a;
      38577: inst = 32'h8220000;
      38578: inst = 32'h10408000;
      38579: inst = 32'hc40518b;
      38580: inst = 32'h8220000;
      38581: inst = 32'h10408000;
      38582: inst = 32'hc40518c;
      38583: inst = 32'h8220000;
      38584: inst = 32'h10408000;
      38585: inst = 32'hc40518d;
      38586: inst = 32'h8220000;
      38587: inst = 32'h10408000;
      38588: inst = 32'hc40518e;
      38589: inst = 32'h8220000;
      38590: inst = 32'h10408000;
      38591: inst = 32'hc40518f;
      38592: inst = 32'h8220000;
      38593: inst = 32'h10408000;
      38594: inst = 32'hc405190;
      38595: inst = 32'h8220000;
      38596: inst = 32'h10408000;
      38597: inst = 32'hc405191;
      38598: inst = 32'h8220000;
      38599: inst = 32'h10408000;
      38600: inst = 32'hc405192;
      38601: inst = 32'h8220000;
      38602: inst = 32'h10408000;
      38603: inst = 32'hc405193;
      38604: inst = 32'h8220000;
      38605: inst = 32'h10408000;
      38606: inst = 32'hc405194;
      38607: inst = 32'h8220000;
      38608: inst = 32'h10408000;
      38609: inst = 32'hc405195;
      38610: inst = 32'h8220000;
      38611: inst = 32'h10408000;
      38612: inst = 32'hc405199;
      38613: inst = 32'h8220000;
      38614: inst = 32'h10408000;
      38615: inst = 32'hc40519a;
      38616: inst = 32'h8220000;
      38617: inst = 32'h10408000;
      38618: inst = 32'hc40519b;
      38619: inst = 32'h8220000;
      38620: inst = 32'h10408000;
      38621: inst = 32'hc40519c;
      38622: inst = 32'h8220000;
      38623: inst = 32'h10408000;
      38624: inst = 32'hc40519d;
      38625: inst = 32'h8220000;
      38626: inst = 32'h10408000;
      38627: inst = 32'hc40519e;
      38628: inst = 32'h8220000;
      38629: inst = 32'h10408000;
      38630: inst = 32'hc40519f;
      38631: inst = 32'h8220000;
      38632: inst = 32'h10408000;
      38633: inst = 32'hc4051a0;
      38634: inst = 32'h8220000;
      38635: inst = 32'h10408000;
      38636: inst = 32'hc4051a1;
      38637: inst = 32'h8220000;
      38638: inst = 32'h10408000;
      38639: inst = 32'hc4051a2;
      38640: inst = 32'h8220000;
      38641: inst = 32'h10408000;
      38642: inst = 32'hc4051a3;
      38643: inst = 32'h8220000;
      38644: inst = 32'h10408000;
      38645: inst = 32'hc4051a4;
      38646: inst = 32'h8220000;
      38647: inst = 32'h10408000;
      38648: inst = 32'hc4051a5;
      38649: inst = 32'h8220000;
      38650: inst = 32'h10408000;
      38651: inst = 32'hc4051a6;
      38652: inst = 32'h8220000;
      38653: inst = 32'h10408000;
      38654: inst = 32'hc4051a7;
      38655: inst = 32'h8220000;
      38656: inst = 32'h10408000;
      38657: inst = 32'hc4051a8;
      38658: inst = 32'h8220000;
      38659: inst = 32'h10408000;
      38660: inst = 32'hc4051a9;
      38661: inst = 32'h8220000;
      38662: inst = 32'h10408000;
      38663: inst = 32'hc4051aa;
      38664: inst = 32'h8220000;
      38665: inst = 32'h10408000;
      38666: inst = 32'hc4051ab;
      38667: inst = 32'h8220000;
      38668: inst = 32'h10408000;
      38669: inst = 32'hc4051ac;
      38670: inst = 32'h8220000;
      38671: inst = 32'h10408000;
      38672: inst = 32'hc4051ad;
      38673: inst = 32'h8220000;
      38674: inst = 32'h10408000;
      38675: inst = 32'hc4051ae;
      38676: inst = 32'h8220000;
      38677: inst = 32'h10408000;
      38678: inst = 32'hc4051af;
      38679: inst = 32'h8220000;
      38680: inst = 32'h10408000;
      38681: inst = 32'hc4051b0;
      38682: inst = 32'h8220000;
      38683: inst = 32'h10408000;
      38684: inst = 32'hc4051b1;
      38685: inst = 32'h8220000;
      38686: inst = 32'h10408000;
      38687: inst = 32'hc4051b2;
      38688: inst = 32'h8220000;
      38689: inst = 32'h10408000;
      38690: inst = 32'hc4051b3;
      38691: inst = 32'h8220000;
      38692: inst = 32'h10408000;
      38693: inst = 32'hc4051b4;
      38694: inst = 32'h8220000;
      38695: inst = 32'h10408000;
      38696: inst = 32'hc4051b5;
      38697: inst = 32'h8220000;
      38698: inst = 32'h10408000;
      38699: inst = 32'hc4051b6;
      38700: inst = 32'h8220000;
      38701: inst = 32'h10408000;
      38702: inst = 32'hc4051b7;
      38703: inst = 32'h8220000;
      38704: inst = 32'h10408000;
      38705: inst = 32'hc4051b8;
      38706: inst = 32'h8220000;
      38707: inst = 32'h10408000;
      38708: inst = 32'hc4051b9;
      38709: inst = 32'h8220000;
      38710: inst = 32'h10408000;
      38711: inst = 32'hc4051ba;
      38712: inst = 32'h8220000;
      38713: inst = 32'h10408000;
      38714: inst = 32'hc4051bb;
      38715: inst = 32'h8220000;
      38716: inst = 32'h10408000;
      38717: inst = 32'hc4051bc;
      38718: inst = 32'h8220000;
      38719: inst = 32'h10408000;
      38720: inst = 32'hc4051bd;
      38721: inst = 32'h8220000;
      38722: inst = 32'h10408000;
      38723: inst = 32'hc4051be;
      38724: inst = 32'h8220000;
      38725: inst = 32'h10408000;
      38726: inst = 32'hc4051bf;
      38727: inst = 32'h8220000;
      38728: inst = 32'h10408000;
      38729: inst = 32'hc4051c0;
      38730: inst = 32'h8220000;
      38731: inst = 32'h10408000;
      38732: inst = 32'hc4051c1;
      38733: inst = 32'h8220000;
      38734: inst = 32'h10408000;
      38735: inst = 32'hc4051c2;
      38736: inst = 32'h8220000;
      38737: inst = 32'h10408000;
      38738: inst = 32'hc4051c3;
      38739: inst = 32'h8220000;
      38740: inst = 32'h10408000;
      38741: inst = 32'hc4051c4;
      38742: inst = 32'h8220000;
      38743: inst = 32'h10408000;
      38744: inst = 32'hc4051c5;
      38745: inst = 32'h8220000;
      38746: inst = 32'h10408000;
      38747: inst = 32'hc4051c6;
      38748: inst = 32'h8220000;
      38749: inst = 32'h10408000;
      38750: inst = 32'hc4051c7;
      38751: inst = 32'h8220000;
      38752: inst = 32'h10408000;
      38753: inst = 32'hc4051c8;
      38754: inst = 32'h8220000;
      38755: inst = 32'h10408000;
      38756: inst = 32'hc4051c9;
      38757: inst = 32'h8220000;
      38758: inst = 32'h10408000;
      38759: inst = 32'hc4051ca;
      38760: inst = 32'h8220000;
      38761: inst = 32'h10408000;
      38762: inst = 32'hc4051cb;
      38763: inst = 32'h8220000;
      38764: inst = 32'h10408000;
      38765: inst = 32'hc4051cc;
      38766: inst = 32'h8220000;
      38767: inst = 32'h10408000;
      38768: inst = 32'hc4051cd;
      38769: inst = 32'h8220000;
      38770: inst = 32'h10408000;
      38771: inst = 32'hc4051ce;
      38772: inst = 32'h8220000;
      38773: inst = 32'h10408000;
      38774: inst = 32'hc4051cf;
      38775: inst = 32'h8220000;
      38776: inst = 32'h10408000;
      38777: inst = 32'hc4051d0;
      38778: inst = 32'h8220000;
      38779: inst = 32'h10408000;
      38780: inst = 32'hc4051d1;
      38781: inst = 32'h8220000;
      38782: inst = 32'h10408000;
      38783: inst = 32'hc4051d2;
      38784: inst = 32'h8220000;
      38785: inst = 32'h10408000;
      38786: inst = 32'hc4051d3;
      38787: inst = 32'h8220000;
      38788: inst = 32'h10408000;
      38789: inst = 32'hc4051d4;
      38790: inst = 32'h8220000;
      38791: inst = 32'h10408000;
      38792: inst = 32'hc4051d5;
      38793: inst = 32'h8220000;
      38794: inst = 32'h10408000;
      38795: inst = 32'hc4051d6;
      38796: inst = 32'h8220000;
      38797: inst = 32'h10408000;
      38798: inst = 32'hc4051d7;
      38799: inst = 32'h8220000;
      38800: inst = 32'h10408000;
      38801: inst = 32'hc4051d8;
      38802: inst = 32'h8220000;
      38803: inst = 32'h10408000;
      38804: inst = 32'hc4051d9;
      38805: inst = 32'h8220000;
      38806: inst = 32'h10408000;
      38807: inst = 32'hc4051da;
      38808: inst = 32'h8220000;
      38809: inst = 32'h10408000;
      38810: inst = 32'hc4051db;
      38811: inst = 32'h8220000;
      38812: inst = 32'h10408000;
      38813: inst = 32'hc4051dc;
      38814: inst = 32'h8220000;
      38815: inst = 32'h10408000;
      38816: inst = 32'hc4051e3;
      38817: inst = 32'h8220000;
      38818: inst = 32'h10408000;
      38819: inst = 32'hc4051e4;
      38820: inst = 32'h8220000;
      38821: inst = 32'h10408000;
      38822: inst = 32'hc4051e5;
      38823: inst = 32'h8220000;
      38824: inst = 32'h10408000;
      38825: inst = 32'hc4051e6;
      38826: inst = 32'h8220000;
      38827: inst = 32'h10408000;
      38828: inst = 32'hc4051e7;
      38829: inst = 32'h8220000;
      38830: inst = 32'h10408000;
      38831: inst = 32'hc4051e8;
      38832: inst = 32'h8220000;
      38833: inst = 32'h10408000;
      38834: inst = 32'hc4051e9;
      38835: inst = 32'h8220000;
      38836: inst = 32'h10408000;
      38837: inst = 32'hc4051ea;
      38838: inst = 32'h8220000;
      38839: inst = 32'h10408000;
      38840: inst = 32'hc4051eb;
      38841: inst = 32'h8220000;
      38842: inst = 32'h10408000;
      38843: inst = 32'hc4051ec;
      38844: inst = 32'h8220000;
      38845: inst = 32'h10408000;
      38846: inst = 32'hc4051ed;
      38847: inst = 32'h8220000;
      38848: inst = 32'h10408000;
      38849: inst = 32'hc4051ee;
      38850: inst = 32'h8220000;
      38851: inst = 32'h10408000;
      38852: inst = 32'hc4051ef;
      38853: inst = 32'h8220000;
      38854: inst = 32'h10408000;
      38855: inst = 32'hc4051f0;
      38856: inst = 32'h8220000;
      38857: inst = 32'h10408000;
      38858: inst = 32'hc4051f1;
      38859: inst = 32'h8220000;
      38860: inst = 32'h10408000;
      38861: inst = 32'hc4051f2;
      38862: inst = 32'h8220000;
      38863: inst = 32'h10408000;
      38864: inst = 32'hc4051f3;
      38865: inst = 32'h8220000;
      38866: inst = 32'h10408000;
      38867: inst = 32'hc4051f4;
      38868: inst = 32'h8220000;
      38869: inst = 32'h10408000;
      38870: inst = 32'hc4051f5;
      38871: inst = 32'h8220000;
      38872: inst = 32'h10408000;
      38873: inst = 32'hc4051f9;
      38874: inst = 32'h8220000;
      38875: inst = 32'h10408000;
      38876: inst = 32'hc4051fa;
      38877: inst = 32'h8220000;
      38878: inst = 32'h10408000;
      38879: inst = 32'hc4051fb;
      38880: inst = 32'h8220000;
      38881: inst = 32'h10408000;
      38882: inst = 32'hc4051fc;
      38883: inst = 32'h8220000;
      38884: inst = 32'h10408000;
      38885: inst = 32'hc4051fd;
      38886: inst = 32'h8220000;
      38887: inst = 32'h10408000;
      38888: inst = 32'hc4051fe;
      38889: inst = 32'h8220000;
      38890: inst = 32'h10408000;
      38891: inst = 32'hc4051ff;
      38892: inst = 32'h8220000;
      38893: inst = 32'h10408000;
      38894: inst = 32'hc405200;
      38895: inst = 32'h8220000;
      38896: inst = 32'h10408000;
      38897: inst = 32'hc405201;
      38898: inst = 32'h8220000;
      38899: inst = 32'h10408000;
      38900: inst = 32'hc405202;
      38901: inst = 32'h8220000;
      38902: inst = 32'h10408000;
      38903: inst = 32'hc405203;
      38904: inst = 32'h8220000;
      38905: inst = 32'h10408000;
      38906: inst = 32'hc405204;
      38907: inst = 32'h8220000;
      38908: inst = 32'h10408000;
      38909: inst = 32'hc405205;
      38910: inst = 32'h8220000;
      38911: inst = 32'h10408000;
      38912: inst = 32'hc405206;
      38913: inst = 32'h8220000;
      38914: inst = 32'h10408000;
      38915: inst = 32'hc405207;
      38916: inst = 32'h8220000;
      38917: inst = 32'h10408000;
      38918: inst = 32'hc405208;
      38919: inst = 32'h8220000;
      38920: inst = 32'h10408000;
      38921: inst = 32'hc405209;
      38922: inst = 32'h8220000;
      38923: inst = 32'h10408000;
      38924: inst = 32'hc40520a;
      38925: inst = 32'h8220000;
      38926: inst = 32'h10408000;
      38927: inst = 32'hc40520b;
      38928: inst = 32'h8220000;
      38929: inst = 32'h10408000;
      38930: inst = 32'hc40520c;
      38931: inst = 32'h8220000;
      38932: inst = 32'h10408000;
      38933: inst = 32'hc40520d;
      38934: inst = 32'h8220000;
      38935: inst = 32'h10408000;
      38936: inst = 32'hc40520e;
      38937: inst = 32'h8220000;
      38938: inst = 32'h10408000;
      38939: inst = 32'hc40520f;
      38940: inst = 32'h8220000;
      38941: inst = 32'h10408000;
      38942: inst = 32'hc405210;
      38943: inst = 32'h8220000;
      38944: inst = 32'h10408000;
      38945: inst = 32'hc405211;
      38946: inst = 32'h8220000;
      38947: inst = 32'h10408000;
      38948: inst = 32'hc405212;
      38949: inst = 32'h8220000;
      38950: inst = 32'h10408000;
      38951: inst = 32'hc405213;
      38952: inst = 32'h8220000;
      38953: inst = 32'h10408000;
      38954: inst = 32'hc405214;
      38955: inst = 32'h8220000;
      38956: inst = 32'h10408000;
      38957: inst = 32'hc405215;
      38958: inst = 32'h8220000;
      38959: inst = 32'h10408000;
      38960: inst = 32'hc405216;
      38961: inst = 32'h8220000;
      38962: inst = 32'h10408000;
      38963: inst = 32'hc405217;
      38964: inst = 32'h8220000;
      38965: inst = 32'h10408000;
      38966: inst = 32'hc405218;
      38967: inst = 32'h8220000;
      38968: inst = 32'h10408000;
      38969: inst = 32'hc405219;
      38970: inst = 32'h8220000;
      38971: inst = 32'h10408000;
      38972: inst = 32'hc40521a;
      38973: inst = 32'h8220000;
      38974: inst = 32'h10408000;
      38975: inst = 32'hc40521b;
      38976: inst = 32'h8220000;
      38977: inst = 32'h10408000;
      38978: inst = 32'hc40521c;
      38979: inst = 32'h8220000;
      38980: inst = 32'h10408000;
      38981: inst = 32'hc40521d;
      38982: inst = 32'h8220000;
      38983: inst = 32'h10408000;
      38984: inst = 32'hc40521e;
      38985: inst = 32'h8220000;
      38986: inst = 32'h10408000;
      38987: inst = 32'hc40521f;
      38988: inst = 32'h8220000;
      38989: inst = 32'h10408000;
      38990: inst = 32'hc405220;
      38991: inst = 32'h8220000;
      38992: inst = 32'h10408000;
      38993: inst = 32'hc405221;
      38994: inst = 32'h8220000;
      38995: inst = 32'h10408000;
      38996: inst = 32'hc405222;
      38997: inst = 32'h8220000;
      38998: inst = 32'h10408000;
      38999: inst = 32'hc405223;
      39000: inst = 32'h8220000;
      39001: inst = 32'h10408000;
      39002: inst = 32'hc405224;
      39003: inst = 32'h8220000;
      39004: inst = 32'h10408000;
      39005: inst = 32'hc405225;
      39006: inst = 32'h8220000;
      39007: inst = 32'h10408000;
      39008: inst = 32'hc405226;
      39009: inst = 32'h8220000;
      39010: inst = 32'h10408000;
      39011: inst = 32'hc405227;
      39012: inst = 32'h8220000;
      39013: inst = 32'h10408000;
      39014: inst = 32'hc405228;
      39015: inst = 32'h8220000;
      39016: inst = 32'h10408000;
      39017: inst = 32'hc405229;
      39018: inst = 32'h8220000;
      39019: inst = 32'h10408000;
      39020: inst = 32'hc40522a;
      39021: inst = 32'h8220000;
      39022: inst = 32'h10408000;
      39023: inst = 32'hc40522b;
      39024: inst = 32'h8220000;
      39025: inst = 32'h10408000;
      39026: inst = 32'hc40522c;
      39027: inst = 32'h8220000;
      39028: inst = 32'h10408000;
      39029: inst = 32'hc40522d;
      39030: inst = 32'h8220000;
      39031: inst = 32'h10408000;
      39032: inst = 32'hc40522e;
      39033: inst = 32'h8220000;
      39034: inst = 32'h10408000;
      39035: inst = 32'hc40522f;
      39036: inst = 32'h8220000;
      39037: inst = 32'h10408000;
      39038: inst = 32'hc405230;
      39039: inst = 32'h8220000;
      39040: inst = 32'h10408000;
      39041: inst = 32'hc405231;
      39042: inst = 32'h8220000;
      39043: inst = 32'h10408000;
      39044: inst = 32'hc405232;
      39045: inst = 32'h8220000;
      39046: inst = 32'h10408000;
      39047: inst = 32'hc405233;
      39048: inst = 32'h8220000;
      39049: inst = 32'h10408000;
      39050: inst = 32'hc405234;
      39051: inst = 32'h8220000;
      39052: inst = 32'h10408000;
      39053: inst = 32'hc405235;
      39054: inst = 32'h8220000;
      39055: inst = 32'h10408000;
      39056: inst = 32'hc405236;
      39057: inst = 32'h8220000;
      39058: inst = 32'h10408000;
      39059: inst = 32'hc405237;
      39060: inst = 32'h8220000;
      39061: inst = 32'h10408000;
      39062: inst = 32'hc405238;
      39063: inst = 32'h8220000;
      39064: inst = 32'h10408000;
      39065: inst = 32'hc405239;
      39066: inst = 32'h8220000;
      39067: inst = 32'h10408000;
      39068: inst = 32'hc40523a;
      39069: inst = 32'h8220000;
      39070: inst = 32'h10408000;
      39071: inst = 32'hc40523b;
      39072: inst = 32'h8220000;
      39073: inst = 32'h10408000;
      39074: inst = 32'hc40523c;
      39075: inst = 32'h8220000;
      39076: inst = 32'h10408000;
      39077: inst = 32'hc405243;
      39078: inst = 32'h8220000;
      39079: inst = 32'h10408000;
      39080: inst = 32'hc405244;
      39081: inst = 32'h8220000;
      39082: inst = 32'h10408000;
      39083: inst = 32'hc405245;
      39084: inst = 32'h8220000;
      39085: inst = 32'h10408000;
      39086: inst = 32'hc405246;
      39087: inst = 32'h8220000;
      39088: inst = 32'h10408000;
      39089: inst = 32'hc405247;
      39090: inst = 32'h8220000;
      39091: inst = 32'h10408000;
      39092: inst = 32'hc405248;
      39093: inst = 32'h8220000;
      39094: inst = 32'h10408000;
      39095: inst = 32'hc405249;
      39096: inst = 32'h8220000;
      39097: inst = 32'h10408000;
      39098: inst = 32'hc40524a;
      39099: inst = 32'h8220000;
      39100: inst = 32'h10408000;
      39101: inst = 32'hc40524b;
      39102: inst = 32'h8220000;
      39103: inst = 32'h10408000;
      39104: inst = 32'hc40524c;
      39105: inst = 32'h8220000;
      39106: inst = 32'h10408000;
      39107: inst = 32'hc40524d;
      39108: inst = 32'h8220000;
      39109: inst = 32'h10408000;
      39110: inst = 32'hc40524e;
      39111: inst = 32'h8220000;
      39112: inst = 32'h10408000;
      39113: inst = 32'hc40524f;
      39114: inst = 32'h8220000;
      39115: inst = 32'h10408000;
      39116: inst = 32'hc405250;
      39117: inst = 32'h8220000;
      39118: inst = 32'h10408000;
      39119: inst = 32'hc405251;
      39120: inst = 32'h8220000;
      39121: inst = 32'h10408000;
      39122: inst = 32'hc405252;
      39123: inst = 32'h8220000;
      39124: inst = 32'h10408000;
      39125: inst = 32'hc405253;
      39126: inst = 32'h8220000;
      39127: inst = 32'h10408000;
      39128: inst = 32'hc405254;
      39129: inst = 32'h8220000;
      39130: inst = 32'h10408000;
      39131: inst = 32'hc405255;
      39132: inst = 32'h8220000;
      39133: inst = 32'h10408000;
      39134: inst = 32'hc405259;
      39135: inst = 32'h8220000;
      39136: inst = 32'h10408000;
      39137: inst = 32'hc40525a;
      39138: inst = 32'h8220000;
      39139: inst = 32'h10408000;
      39140: inst = 32'hc40525b;
      39141: inst = 32'h8220000;
      39142: inst = 32'h10408000;
      39143: inst = 32'hc40525c;
      39144: inst = 32'h8220000;
      39145: inst = 32'h10408000;
      39146: inst = 32'hc40525d;
      39147: inst = 32'h8220000;
      39148: inst = 32'h10408000;
      39149: inst = 32'hc40525e;
      39150: inst = 32'h8220000;
      39151: inst = 32'h10408000;
      39152: inst = 32'hc40525f;
      39153: inst = 32'h8220000;
      39154: inst = 32'h10408000;
      39155: inst = 32'hc405260;
      39156: inst = 32'h8220000;
      39157: inst = 32'h10408000;
      39158: inst = 32'hc405261;
      39159: inst = 32'h8220000;
      39160: inst = 32'h10408000;
      39161: inst = 32'hc405262;
      39162: inst = 32'h8220000;
      39163: inst = 32'h10408000;
      39164: inst = 32'hc405263;
      39165: inst = 32'h8220000;
      39166: inst = 32'h10408000;
      39167: inst = 32'hc405264;
      39168: inst = 32'h8220000;
      39169: inst = 32'h10408000;
      39170: inst = 32'hc405265;
      39171: inst = 32'h8220000;
      39172: inst = 32'h10408000;
      39173: inst = 32'hc405266;
      39174: inst = 32'h8220000;
      39175: inst = 32'h10408000;
      39176: inst = 32'hc405267;
      39177: inst = 32'h8220000;
      39178: inst = 32'h10408000;
      39179: inst = 32'hc405268;
      39180: inst = 32'h8220000;
      39181: inst = 32'h10408000;
      39182: inst = 32'hc405269;
      39183: inst = 32'h8220000;
      39184: inst = 32'h10408000;
      39185: inst = 32'hc40526a;
      39186: inst = 32'h8220000;
      39187: inst = 32'h10408000;
      39188: inst = 32'hc40526b;
      39189: inst = 32'h8220000;
      39190: inst = 32'h10408000;
      39191: inst = 32'hc40526c;
      39192: inst = 32'h8220000;
      39193: inst = 32'h10408000;
      39194: inst = 32'hc40526d;
      39195: inst = 32'h8220000;
      39196: inst = 32'h10408000;
      39197: inst = 32'hc40526e;
      39198: inst = 32'h8220000;
      39199: inst = 32'h10408000;
      39200: inst = 32'hc40526f;
      39201: inst = 32'h8220000;
      39202: inst = 32'h10408000;
      39203: inst = 32'hc405270;
      39204: inst = 32'h8220000;
      39205: inst = 32'h10408000;
      39206: inst = 32'hc405271;
      39207: inst = 32'h8220000;
      39208: inst = 32'h10408000;
      39209: inst = 32'hc405272;
      39210: inst = 32'h8220000;
      39211: inst = 32'h10408000;
      39212: inst = 32'hc405273;
      39213: inst = 32'h8220000;
      39214: inst = 32'h10408000;
      39215: inst = 32'hc405274;
      39216: inst = 32'h8220000;
      39217: inst = 32'h10408000;
      39218: inst = 32'hc405275;
      39219: inst = 32'h8220000;
      39220: inst = 32'h10408000;
      39221: inst = 32'hc405276;
      39222: inst = 32'h8220000;
      39223: inst = 32'h10408000;
      39224: inst = 32'hc405277;
      39225: inst = 32'h8220000;
      39226: inst = 32'h10408000;
      39227: inst = 32'hc405278;
      39228: inst = 32'h8220000;
      39229: inst = 32'h10408000;
      39230: inst = 32'hc405279;
      39231: inst = 32'h8220000;
      39232: inst = 32'h10408000;
      39233: inst = 32'hc40527a;
      39234: inst = 32'h8220000;
      39235: inst = 32'h10408000;
      39236: inst = 32'hc40527b;
      39237: inst = 32'h8220000;
      39238: inst = 32'h10408000;
      39239: inst = 32'hc40527c;
      39240: inst = 32'h8220000;
      39241: inst = 32'h10408000;
      39242: inst = 32'hc40527d;
      39243: inst = 32'h8220000;
      39244: inst = 32'h10408000;
      39245: inst = 32'hc40527e;
      39246: inst = 32'h8220000;
      39247: inst = 32'h10408000;
      39248: inst = 32'hc40527f;
      39249: inst = 32'h8220000;
      39250: inst = 32'h10408000;
      39251: inst = 32'hc405280;
      39252: inst = 32'h8220000;
      39253: inst = 32'h10408000;
      39254: inst = 32'hc405281;
      39255: inst = 32'h8220000;
      39256: inst = 32'h10408000;
      39257: inst = 32'hc405282;
      39258: inst = 32'h8220000;
      39259: inst = 32'h10408000;
      39260: inst = 32'hc405283;
      39261: inst = 32'h8220000;
      39262: inst = 32'h10408000;
      39263: inst = 32'hc405284;
      39264: inst = 32'h8220000;
      39265: inst = 32'h10408000;
      39266: inst = 32'hc405285;
      39267: inst = 32'h8220000;
      39268: inst = 32'h10408000;
      39269: inst = 32'hc405286;
      39270: inst = 32'h8220000;
      39271: inst = 32'h10408000;
      39272: inst = 32'hc405287;
      39273: inst = 32'h8220000;
      39274: inst = 32'h10408000;
      39275: inst = 32'hc405288;
      39276: inst = 32'h8220000;
      39277: inst = 32'h10408000;
      39278: inst = 32'hc405289;
      39279: inst = 32'h8220000;
      39280: inst = 32'h10408000;
      39281: inst = 32'hc40528a;
      39282: inst = 32'h8220000;
      39283: inst = 32'h10408000;
      39284: inst = 32'hc40528b;
      39285: inst = 32'h8220000;
      39286: inst = 32'h10408000;
      39287: inst = 32'hc40528c;
      39288: inst = 32'h8220000;
      39289: inst = 32'h10408000;
      39290: inst = 32'hc40528d;
      39291: inst = 32'h8220000;
      39292: inst = 32'h10408000;
      39293: inst = 32'hc40528e;
      39294: inst = 32'h8220000;
      39295: inst = 32'h10408000;
      39296: inst = 32'hc40528f;
      39297: inst = 32'h8220000;
      39298: inst = 32'h10408000;
      39299: inst = 32'hc405290;
      39300: inst = 32'h8220000;
      39301: inst = 32'h10408000;
      39302: inst = 32'hc405291;
      39303: inst = 32'h8220000;
      39304: inst = 32'h10408000;
      39305: inst = 32'hc405292;
      39306: inst = 32'h8220000;
      39307: inst = 32'h10408000;
      39308: inst = 32'hc405293;
      39309: inst = 32'h8220000;
      39310: inst = 32'h10408000;
      39311: inst = 32'hc405294;
      39312: inst = 32'h8220000;
      39313: inst = 32'h10408000;
      39314: inst = 32'hc405295;
      39315: inst = 32'h8220000;
      39316: inst = 32'h10408000;
      39317: inst = 32'hc405296;
      39318: inst = 32'h8220000;
      39319: inst = 32'h10408000;
      39320: inst = 32'hc405297;
      39321: inst = 32'h8220000;
      39322: inst = 32'h10408000;
      39323: inst = 32'hc405298;
      39324: inst = 32'h8220000;
      39325: inst = 32'h10408000;
      39326: inst = 32'hc405299;
      39327: inst = 32'h8220000;
      39328: inst = 32'h10408000;
      39329: inst = 32'hc40529a;
      39330: inst = 32'h8220000;
      39331: inst = 32'h10408000;
      39332: inst = 32'hc40529b;
      39333: inst = 32'h8220000;
      39334: inst = 32'h10408000;
      39335: inst = 32'hc40529c;
      39336: inst = 32'h8220000;
      39337: inst = 32'h10408000;
      39338: inst = 32'hc4052a3;
      39339: inst = 32'h8220000;
      39340: inst = 32'h10408000;
      39341: inst = 32'hc4052a4;
      39342: inst = 32'h8220000;
      39343: inst = 32'h10408000;
      39344: inst = 32'hc4052a5;
      39345: inst = 32'h8220000;
      39346: inst = 32'h10408000;
      39347: inst = 32'hc4052a6;
      39348: inst = 32'h8220000;
      39349: inst = 32'h10408000;
      39350: inst = 32'hc4052a7;
      39351: inst = 32'h8220000;
      39352: inst = 32'h10408000;
      39353: inst = 32'hc4052a8;
      39354: inst = 32'h8220000;
      39355: inst = 32'h10408000;
      39356: inst = 32'hc4052a9;
      39357: inst = 32'h8220000;
      39358: inst = 32'h10408000;
      39359: inst = 32'hc4052aa;
      39360: inst = 32'h8220000;
      39361: inst = 32'h10408000;
      39362: inst = 32'hc4052ab;
      39363: inst = 32'h8220000;
      39364: inst = 32'h10408000;
      39365: inst = 32'hc4052ac;
      39366: inst = 32'h8220000;
      39367: inst = 32'h10408000;
      39368: inst = 32'hc4052ad;
      39369: inst = 32'h8220000;
      39370: inst = 32'h10408000;
      39371: inst = 32'hc4052ae;
      39372: inst = 32'h8220000;
      39373: inst = 32'h10408000;
      39374: inst = 32'hc4052af;
      39375: inst = 32'h8220000;
      39376: inst = 32'h10408000;
      39377: inst = 32'hc4052b0;
      39378: inst = 32'h8220000;
      39379: inst = 32'h10408000;
      39380: inst = 32'hc4052b1;
      39381: inst = 32'h8220000;
      39382: inst = 32'h10408000;
      39383: inst = 32'hc4052b2;
      39384: inst = 32'h8220000;
      39385: inst = 32'h10408000;
      39386: inst = 32'hc4052b3;
      39387: inst = 32'h8220000;
      39388: inst = 32'h10408000;
      39389: inst = 32'hc4052b4;
      39390: inst = 32'h8220000;
      39391: inst = 32'h10408000;
      39392: inst = 32'hc4052b5;
      39393: inst = 32'h8220000;
      39394: inst = 32'h10408000;
      39395: inst = 32'hc4052b9;
      39396: inst = 32'h8220000;
      39397: inst = 32'h10408000;
      39398: inst = 32'hc4052ba;
      39399: inst = 32'h8220000;
      39400: inst = 32'h10408000;
      39401: inst = 32'hc4052bb;
      39402: inst = 32'h8220000;
      39403: inst = 32'h10408000;
      39404: inst = 32'hc4052bc;
      39405: inst = 32'h8220000;
      39406: inst = 32'h10408000;
      39407: inst = 32'hc4052bd;
      39408: inst = 32'h8220000;
      39409: inst = 32'h10408000;
      39410: inst = 32'hc4052be;
      39411: inst = 32'h8220000;
      39412: inst = 32'h10408000;
      39413: inst = 32'hc4052bf;
      39414: inst = 32'h8220000;
      39415: inst = 32'h10408000;
      39416: inst = 32'hc4052c0;
      39417: inst = 32'h8220000;
      39418: inst = 32'h10408000;
      39419: inst = 32'hc4052c1;
      39420: inst = 32'h8220000;
      39421: inst = 32'h10408000;
      39422: inst = 32'hc4052c2;
      39423: inst = 32'h8220000;
      39424: inst = 32'h10408000;
      39425: inst = 32'hc4052c3;
      39426: inst = 32'h8220000;
      39427: inst = 32'h10408000;
      39428: inst = 32'hc4052c4;
      39429: inst = 32'h8220000;
      39430: inst = 32'h10408000;
      39431: inst = 32'hc4052c5;
      39432: inst = 32'h8220000;
      39433: inst = 32'h10408000;
      39434: inst = 32'hc4052c6;
      39435: inst = 32'h8220000;
      39436: inst = 32'h10408000;
      39437: inst = 32'hc4052c7;
      39438: inst = 32'h8220000;
      39439: inst = 32'h10408000;
      39440: inst = 32'hc4052c8;
      39441: inst = 32'h8220000;
      39442: inst = 32'h10408000;
      39443: inst = 32'hc4052c9;
      39444: inst = 32'h8220000;
      39445: inst = 32'h10408000;
      39446: inst = 32'hc4052ca;
      39447: inst = 32'h8220000;
      39448: inst = 32'h10408000;
      39449: inst = 32'hc4052cb;
      39450: inst = 32'h8220000;
      39451: inst = 32'h10408000;
      39452: inst = 32'hc4052cc;
      39453: inst = 32'h8220000;
      39454: inst = 32'h10408000;
      39455: inst = 32'hc4052cd;
      39456: inst = 32'h8220000;
      39457: inst = 32'h10408000;
      39458: inst = 32'hc4052ce;
      39459: inst = 32'h8220000;
      39460: inst = 32'h10408000;
      39461: inst = 32'hc4052cf;
      39462: inst = 32'h8220000;
      39463: inst = 32'h10408000;
      39464: inst = 32'hc4052d0;
      39465: inst = 32'h8220000;
      39466: inst = 32'h10408000;
      39467: inst = 32'hc4052d1;
      39468: inst = 32'h8220000;
      39469: inst = 32'h10408000;
      39470: inst = 32'hc4052d2;
      39471: inst = 32'h8220000;
      39472: inst = 32'h10408000;
      39473: inst = 32'hc4052d3;
      39474: inst = 32'h8220000;
      39475: inst = 32'h10408000;
      39476: inst = 32'hc4052d4;
      39477: inst = 32'h8220000;
      39478: inst = 32'h10408000;
      39479: inst = 32'hc4052d5;
      39480: inst = 32'h8220000;
      39481: inst = 32'h10408000;
      39482: inst = 32'hc4052d6;
      39483: inst = 32'h8220000;
      39484: inst = 32'h10408000;
      39485: inst = 32'hc4052d7;
      39486: inst = 32'h8220000;
      39487: inst = 32'h10408000;
      39488: inst = 32'hc4052d8;
      39489: inst = 32'h8220000;
      39490: inst = 32'h10408000;
      39491: inst = 32'hc4052d9;
      39492: inst = 32'h8220000;
      39493: inst = 32'h10408000;
      39494: inst = 32'hc4052da;
      39495: inst = 32'h8220000;
      39496: inst = 32'h10408000;
      39497: inst = 32'hc4052db;
      39498: inst = 32'h8220000;
      39499: inst = 32'h10408000;
      39500: inst = 32'hc4052dc;
      39501: inst = 32'h8220000;
      39502: inst = 32'h10408000;
      39503: inst = 32'hc4052dd;
      39504: inst = 32'h8220000;
      39505: inst = 32'h10408000;
      39506: inst = 32'hc4052de;
      39507: inst = 32'h8220000;
      39508: inst = 32'h10408000;
      39509: inst = 32'hc4052df;
      39510: inst = 32'h8220000;
      39511: inst = 32'h10408000;
      39512: inst = 32'hc4052e0;
      39513: inst = 32'h8220000;
      39514: inst = 32'h10408000;
      39515: inst = 32'hc4052e1;
      39516: inst = 32'h8220000;
      39517: inst = 32'h10408000;
      39518: inst = 32'hc4052e2;
      39519: inst = 32'h8220000;
      39520: inst = 32'h10408000;
      39521: inst = 32'hc4052e3;
      39522: inst = 32'h8220000;
      39523: inst = 32'h10408000;
      39524: inst = 32'hc4052e4;
      39525: inst = 32'h8220000;
      39526: inst = 32'h10408000;
      39527: inst = 32'hc4052e5;
      39528: inst = 32'h8220000;
      39529: inst = 32'h10408000;
      39530: inst = 32'hc4052e6;
      39531: inst = 32'h8220000;
      39532: inst = 32'h10408000;
      39533: inst = 32'hc4052e7;
      39534: inst = 32'h8220000;
      39535: inst = 32'h10408000;
      39536: inst = 32'hc4052e8;
      39537: inst = 32'h8220000;
      39538: inst = 32'h10408000;
      39539: inst = 32'hc4052e9;
      39540: inst = 32'h8220000;
      39541: inst = 32'h10408000;
      39542: inst = 32'hc4052ea;
      39543: inst = 32'h8220000;
      39544: inst = 32'h10408000;
      39545: inst = 32'hc4052eb;
      39546: inst = 32'h8220000;
      39547: inst = 32'h10408000;
      39548: inst = 32'hc4052ec;
      39549: inst = 32'h8220000;
      39550: inst = 32'h10408000;
      39551: inst = 32'hc4052ed;
      39552: inst = 32'h8220000;
      39553: inst = 32'h10408000;
      39554: inst = 32'hc4052ee;
      39555: inst = 32'h8220000;
      39556: inst = 32'h10408000;
      39557: inst = 32'hc4052ef;
      39558: inst = 32'h8220000;
      39559: inst = 32'h10408000;
      39560: inst = 32'hc4052f0;
      39561: inst = 32'h8220000;
      39562: inst = 32'h10408000;
      39563: inst = 32'hc4052f1;
      39564: inst = 32'h8220000;
      39565: inst = 32'h10408000;
      39566: inst = 32'hc4052f2;
      39567: inst = 32'h8220000;
      39568: inst = 32'h10408000;
      39569: inst = 32'hc4052f3;
      39570: inst = 32'h8220000;
      39571: inst = 32'h10408000;
      39572: inst = 32'hc4052f4;
      39573: inst = 32'h8220000;
      39574: inst = 32'h10408000;
      39575: inst = 32'hc4052f5;
      39576: inst = 32'h8220000;
      39577: inst = 32'h10408000;
      39578: inst = 32'hc4052f6;
      39579: inst = 32'h8220000;
      39580: inst = 32'h10408000;
      39581: inst = 32'hc4052f7;
      39582: inst = 32'h8220000;
      39583: inst = 32'h10408000;
      39584: inst = 32'hc4052f8;
      39585: inst = 32'h8220000;
      39586: inst = 32'h10408000;
      39587: inst = 32'hc4052f9;
      39588: inst = 32'h8220000;
      39589: inst = 32'h10408000;
      39590: inst = 32'hc4052fa;
      39591: inst = 32'h8220000;
      39592: inst = 32'h10408000;
      39593: inst = 32'hc4052fb;
      39594: inst = 32'h8220000;
      39595: inst = 32'h10408000;
      39596: inst = 32'hc4052fc;
      39597: inst = 32'h8220000;
      39598: inst = 32'h10408000;
      39599: inst = 32'hc405303;
      39600: inst = 32'h8220000;
      39601: inst = 32'h10408000;
      39602: inst = 32'hc405304;
      39603: inst = 32'h8220000;
      39604: inst = 32'h10408000;
      39605: inst = 32'hc405305;
      39606: inst = 32'h8220000;
      39607: inst = 32'h10408000;
      39608: inst = 32'hc405306;
      39609: inst = 32'h8220000;
      39610: inst = 32'h10408000;
      39611: inst = 32'hc405307;
      39612: inst = 32'h8220000;
      39613: inst = 32'h10408000;
      39614: inst = 32'hc405308;
      39615: inst = 32'h8220000;
      39616: inst = 32'h10408000;
      39617: inst = 32'hc405309;
      39618: inst = 32'h8220000;
      39619: inst = 32'h10408000;
      39620: inst = 32'hc40530a;
      39621: inst = 32'h8220000;
      39622: inst = 32'h10408000;
      39623: inst = 32'hc40530b;
      39624: inst = 32'h8220000;
      39625: inst = 32'h10408000;
      39626: inst = 32'hc40530c;
      39627: inst = 32'h8220000;
      39628: inst = 32'h10408000;
      39629: inst = 32'hc40530d;
      39630: inst = 32'h8220000;
      39631: inst = 32'h10408000;
      39632: inst = 32'hc40530e;
      39633: inst = 32'h8220000;
      39634: inst = 32'h10408000;
      39635: inst = 32'hc40530f;
      39636: inst = 32'h8220000;
      39637: inst = 32'h10408000;
      39638: inst = 32'hc405310;
      39639: inst = 32'h8220000;
      39640: inst = 32'h10408000;
      39641: inst = 32'hc405311;
      39642: inst = 32'h8220000;
      39643: inst = 32'h10408000;
      39644: inst = 32'hc405312;
      39645: inst = 32'h8220000;
      39646: inst = 32'h10408000;
      39647: inst = 32'hc405313;
      39648: inst = 32'h8220000;
      39649: inst = 32'h10408000;
      39650: inst = 32'hc405314;
      39651: inst = 32'h8220000;
      39652: inst = 32'h10408000;
      39653: inst = 32'hc405315;
      39654: inst = 32'h8220000;
      39655: inst = 32'h10408000;
      39656: inst = 32'hc405319;
      39657: inst = 32'h8220000;
      39658: inst = 32'h10408000;
      39659: inst = 32'hc40531a;
      39660: inst = 32'h8220000;
      39661: inst = 32'h10408000;
      39662: inst = 32'hc40531b;
      39663: inst = 32'h8220000;
      39664: inst = 32'h10408000;
      39665: inst = 32'hc40531c;
      39666: inst = 32'h8220000;
      39667: inst = 32'h10408000;
      39668: inst = 32'hc40531d;
      39669: inst = 32'h8220000;
      39670: inst = 32'h10408000;
      39671: inst = 32'hc40531e;
      39672: inst = 32'h8220000;
      39673: inst = 32'h10408000;
      39674: inst = 32'hc40531f;
      39675: inst = 32'h8220000;
      39676: inst = 32'h10408000;
      39677: inst = 32'hc405320;
      39678: inst = 32'h8220000;
      39679: inst = 32'h10408000;
      39680: inst = 32'hc405321;
      39681: inst = 32'h8220000;
      39682: inst = 32'h10408000;
      39683: inst = 32'hc405322;
      39684: inst = 32'h8220000;
      39685: inst = 32'h10408000;
      39686: inst = 32'hc405323;
      39687: inst = 32'h8220000;
      39688: inst = 32'h10408000;
      39689: inst = 32'hc405324;
      39690: inst = 32'h8220000;
      39691: inst = 32'h10408000;
      39692: inst = 32'hc405325;
      39693: inst = 32'h8220000;
      39694: inst = 32'h10408000;
      39695: inst = 32'hc405326;
      39696: inst = 32'h8220000;
      39697: inst = 32'h10408000;
      39698: inst = 32'hc405327;
      39699: inst = 32'h8220000;
      39700: inst = 32'h10408000;
      39701: inst = 32'hc405328;
      39702: inst = 32'h8220000;
      39703: inst = 32'h10408000;
      39704: inst = 32'hc405329;
      39705: inst = 32'h8220000;
      39706: inst = 32'h10408000;
      39707: inst = 32'hc40532a;
      39708: inst = 32'h8220000;
      39709: inst = 32'h10408000;
      39710: inst = 32'hc40532b;
      39711: inst = 32'h8220000;
      39712: inst = 32'h10408000;
      39713: inst = 32'hc40532c;
      39714: inst = 32'h8220000;
      39715: inst = 32'h10408000;
      39716: inst = 32'hc40532d;
      39717: inst = 32'h8220000;
      39718: inst = 32'h10408000;
      39719: inst = 32'hc40532e;
      39720: inst = 32'h8220000;
      39721: inst = 32'h10408000;
      39722: inst = 32'hc40532f;
      39723: inst = 32'h8220000;
      39724: inst = 32'h10408000;
      39725: inst = 32'hc405330;
      39726: inst = 32'h8220000;
      39727: inst = 32'h10408000;
      39728: inst = 32'hc405331;
      39729: inst = 32'h8220000;
      39730: inst = 32'h10408000;
      39731: inst = 32'hc405332;
      39732: inst = 32'h8220000;
      39733: inst = 32'h10408000;
      39734: inst = 32'hc405333;
      39735: inst = 32'h8220000;
      39736: inst = 32'h10408000;
      39737: inst = 32'hc405334;
      39738: inst = 32'h8220000;
      39739: inst = 32'h10408000;
      39740: inst = 32'hc405335;
      39741: inst = 32'h8220000;
      39742: inst = 32'h10408000;
      39743: inst = 32'hc405336;
      39744: inst = 32'h8220000;
      39745: inst = 32'h10408000;
      39746: inst = 32'hc405337;
      39747: inst = 32'h8220000;
      39748: inst = 32'h10408000;
      39749: inst = 32'hc405338;
      39750: inst = 32'h8220000;
      39751: inst = 32'h10408000;
      39752: inst = 32'hc405339;
      39753: inst = 32'h8220000;
      39754: inst = 32'h10408000;
      39755: inst = 32'hc40533a;
      39756: inst = 32'h8220000;
      39757: inst = 32'h10408000;
      39758: inst = 32'hc40533b;
      39759: inst = 32'h8220000;
      39760: inst = 32'h10408000;
      39761: inst = 32'hc40533c;
      39762: inst = 32'h8220000;
      39763: inst = 32'h10408000;
      39764: inst = 32'hc40533d;
      39765: inst = 32'h8220000;
      39766: inst = 32'h10408000;
      39767: inst = 32'hc40533e;
      39768: inst = 32'h8220000;
      39769: inst = 32'h10408000;
      39770: inst = 32'hc40533f;
      39771: inst = 32'h8220000;
      39772: inst = 32'h10408000;
      39773: inst = 32'hc405340;
      39774: inst = 32'h8220000;
      39775: inst = 32'h10408000;
      39776: inst = 32'hc405341;
      39777: inst = 32'h8220000;
      39778: inst = 32'h10408000;
      39779: inst = 32'hc405342;
      39780: inst = 32'h8220000;
      39781: inst = 32'h10408000;
      39782: inst = 32'hc405343;
      39783: inst = 32'h8220000;
      39784: inst = 32'h10408000;
      39785: inst = 32'hc405344;
      39786: inst = 32'h8220000;
      39787: inst = 32'h10408000;
      39788: inst = 32'hc405345;
      39789: inst = 32'h8220000;
      39790: inst = 32'h10408000;
      39791: inst = 32'hc405346;
      39792: inst = 32'h8220000;
      39793: inst = 32'h10408000;
      39794: inst = 32'hc405347;
      39795: inst = 32'h8220000;
      39796: inst = 32'h10408000;
      39797: inst = 32'hc405348;
      39798: inst = 32'h8220000;
      39799: inst = 32'h10408000;
      39800: inst = 32'hc405349;
      39801: inst = 32'h8220000;
      39802: inst = 32'h10408000;
      39803: inst = 32'hc40534a;
      39804: inst = 32'h8220000;
      39805: inst = 32'h10408000;
      39806: inst = 32'hc40534b;
      39807: inst = 32'h8220000;
      39808: inst = 32'h10408000;
      39809: inst = 32'hc40534c;
      39810: inst = 32'h8220000;
      39811: inst = 32'h10408000;
      39812: inst = 32'hc40534d;
      39813: inst = 32'h8220000;
      39814: inst = 32'h10408000;
      39815: inst = 32'hc40534e;
      39816: inst = 32'h8220000;
      39817: inst = 32'h10408000;
      39818: inst = 32'hc40534f;
      39819: inst = 32'h8220000;
      39820: inst = 32'h10408000;
      39821: inst = 32'hc405350;
      39822: inst = 32'h8220000;
      39823: inst = 32'h10408000;
      39824: inst = 32'hc405351;
      39825: inst = 32'h8220000;
      39826: inst = 32'h10408000;
      39827: inst = 32'hc40535c;
      39828: inst = 32'h8220000;
      39829: inst = 32'h10408000;
      39830: inst = 32'hc405363;
      39831: inst = 32'h8220000;
      39832: inst = 32'h10408000;
      39833: inst = 32'hc405364;
      39834: inst = 32'h8220000;
      39835: inst = 32'h10408000;
      39836: inst = 32'hc405365;
      39837: inst = 32'h8220000;
      39838: inst = 32'h10408000;
      39839: inst = 32'hc405366;
      39840: inst = 32'h8220000;
      39841: inst = 32'h10408000;
      39842: inst = 32'hc405367;
      39843: inst = 32'h8220000;
      39844: inst = 32'h10408000;
      39845: inst = 32'hc405368;
      39846: inst = 32'h8220000;
      39847: inst = 32'h10408000;
      39848: inst = 32'hc405369;
      39849: inst = 32'h8220000;
      39850: inst = 32'h10408000;
      39851: inst = 32'hc40536a;
      39852: inst = 32'h8220000;
      39853: inst = 32'h10408000;
      39854: inst = 32'hc40536b;
      39855: inst = 32'h8220000;
      39856: inst = 32'h10408000;
      39857: inst = 32'hc40536c;
      39858: inst = 32'h8220000;
      39859: inst = 32'h10408000;
      39860: inst = 32'hc40536d;
      39861: inst = 32'h8220000;
      39862: inst = 32'h10408000;
      39863: inst = 32'hc40536e;
      39864: inst = 32'h8220000;
      39865: inst = 32'h10408000;
      39866: inst = 32'hc40536f;
      39867: inst = 32'h8220000;
      39868: inst = 32'h10408000;
      39869: inst = 32'hc405370;
      39870: inst = 32'h8220000;
      39871: inst = 32'h10408000;
      39872: inst = 32'hc405371;
      39873: inst = 32'h8220000;
      39874: inst = 32'h10408000;
      39875: inst = 32'hc405372;
      39876: inst = 32'h8220000;
      39877: inst = 32'h10408000;
      39878: inst = 32'hc405373;
      39879: inst = 32'h8220000;
      39880: inst = 32'h10408000;
      39881: inst = 32'hc405374;
      39882: inst = 32'h8220000;
      39883: inst = 32'h10408000;
      39884: inst = 32'hc405375;
      39885: inst = 32'h8220000;
      39886: inst = 32'h10408000;
      39887: inst = 32'hc405379;
      39888: inst = 32'h8220000;
      39889: inst = 32'h10408000;
      39890: inst = 32'hc40537a;
      39891: inst = 32'h8220000;
      39892: inst = 32'h10408000;
      39893: inst = 32'hc40537b;
      39894: inst = 32'h8220000;
      39895: inst = 32'h10408000;
      39896: inst = 32'hc40537c;
      39897: inst = 32'h8220000;
      39898: inst = 32'h10408000;
      39899: inst = 32'hc40537d;
      39900: inst = 32'h8220000;
      39901: inst = 32'h10408000;
      39902: inst = 32'hc40537e;
      39903: inst = 32'h8220000;
      39904: inst = 32'h10408000;
      39905: inst = 32'hc40537f;
      39906: inst = 32'h8220000;
      39907: inst = 32'h10408000;
      39908: inst = 32'hc405380;
      39909: inst = 32'h8220000;
      39910: inst = 32'h10408000;
      39911: inst = 32'hc405381;
      39912: inst = 32'h8220000;
      39913: inst = 32'h10408000;
      39914: inst = 32'hc405382;
      39915: inst = 32'h8220000;
      39916: inst = 32'h10408000;
      39917: inst = 32'hc405383;
      39918: inst = 32'h8220000;
      39919: inst = 32'h10408000;
      39920: inst = 32'hc405384;
      39921: inst = 32'h8220000;
      39922: inst = 32'h10408000;
      39923: inst = 32'hc405385;
      39924: inst = 32'h8220000;
      39925: inst = 32'h10408000;
      39926: inst = 32'hc405386;
      39927: inst = 32'h8220000;
      39928: inst = 32'h10408000;
      39929: inst = 32'hc405387;
      39930: inst = 32'h8220000;
      39931: inst = 32'h10408000;
      39932: inst = 32'hc405388;
      39933: inst = 32'h8220000;
      39934: inst = 32'h10408000;
      39935: inst = 32'hc405389;
      39936: inst = 32'h8220000;
      39937: inst = 32'h10408000;
      39938: inst = 32'hc40538a;
      39939: inst = 32'h8220000;
      39940: inst = 32'h10408000;
      39941: inst = 32'hc40538b;
      39942: inst = 32'h8220000;
      39943: inst = 32'h10408000;
      39944: inst = 32'hc40538c;
      39945: inst = 32'h8220000;
      39946: inst = 32'h10408000;
      39947: inst = 32'hc40538d;
      39948: inst = 32'h8220000;
      39949: inst = 32'h10408000;
      39950: inst = 32'hc40538e;
      39951: inst = 32'h8220000;
      39952: inst = 32'h10408000;
      39953: inst = 32'hc40538f;
      39954: inst = 32'h8220000;
      39955: inst = 32'h10408000;
      39956: inst = 32'hc405390;
      39957: inst = 32'h8220000;
      39958: inst = 32'h10408000;
      39959: inst = 32'hc405391;
      39960: inst = 32'h8220000;
      39961: inst = 32'h10408000;
      39962: inst = 32'hc405392;
      39963: inst = 32'h8220000;
      39964: inst = 32'h10408000;
      39965: inst = 32'hc405393;
      39966: inst = 32'h8220000;
      39967: inst = 32'h10408000;
      39968: inst = 32'hc405394;
      39969: inst = 32'h8220000;
      39970: inst = 32'h10408000;
      39971: inst = 32'hc405395;
      39972: inst = 32'h8220000;
      39973: inst = 32'h10408000;
      39974: inst = 32'hc405396;
      39975: inst = 32'h8220000;
      39976: inst = 32'h10408000;
      39977: inst = 32'hc405397;
      39978: inst = 32'h8220000;
      39979: inst = 32'h10408000;
      39980: inst = 32'hc405398;
      39981: inst = 32'h8220000;
      39982: inst = 32'h10408000;
      39983: inst = 32'hc405399;
      39984: inst = 32'h8220000;
      39985: inst = 32'h10408000;
      39986: inst = 32'hc40539a;
      39987: inst = 32'h8220000;
      39988: inst = 32'h10408000;
      39989: inst = 32'hc40539b;
      39990: inst = 32'h8220000;
      39991: inst = 32'h10408000;
      39992: inst = 32'hc40539c;
      39993: inst = 32'h8220000;
      39994: inst = 32'h10408000;
      39995: inst = 32'hc40539d;
      39996: inst = 32'h8220000;
      39997: inst = 32'h10408000;
      39998: inst = 32'hc40539e;
      39999: inst = 32'h8220000;
      40000: inst = 32'h10408000;
      40001: inst = 32'hc40539f;
      40002: inst = 32'h8220000;
      40003: inst = 32'h10408000;
      40004: inst = 32'hc4053a0;
      40005: inst = 32'h8220000;
      40006: inst = 32'h10408000;
      40007: inst = 32'hc4053a1;
      40008: inst = 32'h8220000;
      40009: inst = 32'h10408000;
      40010: inst = 32'hc4053a2;
      40011: inst = 32'h8220000;
      40012: inst = 32'h10408000;
      40013: inst = 32'hc4053a3;
      40014: inst = 32'h8220000;
      40015: inst = 32'h10408000;
      40016: inst = 32'hc4053a4;
      40017: inst = 32'h8220000;
      40018: inst = 32'h10408000;
      40019: inst = 32'hc4053a5;
      40020: inst = 32'h8220000;
      40021: inst = 32'h10408000;
      40022: inst = 32'hc4053a6;
      40023: inst = 32'h8220000;
      40024: inst = 32'h10408000;
      40025: inst = 32'hc4053a7;
      40026: inst = 32'h8220000;
      40027: inst = 32'h10408000;
      40028: inst = 32'hc4053a8;
      40029: inst = 32'h8220000;
      40030: inst = 32'h10408000;
      40031: inst = 32'hc4053a9;
      40032: inst = 32'h8220000;
      40033: inst = 32'h10408000;
      40034: inst = 32'hc4053aa;
      40035: inst = 32'h8220000;
      40036: inst = 32'h10408000;
      40037: inst = 32'hc4053ab;
      40038: inst = 32'h8220000;
      40039: inst = 32'h10408000;
      40040: inst = 32'hc4053ac;
      40041: inst = 32'h8220000;
      40042: inst = 32'h10408000;
      40043: inst = 32'hc4053ad;
      40044: inst = 32'h8220000;
      40045: inst = 32'h10408000;
      40046: inst = 32'hc4053ae;
      40047: inst = 32'h8220000;
      40048: inst = 32'h10408000;
      40049: inst = 32'hc4053af;
      40050: inst = 32'h8220000;
      40051: inst = 32'h10408000;
      40052: inst = 32'hc4053b0;
      40053: inst = 32'h8220000;
      40054: inst = 32'h10408000;
      40055: inst = 32'hc4053b1;
      40056: inst = 32'h8220000;
      40057: inst = 32'h10408000;
      40058: inst = 32'hc4053bc;
      40059: inst = 32'h8220000;
      40060: inst = 32'h10408000;
      40061: inst = 32'hc4053c3;
      40062: inst = 32'h8220000;
      40063: inst = 32'h10408000;
      40064: inst = 32'hc4053c4;
      40065: inst = 32'h8220000;
      40066: inst = 32'h10408000;
      40067: inst = 32'hc4053c5;
      40068: inst = 32'h8220000;
      40069: inst = 32'h10408000;
      40070: inst = 32'hc4053c6;
      40071: inst = 32'h8220000;
      40072: inst = 32'h10408000;
      40073: inst = 32'hc4053c7;
      40074: inst = 32'h8220000;
      40075: inst = 32'h10408000;
      40076: inst = 32'hc4053cf;
      40077: inst = 32'h8220000;
      40078: inst = 32'h10408000;
      40079: inst = 32'hc4053d0;
      40080: inst = 32'h8220000;
      40081: inst = 32'h10408000;
      40082: inst = 32'hc4053d1;
      40083: inst = 32'h8220000;
      40084: inst = 32'h10408000;
      40085: inst = 32'hc4053d2;
      40086: inst = 32'h8220000;
      40087: inst = 32'h10408000;
      40088: inst = 32'hc4053d3;
      40089: inst = 32'h8220000;
      40090: inst = 32'h10408000;
      40091: inst = 32'hc4053d4;
      40092: inst = 32'h8220000;
      40093: inst = 32'h10408000;
      40094: inst = 32'hc4053d5;
      40095: inst = 32'h8220000;
      40096: inst = 32'h10408000;
      40097: inst = 32'hc4053d9;
      40098: inst = 32'h8220000;
      40099: inst = 32'h10408000;
      40100: inst = 32'hc4053da;
      40101: inst = 32'h8220000;
      40102: inst = 32'h10408000;
      40103: inst = 32'hc4053db;
      40104: inst = 32'h8220000;
      40105: inst = 32'h10408000;
      40106: inst = 32'hc4053dc;
      40107: inst = 32'h8220000;
      40108: inst = 32'h10408000;
      40109: inst = 32'hc4053dd;
      40110: inst = 32'h8220000;
      40111: inst = 32'h10408000;
      40112: inst = 32'hc4053de;
      40113: inst = 32'h8220000;
      40114: inst = 32'h10408000;
      40115: inst = 32'hc4053df;
      40116: inst = 32'h8220000;
      40117: inst = 32'h10408000;
      40118: inst = 32'hc4053e0;
      40119: inst = 32'h8220000;
      40120: inst = 32'h10408000;
      40121: inst = 32'hc4053e1;
      40122: inst = 32'h8220000;
      40123: inst = 32'h10408000;
      40124: inst = 32'hc4053e2;
      40125: inst = 32'h8220000;
      40126: inst = 32'h10408000;
      40127: inst = 32'hc4053e3;
      40128: inst = 32'h8220000;
      40129: inst = 32'h10408000;
      40130: inst = 32'hc4053e4;
      40131: inst = 32'h8220000;
      40132: inst = 32'h10408000;
      40133: inst = 32'hc4053e5;
      40134: inst = 32'h8220000;
      40135: inst = 32'h10408000;
      40136: inst = 32'hc4053e6;
      40137: inst = 32'h8220000;
      40138: inst = 32'h10408000;
      40139: inst = 32'hc4053e7;
      40140: inst = 32'h8220000;
      40141: inst = 32'h10408000;
      40142: inst = 32'hc4053e8;
      40143: inst = 32'h8220000;
      40144: inst = 32'h10408000;
      40145: inst = 32'hc4053e9;
      40146: inst = 32'h8220000;
      40147: inst = 32'h10408000;
      40148: inst = 32'hc4053ea;
      40149: inst = 32'h8220000;
      40150: inst = 32'h10408000;
      40151: inst = 32'hc4053eb;
      40152: inst = 32'h8220000;
      40153: inst = 32'h10408000;
      40154: inst = 32'hc4053ec;
      40155: inst = 32'h8220000;
      40156: inst = 32'h10408000;
      40157: inst = 32'hc4053ed;
      40158: inst = 32'h8220000;
      40159: inst = 32'h10408000;
      40160: inst = 32'hc4053ee;
      40161: inst = 32'h8220000;
      40162: inst = 32'h10408000;
      40163: inst = 32'hc4053ef;
      40164: inst = 32'h8220000;
      40165: inst = 32'h10408000;
      40166: inst = 32'hc4053f0;
      40167: inst = 32'h8220000;
      40168: inst = 32'h10408000;
      40169: inst = 32'hc4053f1;
      40170: inst = 32'h8220000;
      40171: inst = 32'h10408000;
      40172: inst = 32'hc4053f2;
      40173: inst = 32'h8220000;
      40174: inst = 32'h10408000;
      40175: inst = 32'hc4053f3;
      40176: inst = 32'h8220000;
      40177: inst = 32'h10408000;
      40178: inst = 32'hc4053f4;
      40179: inst = 32'h8220000;
      40180: inst = 32'h10408000;
      40181: inst = 32'hc4053f5;
      40182: inst = 32'h8220000;
      40183: inst = 32'h10408000;
      40184: inst = 32'hc4053f6;
      40185: inst = 32'h8220000;
      40186: inst = 32'h10408000;
      40187: inst = 32'hc4053f7;
      40188: inst = 32'h8220000;
      40189: inst = 32'h10408000;
      40190: inst = 32'hc4053f8;
      40191: inst = 32'h8220000;
      40192: inst = 32'h10408000;
      40193: inst = 32'hc4053f9;
      40194: inst = 32'h8220000;
      40195: inst = 32'h10408000;
      40196: inst = 32'hc4053fa;
      40197: inst = 32'h8220000;
      40198: inst = 32'h10408000;
      40199: inst = 32'hc4053fb;
      40200: inst = 32'h8220000;
      40201: inst = 32'h10408000;
      40202: inst = 32'hc4053fc;
      40203: inst = 32'h8220000;
      40204: inst = 32'h10408000;
      40205: inst = 32'hc4053fd;
      40206: inst = 32'h8220000;
      40207: inst = 32'h10408000;
      40208: inst = 32'hc4053fe;
      40209: inst = 32'h8220000;
      40210: inst = 32'h10408000;
      40211: inst = 32'hc4053ff;
      40212: inst = 32'h8220000;
      40213: inst = 32'h10408000;
      40214: inst = 32'hc405400;
      40215: inst = 32'h8220000;
      40216: inst = 32'h10408000;
      40217: inst = 32'hc405401;
      40218: inst = 32'h8220000;
      40219: inst = 32'h10408000;
      40220: inst = 32'hc405402;
      40221: inst = 32'h8220000;
      40222: inst = 32'h10408000;
      40223: inst = 32'hc405403;
      40224: inst = 32'h8220000;
      40225: inst = 32'h10408000;
      40226: inst = 32'hc405404;
      40227: inst = 32'h8220000;
      40228: inst = 32'h10408000;
      40229: inst = 32'hc405405;
      40230: inst = 32'h8220000;
      40231: inst = 32'h10408000;
      40232: inst = 32'hc405406;
      40233: inst = 32'h8220000;
      40234: inst = 32'h10408000;
      40235: inst = 32'hc405407;
      40236: inst = 32'h8220000;
      40237: inst = 32'h10408000;
      40238: inst = 32'hc405408;
      40239: inst = 32'h8220000;
      40240: inst = 32'h10408000;
      40241: inst = 32'hc405409;
      40242: inst = 32'h8220000;
      40243: inst = 32'h10408000;
      40244: inst = 32'hc40540a;
      40245: inst = 32'h8220000;
      40246: inst = 32'h10408000;
      40247: inst = 32'hc40540b;
      40248: inst = 32'h8220000;
      40249: inst = 32'h10408000;
      40250: inst = 32'hc40540c;
      40251: inst = 32'h8220000;
      40252: inst = 32'h10408000;
      40253: inst = 32'hc40540d;
      40254: inst = 32'h8220000;
      40255: inst = 32'h10408000;
      40256: inst = 32'hc40540e;
      40257: inst = 32'h8220000;
      40258: inst = 32'h10408000;
      40259: inst = 32'hc40540f;
      40260: inst = 32'h8220000;
      40261: inst = 32'h10408000;
      40262: inst = 32'hc405410;
      40263: inst = 32'h8220000;
      40264: inst = 32'h10408000;
      40265: inst = 32'hc405411;
      40266: inst = 32'h8220000;
      40267: inst = 32'h10408000;
      40268: inst = 32'hc40541c;
      40269: inst = 32'h8220000;
      40270: inst = 32'h10408000;
      40271: inst = 32'hc405423;
      40272: inst = 32'h8220000;
      40273: inst = 32'h10408000;
      40274: inst = 32'hc405424;
      40275: inst = 32'h8220000;
      40276: inst = 32'h10408000;
      40277: inst = 32'hc405425;
      40278: inst = 32'h8220000;
      40279: inst = 32'h10408000;
      40280: inst = 32'hc405426;
      40281: inst = 32'h8220000;
      40282: inst = 32'h10408000;
      40283: inst = 32'hc405430;
      40284: inst = 32'h8220000;
      40285: inst = 32'h10408000;
      40286: inst = 32'hc405431;
      40287: inst = 32'h8220000;
      40288: inst = 32'h10408000;
      40289: inst = 32'hc405432;
      40290: inst = 32'h8220000;
      40291: inst = 32'h10408000;
      40292: inst = 32'hc405433;
      40293: inst = 32'h8220000;
      40294: inst = 32'h10408000;
      40295: inst = 32'hc405434;
      40296: inst = 32'h8220000;
      40297: inst = 32'h10408000;
      40298: inst = 32'hc405435;
      40299: inst = 32'h8220000;
      40300: inst = 32'h10408000;
      40301: inst = 32'hc40544a;
      40302: inst = 32'h8220000;
      40303: inst = 32'h10408000;
      40304: inst = 32'hc40544b;
      40305: inst = 32'h8220000;
      40306: inst = 32'h10408000;
      40307: inst = 32'hc40544c;
      40308: inst = 32'h8220000;
      40309: inst = 32'h10408000;
      40310: inst = 32'hc40544d;
      40311: inst = 32'h8220000;
      40312: inst = 32'h10408000;
      40313: inst = 32'hc40544e;
      40314: inst = 32'h8220000;
      40315: inst = 32'h10408000;
      40316: inst = 32'hc40544f;
      40317: inst = 32'h8220000;
      40318: inst = 32'h10408000;
      40319: inst = 32'hc405450;
      40320: inst = 32'h8220000;
      40321: inst = 32'h10408000;
      40322: inst = 32'hc405451;
      40323: inst = 32'h8220000;
      40324: inst = 32'h10408000;
      40325: inst = 32'hc405452;
      40326: inst = 32'h8220000;
      40327: inst = 32'h10408000;
      40328: inst = 32'hc405453;
      40329: inst = 32'h8220000;
      40330: inst = 32'h10408000;
      40331: inst = 32'hc405454;
      40332: inst = 32'h8220000;
      40333: inst = 32'h10408000;
      40334: inst = 32'hc405455;
      40335: inst = 32'h8220000;
      40336: inst = 32'h10408000;
      40337: inst = 32'hc405456;
      40338: inst = 32'h8220000;
      40339: inst = 32'h10408000;
      40340: inst = 32'hc405457;
      40341: inst = 32'h8220000;
      40342: inst = 32'h10408000;
      40343: inst = 32'hc405458;
      40344: inst = 32'h8220000;
      40345: inst = 32'h10408000;
      40346: inst = 32'hc405459;
      40347: inst = 32'h8220000;
      40348: inst = 32'h10408000;
      40349: inst = 32'hc40545a;
      40350: inst = 32'h8220000;
      40351: inst = 32'h10408000;
      40352: inst = 32'hc40545b;
      40353: inst = 32'h8220000;
      40354: inst = 32'h10408000;
      40355: inst = 32'hc40545c;
      40356: inst = 32'h8220000;
      40357: inst = 32'h10408000;
      40358: inst = 32'hc40545d;
      40359: inst = 32'h8220000;
      40360: inst = 32'h10408000;
      40361: inst = 32'hc40545e;
      40362: inst = 32'h8220000;
      40363: inst = 32'h10408000;
      40364: inst = 32'hc40545f;
      40365: inst = 32'h8220000;
      40366: inst = 32'h10408000;
      40367: inst = 32'hc405460;
      40368: inst = 32'h8220000;
      40369: inst = 32'h10408000;
      40370: inst = 32'hc405461;
      40371: inst = 32'h8220000;
      40372: inst = 32'h10408000;
      40373: inst = 32'hc405462;
      40374: inst = 32'h8220000;
      40375: inst = 32'h10408000;
      40376: inst = 32'hc405463;
      40377: inst = 32'h8220000;
      40378: inst = 32'h10408000;
      40379: inst = 32'hc405464;
      40380: inst = 32'h8220000;
      40381: inst = 32'h10408000;
      40382: inst = 32'hc405465;
      40383: inst = 32'h8220000;
      40384: inst = 32'h10408000;
      40385: inst = 32'hc405466;
      40386: inst = 32'h8220000;
      40387: inst = 32'h10408000;
      40388: inst = 32'hc405467;
      40389: inst = 32'h8220000;
      40390: inst = 32'h10408000;
      40391: inst = 32'hc405468;
      40392: inst = 32'h8220000;
      40393: inst = 32'h10408000;
      40394: inst = 32'hc405469;
      40395: inst = 32'h8220000;
      40396: inst = 32'h10408000;
      40397: inst = 32'hc40546a;
      40398: inst = 32'h8220000;
      40399: inst = 32'h10408000;
      40400: inst = 32'hc40546b;
      40401: inst = 32'h8220000;
      40402: inst = 32'h10408000;
      40403: inst = 32'hc40546c;
      40404: inst = 32'h8220000;
      40405: inst = 32'h10408000;
      40406: inst = 32'hc40546d;
      40407: inst = 32'h8220000;
      40408: inst = 32'h10408000;
      40409: inst = 32'hc40546e;
      40410: inst = 32'h8220000;
      40411: inst = 32'h10408000;
      40412: inst = 32'hc40546f;
      40413: inst = 32'h8220000;
      40414: inst = 32'h10408000;
      40415: inst = 32'hc405470;
      40416: inst = 32'h8220000;
      40417: inst = 32'h10408000;
      40418: inst = 32'hc405471;
      40419: inst = 32'h8220000;
      40420: inst = 32'h10408000;
      40421: inst = 32'hc40547c;
      40422: inst = 32'h8220000;
      40423: inst = 32'h10408000;
      40424: inst = 32'hc405483;
      40425: inst = 32'h8220000;
      40426: inst = 32'h10408000;
      40427: inst = 32'hc405484;
      40428: inst = 32'h8220000;
      40429: inst = 32'h10408000;
      40430: inst = 32'hc405485;
      40431: inst = 32'h8220000;
      40432: inst = 32'h10408000;
      40433: inst = 32'hc405486;
      40434: inst = 32'h8220000;
      40435: inst = 32'h10408000;
      40436: inst = 32'hc405490;
      40437: inst = 32'h8220000;
      40438: inst = 32'h10408000;
      40439: inst = 32'hc405491;
      40440: inst = 32'h8220000;
      40441: inst = 32'h10408000;
      40442: inst = 32'hc405492;
      40443: inst = 32'h8220000;
      40444: inst = 32'h10408000;
      40445: inst = 32'hc405493;
      40446: inst = 32'h8220000;
      40447: inst = 32'h10408000;
      40448: inst = 32'hc405494;
      40449: inst = 32'h8220000;
      40450: inst = 32'h10408000;
      40451: inst = 32'hc405495;
      40452: inst = 32'h8220000;
      40453: inst = 32'h10408000;
      40454: inst = 32'hc4054aa;
      40455: inst = 32'h8220000;
      40456: inst = 32'h10408000;
      40457: inst = 32'hc4054ab;
      40458: inst = 32'h8220000;
      40459: inst = 32'h10408000;
      40460: inst = 32'hc4054ac;
      40461: inst = 32'h8220000;
      40462: inst = 32'h10408000;
      40463: inst = 32'hc4054ad;
      40464: inst = 32'h8220000;
      40465: inst = 32'h10408000;
      40466: inst = 32'hc4054ae;
      40467: inst = 32'h8220000;
      40468: inst = 32'h10408000;
      40469: inst = 32'hc4054af;
      40470: inst = 32'h8220000;
      40471: inst = 32'h10408000;
      40472: inst = 32'hc4054b0;
      40473: inst = 32'h8220000;
      40474: inst = 32'h10408000;
      40475: inst = 32'hc4054b1;
      40476: inst = 32'h8220000;
      40477: inst = 32'h10408000;
      40478: inst = 32'hc4054b2;
      40479: inst = 32'h8220000;
      40480: inst = 32'h10408000;
      40481: inst = 32'hc4054b3;
      40482: inst = 32'h8220000;
      40483: inst = 32'h10408000;
      40484: inst = 32'hc4054b4;
      40485: inst = 32'h8220000;
      40486: inst = 32'h10408000;
      40487: inst = 32'hc4054b5;
      40488: inst = 32'h8220000;
      40489: inst = 32'h10408000;
      40490: inst = 32'hc4054b6;
      40491: inst = 32'h8220000;
      40492: inst = 32'h10408000;
      40493: inst = 32'hc4054b7;
      40494: inst = 32'h8220000;
      40495: inst = 32'h10408000;
      40496: inst = 32'hc4054b8;
      40497: inst = 32'h8220000;
      40498: inst = 32'h10408000;
      40499: inst = 32'hc4054b9;
      40500: inst = 32'h8220000;
      40501: inst = 32'h10408000;
      40502: inst = 32'hc4054ba;
      40503: inst = 32'h8220000;
      40504: inst = 32'h10408000;
      40505: inst = 32'hc4054bb;
      40506: inst = 32'h8220000;
      40507: inst = 32'h10408000;
      40508: inst = 32'hc4054bc;
      40509: inst = 32'h8220000;
      40510: inst = 32'h10408000;
      40511: inst = 32'hc4054bd;
      40512: inst = 32'h8220000;
      40513: inst = 32'h10408000;
      40514: inst = 32'hc4054be;
      40515: inst = 32'h8220000;
      40516: inst = 32'h10408000;
      40517: inst = 32'hc4054bf;
      40518: inst = 32'h8220000;
      40519: inst = 32'h10408000;
      40520: inst = 32'hc4054c0;
      40521: inst = 32'h8220000;
      40522: inst = 32'h10408000;
      40523: inst = 32'hc4054c1;
      40524: inst = 32'h8220000;
      40525: inst = 32'h10408000;
      40526: inst = 32'hc4054c2;
      40527: inst = 32'h8220000;
      40528: inst = 32'h10408000;
      40529: inst = 32'hc4054c3;
      40530: inst = 32'h8220000;
      40531: inst = 32'h10408000;
      40532: inst = 32'hc4054c4;
      40533: inst = 32'h8220000;
      40534: inst = 32'h10408000;
      40535: inst = 32'hc4054c5;
      40536: inst = 32'h8220000;
      40537: inst = 32'h10408000;
      40538: inst = 32'hc4054c6;
      40539: inst = 32'h8220000;
      40540: inst = 32'h10408000;
      40541: inst = 32'hc4054c7;
      40542: inst = 32'h8220000;
      40543: inst = 32'h10408000;
      40544: inst = 32'hc4054c8;
      40545: inst = 32'h8220000;
      40546: inst = 32'h10408000;
      40547: inst = 32'hc4054c9;
      40548: inst = 32'h8220000;
      40549: inst = 32'h10408000;
      40550: inst = 32'hc4054ca;
      40551: inst = 32'h8220000;
      40552: inst = 32'h10408000;
      40553: inst = 32'hc4054cb;
      40554: inst = 32'h8220000;
      40555: inst = 32'h10408000;
      40556: inst = 32'hc4054cc;
      40557: inst = 32'h8220000;
      40558: inst = 32'h10408000;
      40559: inst = 32'hc4054cd;
      40560: inst = 32'h8220000;
      40561: inst = 32'h10408000;
      40562: inst = 32'hc4054ce;
      40563: inst = 32'h8220000;
      40564: inst = 32'h10408000;
      40565: inst = 32'hc4054cf;
      40566: inst = 32'h8220000;
      40567: inst = 32'h10408000;
      40568: inst = 32'hc4054d0;
      40569: inst = 32'h8220000;
      40570: inst = 32'h10408000;
      40571: inst = 32'hc4054d1;
      40572: inst = 32'h8220000;
      40573: inst = 32'h10408000;
      40574: inst = 32'hc4054dc;
      40575: inst = 32'h8220000;
      40576: inst = 32'h10408000;
      40577: inst = 32'hc4054e3;
      40578: inst = 32'h8220000;
      40579: inst = 32'h10408000;
      40580: inst = 32'hc4054e4;
      40581: inst = 32'h8220000;
      40582: inst = 32'h10408000;
      40583: inst = 32'hc4054e5;
      40584: inst = 32'h8220000;
      40585: inst = 32'h10408000;
      40586: inst = 32'hc4054e6;
      40587: inst = 32'h8220000;
      40588: inst = 32'h10408000;
      40589: inst = 32'hc4054f0;
      40590: inst = 32'h8220000;
      40591: inst = 32'h10408000;
      40592: inst = 32'hc4054f1;
      40593: inst = 32'h8220000;
      40594: inst = 32'h10408000;
      40595: inst = 32'hc4054f2;
      40596: inst = 32'h8220000;
      40597: inst = 32'h10408000;
      40598: inst = 32'hc4054f3;
      40599: inst = 32'h8220000;
      40600: inst = 32'h10408000;
      40601: inst = 32'hc4054f4;
      40602: inst = 32'h8220000;
      40603: inst = 32'h10408000;
      40604: inst = 32'hc4054f5;
      40605: inst = 32'h8220000;
      40606: inst = 32'h10408000;
      40607: inst = 32'hc40550a;
      40608: inst = 32'h8220000;
      40609: inst = 32'h10408000;
      40610: inst = 32'hc40550b;
      40611: inst = 32'h8220000;
      40612: inst = 32'h10408000;
      40613: inst = 32'hc40550c;
      40614: inst = 32'h8220000;
      40615: inst = 32'h10408000;
      40616: inst = 32'hc40550d;
      40617: inst = 32'h8220000;
      40618: inst = 32'h10408000;
      40619: inst = 32'hc40550e;
      40620: inst = 32'h8220000;
      40621: inst = 32'h10408000;
      40622: inst = 32'hc40550f;
      40623: inst = 32'h8220000;
      40624: inst = 32'h10408000;
      40625: inst = 32'hc405510;
      40626: inst = 32'h8220000;
      40627: inst = 32'h10408000;
      40628: inst = 32'hc405511;
      40629: inst = 32'h8220000;
      40630: inst = 32'h10408000;
      40631: inst = 32'hc405512;
      40632: inst = 32'h8220000;
      40633: inst = 32'h10408000;
      40634: inst = 32'hc405513;
      40635: inst = 32'h8220000;
      40636: inst = 32'h10408000;
      40637: inst = 32'hc405514;
      40638: inst = 32'h8220000;
      40639: inst = 32'h10408000;
      40640: inst = 32'hc405515;
      40641: inst = 32'h8220000;
      40642: inst = 32'h10408000;
      40643: inst = 32'hc405516;
      40644: inst = 32'h8220000;
      40645: inst = 32'h10408000;
      40646: inst = 32'hc405517;
      40647: inst = 32'h8220000;
      40648: inst = 32'h10408000;
      40649: inst = 32'hc405518;
      40650: inst = 32'h8220000;
      40651: inst = 32'h10408000;
      40652: inst = 32'hc405519;
      40653: inst = 32'h8220000;
      40654: inst = 32'h10408000;
      40655: inst = 32'hc40551a;
      40656: inst = 32'h8220000;
      40657: inst = 32'h10408000;
      40658: inst = 32'hc40551b;
      40659: inst = 32'h8220000;
      40660: inst = 32'h10408000;
      40661: inst = 32'hc40551c;
      40662: inst = 32'h8220000;
      40663: inst = 32'h10408000;
      40664: inst = 32'hc40551d;
      40665: inst = 32'h8220000;
      40666: inst = 32'h10408000;
      40667: inst = 32'hc40551e;
      40668: inst = 32'h8220000;
      40669: inst = 32'h10408000;
      40670: inst = 32'hc40551f;
      40671: inst = 32'h8220000;
      40672: inst = 32'h10408000;
      40673: inst = 32'hc405520;
      40674: inst = 32'h8220000;
      40675: inst = 32'h10408000;
      40676: inst = 32'hc405521;
      40677: inst = 32'h8220000;
      40678: inst = 32'h10408000;
      40679: inst = 32'hc405522;
      40680: inst = 32'h8220000;
      40681: inst = 32'h10408000;
      40682: inst = 32'hc405523;
      40683: inst = 32'h8220000;
      40684: inst = 32'h10408000;
      40685: inst = 32'hc405524;
      40686: inst = 32'h8220000;
      40687: inst = 32'h10408000;
      40688: inst = 32'hc405525;
      40689: inst = 32'h8220000;
      40690: inst = 32'h10408000;
      40691: inst = 32'hc405526;
      40692: inst = 32'h8220000;
      40693: inst = 32'h10408000;
      40694: inst = 32'hc405527;
      40695: inst = 32'h8220000;
      40696: inst = 32'h10408000;
      40697: inst = 32'hc405528;
      40698: inst = 32'h8220000;
      40699: inst = 32'h10408000;
      40700: inst = 32'hc405529;
      40701: inst = 32'h8220000;
      40702: inst = 32'h10408000;
      40703: inst = 32'hc40552a;
      40704: inst = 32'h8220000;
      40705: inst = 32'h10408000;
      40706: inst = 32'hc40552b;
      40707: inst = 32'h8220000;
      40708: inst = 32'h10408000;
      40709: inst = 32'hc40552c;
      40710: inst = 32'h8220000;
      40711: inst = 32'h10408000;
      40712: inst = 32'hc40552d;
      40713: inst = 32'h8220000;
      40714: inst = 32'h10408000;
      40715: inst = 32'hc40552e;
      40716: inst = 32'h8220000;
      40717: inst = 32'h10408000;
      40718: inst = 32'hc40552f;
      40719: inst = 32'h8220000;
      40720: inst = 32'h10408000;
      40721: inst = 32'hc405530;
      40722: inst = 32'h8220000;
      40723: inst = 32'h10408000;
      40724: inst = 32'hc405531;
      40725: inst = 32'h8220000;
      40726: inst = 32'h10408000;
      40727: inst = 32'hc40553c;
      40728: inst = 32'h8220000;
      40729: inst = 32'h10408000;
      40730: inst = 32'hc405543;
      40731: inst = 32'h8220000;
      40732: inst = 32'h10408000;
      40733: inst = 32'hc405544;
      40734: inst = 32'h8220000;
      40735: inst = 32'h10408000;
      40736: inst = 32'hc405545;
      40737: inst = 32'h8220000;
      40738: inst = 32'h10408000;
      40739: inst = 32'hc405546;
      40740: inst = 32'h8220000;
      40741: inst = 32'h10408000;
      40742: inst = 32'hc405550;
      40743: inst = 32'h8220000;
      40744: inst = 32'h10408000;
      40745: inst = 32'hc405551;
      40746: inst = 32'h8220000;
      40747: inst = 32'h10408000;
      40748: inst = 32'hc405552;
      40749: inst = 32'h8220000;
      40750: inst = 32'h10408000;
      40751: inst = 32'hc405553;
      40752: inst = 32'h8220000;
      40753: inst = 32'h10408000;
      40754: inst = 32'hc405554;
      40755: inst = 32'h8220000;
      40756: inst = 32'h10408000;
      40757: inst = 32'hc405555;
      40758: inst = 32'h8220000;
      40759: inst = 32'h10408000;
      40760: inst = 32'hc405559;
      40761: inst = 32'h8220000;
      40762: inst = 32'h10408000;
      40763: inst = 32'hc40555a;
      40764: inst = 32'h8220000;
      40765: inst = 32'h10408000;
      40766: inst = 32'hc40555b;
      40767: inst = 32'h8220000;
      40768: inst = 32'h10408000;
      40769: inst = 32'hc40555c;
      40770: inst = 32'h8220000;
      40771: inst = 32'h10408000;
      40772: inst = 32'hc40555d;
      40773: inst = 32'h8220000;
      40774: inst = 32'h10408000;
      40775: inst = 32'hc40555e;
      40776: inst = 32'h8220000;
      40777: inst = 32'h10408000;
      40778: inst = 32'hc40555f;
      40779: inst = 32'h8220000;
      40780: inst = 32'h10408000;
      40781: inst = 32'hc405560;
      40782: inst = 32'h8220000;
      40783: inst = 32'h10408000;
      40784: inst = 32'hc405561;
      40785: inst = 32'h8220000;
      40786: inst = 32'h10408000;
      40787: inst = 32'hc405562;
      40788: inst = 32'h8220000;
      40789: inst = 32'h10408000;
      40790: inst = 32'hc405563;
      40791: inst = 32'h8220000;
      40792: inst = 32'h10408000;
      40793: inst = 32'hc405564;
      40794: inst = 32'h8220000;
      40795: inst = 32'h10408000;
      40796: inst = 32'hc405565;
      40797: inst = 32'h8220000;
      40798: inst = 32'h10408000;
      40799: inst = 32'hc405566;
      40800: inst = 32'h8220000;
      40801: inst = 32'h10408000;
      40802: inst = 32'hc405567;
      40803: inst = 32'h8220000;
      40804: inst = 32'h10408000;
      40805: inst = 32'hc405568;
      40806: inst = 32'h8220000;
      40807: inst = 32'h10408000;
      40808: inst = 32'hc405569;
      40809: inst = 32'h8220000;
      40810: inst = 32'h10408000;
      40811: inst = 32'hc40556a;
      40812: inst = 32'h8220000;
      40813: inst = 32'h10408000;
      40814: inst = 32'hc40556b;
      40815: inst = 32'h8220000;
      40816: inst = 32'h10408000;
      40817: inst = 32'hc40556c;
      40818: inst = 32'h8220000;
      40819: inst = 32'h10408000;
      40820: inst = 32'hc40556d;
      40821: inst = 32'h8220000;
      40822: inst = 32'h10408000;
      40823: inst = 32'hc40556e;
      40824: inst = 32'h8220000;
      40825: inst = 32'h10408000;
      40826: inst = 32'hc40556f;
      40827: inst = 32'h8220000;
      40828: inst = 32'h10408000;
      40829: inst = 32'hc405570;
      40830: inst = 32'h8220000;
      40831: inst = 32'h10408000;
      40832: inst = 32'hc405571;
      40833: inst = 32'h8220000;
      40834: inst = 32'h10408000;
      40835: inst = 32'hc405572;
      40836: inst = 32'h8220000;
      40837: inst = 32'h10408000;
      40838: inst = 32'hc405573;
      40839: inst = 32'h8220000;
      40840: inst = 32'h10408000;
      40841: inst = 32'hc405574;
      40842: inst = 32'h8220000;
      40843: inst = 32'h10408000;
      40844: inst = 32'hc405575;
      40845: inst = 32'h8220000;
      40846: inst = 32'h10408000;
      40847: inst = 32'hc405576;
      40848: inst = 32'h8220000;
      40849: inst = 32'h10408000;
      40850: inst = 32'hc405577;
      40851: inst = 32'h8220000;
      40852: inst = 32'h10408000;
      40853: inst = 32'hc405578;
      40854: inst = 32'h8220000;
      40855: inst = 32'h10408000;
      40856: inst = 32'hc405579;
      40857: inst = 32'h8220000;
      40858: inst = 32'h10408000;
      40859: inst = 32'hc40557a;
      40860: inst = 32'h8220000;
      40861: inst = 32'h10408000;
      40862: inst = 32'hc40557b;
      40863: inst = 32'h8220000;
      40864: inst = 32'h10408000;
      40865: inst = 32'hc40557c;
      40866: inst = 32'h8220000;
      40867: inst = 32'h10408000;
      40868: inst = 32'hc40557d;
      40869: inst = 32'h8220000;
      40870: inst = 32'h10408000;
      40871: inst = 32'hc40557e;
      40872: inst = 32'h8220000;
      40873: inst = 32'h10408000;
      40874: inst = 32'hc40557f;
      40875: inst = 32'h8220000;
      40876: inst = 32'h10408000;
      40877: inst = 32'hc405580;
      40878: inst = 32'h8220000;
      40879: inst = 32'h10408000;
      40880: inst = 32'hc405581;
      40881: inst = 32'h8220000;
      40882: inst = 32'h10408000;
      40883: inst = 32'hc405582;
      40884: inst = 32'h8220000;
      40885: inst = 32'h10408000;
      40886: inst = 32'hc405583;
      40887: inst = 32'h8220000;
      40888: inst = 32'h10408000;
      40889: inst = 32'hc405584;
      40890: inst = 32'h8220000;
      40891: inst = 32'h10408000;
      40892: inst = 32'hc405585;
      40893: inst = 32'h8220000;
      40894: inst = 32'h10408000;
      40895: inst = 32'hc405586;
      40896: inst = 32'h8220000;
      40897: inst = 32'h10408000;
      40898: inst = 32'hc405587;
      40899: inst = 32'h8220000;
      40900: inst = 32'h10408000;
      40901: inst = 32'hc405588;
      40902: inst = 32'h8220000;
      40903: inst = 32'h10408000;
      40904: inst = 32'hc405589;
      40905: inst = 32'h8220000;
      40906: inst = 32'h10408000;
      40907: inst = 32'hc40558a;
      40908: inst = 32'h8220000;
      40909: inst = 32'h10408000;
      40910: inst = 32'hc40558b;
      40911: inst = 32'h8220000;
      40912: inst = 32'h10408000;
      40913: inst = 32'hc40558c;
      40914: inst = 32'h8220000;
      40915: inst = 32'h10408000;
      40916: inst = 32'hc40558d;
      40917: inst = 32'h8220000;
      40918: inst = 32'h10408000;
      40919: inst = 32'hc40558e;
      40920: inst = 32'h8220000;
      40921: inst = 32'h10408000;
      40922: inst = 32'hc40558f;
      40923: inst = 32'h8220000;
      40924: inst = 32'h10408000;
      40925: inst = 32'hc405590;
      40926: inst = 32'h8220000;
      40927: inst = 32'h10408000;
      40928: inst = 32'hc405591;
      40929: inst = 32'h8220000;
      40930: inst = 32'h10408000;
      40931: inst = 32'hc40559c;
      40932: inst = 32'h8220000;
      40933: inst = 32'h10408000;
      40934: inst = 32'hc4055a3;
      40935: inst = 32'h8220000;
      40936: inst = 32'h10408000;
      40937: inst = 32'hc4055a4;
      40938: inst = 32'h8220000;
      40939: inst = 32'h10408000;
      40940: inst = 32'hc4055a5;
      40941: inst = 32'h8220000;
      40942: inst = 32'h10408000;
      40943: inst = 32'hc4055a6;
      40944: inst = 32'h8220000;
      40945: inst = 32'h10408000;
      40946: inst = 32'hc4055b0;
      40947: inst = 32'h8220000;
      40948: inst = 32'h10408000;
      40949: inst = 32'hc4055b1;
      40950: inst = 32'h8220000;
      40951: inst = 32'h10408000;
      40952: inst = 32'hc4055b2;
      40953: inst = 32'h8220000;
      40954: inst = 32'h10408000;
      40955: inst = 32'hc4055b3;
      40956: inst = 32'h8220000;
      40957: inst = 32'h10408000;
      40958: inst = 32'hc4055b4;
      40959: inst = 32'h8220000;
      40960: inst = 32'h10408000;
      40961: inst = 32'hc4055b5;
      40962: inst = 32'h8220000;
      40963: inst = 32'h10408000;
      40964: inst = 32'hc4055b9;
      40965: inst = 32'h8220000;
      40966: inst = 32'h10408000;
      40967: inst = 32'hc4055ba;
      40968: inst = 32'h8220000;
      40969: inst = 32'h10408000;
      40970: inst = 32'hc4055bb;
      40971: inst = 32'h8220000;
      40972: inst = 32'h10408000;
      40973: inst = 32'hc4055bc;
      40974: inst = 32'h8220000;
      40975: inst = 32'h10408000;
      40976: inst = 32'hc4055bd;
      40977: inst = 32'h8220000;
      40978: inst = 32'h10408000;
      40979: inst = 32'hc4055be;
      40980: inst = 32'h8220000;
      40981: inst = 32'h10408000;
      40982: inst = 32'hc4055bf;
      40983: inst = 32'h8220000;
      40984: inst = 32'h10408000;
      40985: inst = 32'hc4055c0;
      40986: inst = 32'h8220000;
      40987: inst = 32'h10408000;
      40988: inst = 32'hc4055c1;
      40989: inst = 32'h8220000;
      40990: inst = 32'h10408000;
      40991: inst = 32'hc4055c2;
      40992: inst = 32'h8220000;
      40993: inst = 32'h10408000;
      40994: inst = 32'hc4055c3;
      40995: inst = 32'h8220000;
      40996: inst = 32'h10408000;
      40997: inst = 32'hc4055c4;
      40998: inst = 32'h8220000;
      40999: inst = 32'h10408000;
      41000: inst = 32'hc4055c5;
      41001: inst = 32'h8220000;
      41002: inst = 32'h10408000;
      41003: inst = 32'hc4055c6;
      41004: inst = 32'h8220000;
      41005: inst = 32'h10408000;
      41006: inst = 32'hc4055c7;
      41007: inst = 32'h8220000;
      41008: inst = 32'h10408000;
      41009: inst = 32'hc4055c8;
      41010: inst = 32'h8220000;
      41011: inst = 32'h10408000;
      41012: inst = 32'hc4055c9;
      41013: inst = 32'h8220000;
      41014: inst = 32'h10408000;
      41015: inst = 32'hc4055ca;
      41016: inst = 32'h8220000;
      41017: inst = 32'h10408000;
      41018: inst = 32'hc4055cb;
      41019: inst = 32'h8220000;
      41020: inst = 32'h10408000;
      41021: inst = 32'hc4055cc;
      41022: inst = 32'h8220000;
      41023: inst = 32'h10408000;
      41024: inst = 32'hc4055cd;
      41025: inst = 32'h8220000;
      41026: inst = 32'h10408000;
      41027: inst = 32'hc4055ce;
      41028: inst = 32'h8220000;
      41029: inst = 32'h10408000;
      41030: inst = 32'hc4055cf;
      41031: inst = 32'h8220000;
      41032: inst = 32'h10408000;
      41033: inst = 32'hc4055d0;
      41034: inst = 32'h8220000;
      41035: inst = 32'h10408000;
      41036: inst = 32'hc4055d1;
      41037: inst = 32'h8220000;
      41038: inst = 32'h10408000;
      41039: inst = 32'hc4055d2;
      41040: inst = 32'h8220000;
      41041: inst = 32'h10408000;
      41042: inst = 32'hc4055d3;
      41043: inst = 32'h8220000;
      41044: inst = 32'h10408000;
      41045: inst = 32'hc4055d4;
      41046: inst = 32'h8220000;
      41047: inst = 32'h10408000;
      41048: inst = 32'hc4055d5;
      41049: inst = 32'h8220000;
      41050: inst = 32'h10408000;
      41051: inst = 32'hc4055d6;
      41052: inst = 32'h8220000;
      41053: inst = 32'h10408000;
      41054: inst = 32'hc4055d7;
      41055: inst = 32'h8220000;
      41056: inst = 32'h10408000;
      41057: inst = 32'hc4055d8;
      41058: inst = 32'h8220000;
      41059: inst = 32'h10408000;
      41060: inst = 32'hc4055d9;
      41061: inst = 32'h8220000;
      41062: inst = 32'h10408000;
      41063: inst = 32'hc4055da;
      41064: inst = 32'h8220000;
      41065: inst = 32'h10408000;
      41066: inst = 32'hc4055db;
      41067: inst = 32'h8220000;
      41068: inst = 32'h10408000;
      41069: inst = 32'hc4055dc;
      41070: inst = 32'h8220000;
      41071: inst = 32'h10408000;
      41072: inst = 32'hc4055dd;
      41073: inst = 32'h8220000;
      41074: inst = 32'h10408000;
      41075: inst = 32'hc4055de;
      41076: inst = 32'h8220000;
      41077: inst = 32'h10408000;
      41078: inst = 32'hc4055df;
      41079: inst = 32'h8220000;
      41080: inst = 32'h10408000;
      41081: inst = 32'hc4055e0;
      41082: inst = 32'h8220000;
      41083: inst = 32'h10408000;
      41084: inst = 32'hc4055e1;
      41085: inst = 32'h8220000;
      41086: inst = 32'h10408000;
      41087: inst = 32'hc4055e2;
      41088: inst = 32'h8220000;
      41089: inst = 32'h10408000;
      41090: inst = 32'hc4055e3;
      41091: inst = 32'h8220000;
      41092: inst = 32'h10408000;
      41093: inst = 32'hc4055e4;
      41094: inst = 32'h8220000;
      41095: inst = 32'h10408000;
      41096: inst = 32'hc4055e5;
      41097: inst = 32'h8220000;
      41098: inst = 32'h10408000;
      41099: inst = 32'hc4055e6;
      41100: inst = 32'h8220000;
      41101: inst = 32'h10408000;
      41102: inst = 32'hc4055e7;
      41103: inst = 32'h8220000;
      41104: inst = 32'h10408000;
      41105: inst = 32'hc4055e8;
      41106: inst = 32'h8220000;
      41107: inst = 32'h10408000;
      41108: inst = 32'hc4055e9;
      41109: inst = 32'h8220000;
      41110: inst = 32'h10408000;
      41111: inst = 32'hc4055ea;
      41112: inst = 32'h8220000;
      41113: inst = 32'h10408000;
      41114: inst = 32'hc4055eb;
      41115: inst = 32'h8220000;
      41116: inst = 32'h10408000;
      41117: inst = 32'hc4055ec;
      41118: inst = 32'h8220000;
      41119: inst = 32'h10408000;
      41120: inst = 32'hc4055ed;
      41121: inst = 32'h8220000;
      41122: inst = 32'h10408000;
      41123: inst = 32'hc4055ee;
      41124: inst = 32'h8220000;
      41125: inst = 32'h10408000;
      41126: inst = 32'hc4055ef;
      41127: inst = 32'h8220000;
      41128: inst = 32'h10408000;
      41129: inst = 32'hc4055f0;
      41130: inst = 32'h8220000;
      41131: inst = 32'h10408000;
      41132: inst = 32'hc4055f1;
      41133: inst = 32'h8220000;
      41134: inst = 32'h10408000;
      41135: inst = 32'hc4055fc;
      41136: inst = 32'h8220000;
      41137: inst = 32'h10408000;
      41138: inst = 32'hc405603;
      41139: inst = 32'h8220000;
      41140: inst = 32'h10408000;
      41141: inst = 32'hc405604;
      41142: inst = 32'h8220000;
      41143: inst = 32'h10408000;
      41144: inst = 32'hc405605;
      41145: inst = 32'h8220000;
      41146: inst = 32'h10408000;
      41147: inst = 32'hc405606;
      41148: inst = 32'h8220000;
      41149: inst = 32'h10408000;
      41150: inst = 32'hc405613;
      41151: inst = 32'h8220000;
      41152: inst = 32'h10408000;
      41153: inst = 32'hc405614;
      41154: inst = 32'h8220000;
      41155: inst = 32'h10408000;
      41156: inst = 32'hc405615;
      41157: inst = 32'h8220000;
      41158: inst = 32'h10408000;
      41159: inst = 32'hc405619;
      41160: inst = 32'h8220000;
      41161: inst = 32'h10408000;
      41162: inst = 32'hc40561a;
      41163: inst = 32'h8220000;
      41164: inst = 32'h10408000;
      41165: inst = 32'hc40561b;
      41166: inst = 32'h8220000;
      41167: inst = 32'h10408000;
      41168: inst = 32'hc40561c;
      41169: inst = 32'h8220000;
      41170: inst = 32'h10408000;
      41171: inst = 32'hc40561d;
      41172: inst = 32'h8220000;
      41173: inst = 32'h10408000;
      41174: inst = 32'hc40561e;
      41175: inst = 32'h8220000;
      41176: inst = 32'h10408000;
      41177: inst = 32'hc40561f;
      41178: inst = 32'h8220000;
      41179: inst = 32'h10408000;
      41180: inst = 32'hc405620;
      41181: inst = 32'h8220000;
      41182: inst = 32'h10408000;
      41183: inst = 32'hc405621;
      41184: inst = 32'h8220000;
      41185: inst = 32'h10408000;
      41186: inst = 32'hc405622;
      41187: inst = 32'h8220000;
      41188: inst = 32'h10408000;
      41189: inst = 32'hc405623;
      41190: inst = 32'h8220000;
      41191: inst = 32'h10408000;
      41192: inst = 32'hc405624;
      41193: inst = 32'h8220000;
      41194: inst = 32'h10408000;
      41195: inst = 32'hc405625;
      41196: inst = 32'h8220000;
      41197: inst = 32'h10408000;
      41198: inst = 32'hc405626;
      41199: inst = 32'h8220000;
      41200: inst = 32'h10408000;
      41201: inst = 32'hc405627;
      41202: inst = 32'h8220000;
      41203: inst = 32'h10408000;
      41204: inst = 32'hc405628;
      41205: inst = 32'h8220000;
      41206: inst = 32'h10408000;
      41207: inst = 32'hc405629;
      41208: inst = 32'h8220000;
      41209: inst = 32'h10408000;
      41210: inst = 32'hc40562a;
      41211: inst = 32'h8220000;
      41212: inst = 32'h10408000;
      41213: inst = 32'hc40562b;
      41214: inst = 32'h8220000;
      41215: inst = 32'h10408000;
      41216: inst = 32'hc40562c;
      41217: inst = 32'h8220000;
      41218: inst = 32'h10408000;
      41219: inst = 32'hc40562d;
      41220: inst = 32'h8220000;
      41221: inst = 32'h10408000;
      41222: inst = 32'hc40562e;
      41223: inst = 32'h8220000;
      41224: inst = 32'h10408000;
      41225: inst = 32'hc40562f;
      41226: inst = 32'h8220000;
      41227: inst = 32'h10408000;
      41228: inst = 32'hc405630;
      41229: inst = 32'h8220000;
      41230: inst = 32'h10408000;
      41231: inst = 32'hc405631;
      41232: inst = 32'h8220000;
      41233: inst = 32'h10408000;
      41234: inst = 32'hc405632;
      41235: inst = 32'h8220000;
      41236: inst = 32'h10408000;
      41237: inst = 32'hc405633;
      41238: inst = 32'h8220000;
      41239: inst = 32'h10408000;
      41240: inst = 32'hc405634;
      41241: inst = 32'h8220000;
      41242: inst = 32'h10408000;
      41243: inst = 32'hc405635;
      41244: inst = 32'h8220000;
      41245: inst = 32'h10408000;
      41246: inst = 32'hc405636;
      41247: inst = 32'h8220000;
      41248: inst = 32'h10408000;
      41249: inst = 32'hc405637;
      41250: inst = 32'h8220000;
      41251: inst = 32'h10408000;
      41252: inst = 32'hc405638;
      41253: inst = 32'h8220000;
      41254: inst = 32'h10408000;
      41255: inst = 32'hc405639;
      41256: inst = 32'h8220000;
      41257: inst = 32'h10408000;
      41258: inst = 32'hc40563a;
      41259: inst = 32'h8220000;
      41260: inst = 32'h10408000;
      41261: inst = 32'hc40563b;
      41262: inst = 32'h8220000;
      41263: inst = 32'h10408000;
      41264: inst = 32'hc40563c;
      41265: inst = 32'h8220000;
      41266: inst = 32'h10408000;
      41267: inst = 32'hc40563d;
      41268: inst = 32'h8220000;
      41269: inst = 32'h10408000;
      41270: inst = 32'hc40563e;
      41271: inst = 32'h8220000;
      41272: inst = 32'h10408000;
      41273: inst = 32'hc40563f;
      41274: inst = 32'h8220000;
      41275: inst = 32'h10408000;
      41276: inst = 32'hc405640;
      41277: inst = 32'h8220000;
      41278: inst = 32'h10408000;
      41279: inst = 32'hc405641;
      41280: inst = 32'h8220000;
      41281: inst = 32'h10408000;
      41282: inst = 32'hc405642;
      41283: inst = 32'h8220000;
      41284: inst = 32'h10408000;
      41285: inst = 32'hc405643;
      41286: inst = 32'h8220000;
      41287: inst = 32'h10408000;
      41288: inst = 32'hc405644;
      41289: inst = 32'h8220000;
      41290: inst = 32'h10408000;
      41291: inst = 32'hc405645;
      41292: inst = 32'h8220000;
      41293: inst = 32'h10408000;
      41294: inst = 32'hc405646;
      41295: inst = 32'h8220000;
      41296: inst = 32'h10408000;
      41297: inst = 32'hc405647;
      41298: inst = 32'h8220000;
      41299: inst = 32'h10408000;
      41300: inst = 32'hc405648;
      41301: inst = 32'h8220000;
      41302: inst = 32'h10408000;
      41303: inst = 32'hc405649;
      41304: inst = 32'h8220000;
      41305: inst = 32'h10408000;
      41306: inst = 32'hc40564a;
      41307: inst = 32'h8220000;
      41308: inst = 32'h10408000;
      41309: inst = 32'hc40564b;
      41310: inst = 32'h8220000;
      41311: inst = 32'h10408000;
      41312: inst = 32'hc40564c;
      41313: inst = 32'h8220000;
      41314: inst = 32'h10408000;
      41315: inst = 32'hc40564d;
      41316: inst = 32'h8220000;
      41317: inst = 32'h10408000;
      41318: inst = 32'hc40564e;
      41319: inst = 32'h8220000;
      41320: inst = 32'h10408000;
      41321: inst = 32'hc40564f;
      41322: inst = 32'h8220000;
      41323: inst = 32'h10408000;
      41324: inst = 32'hc405650;
      41325: inst = 32'h8220000;
      41326: inst = 32'h10408000;
      41327: inst = 32'hc405651;
      41328: inst = 32'h8220000;
      41329: inst = 32'h10408000;
      41330: inst = 32'hc40565c;
      41331: inst = 32'h8220000;
      41332: inst = 32'h10408000;
      41333: inst = 32'hc405663;
      41334: inst = 32'h8220000;
      41335: inst = 32'h10408000;
      41336: inst = 32'hc405664;
      41337: inst = 32'h8220000;
      41338: inst = 32'h10408000;
      41339: inst = 32'hc405665;
      41340: inst = 32'h8220000;
      41341: inst = 32'h10408000;
      41342: inst = 32'hc405666;
      41343: inst = 32'h8220000;
      41344: inst = 32'h10408000;
      41345: inst = 32'hc405667;
      41346: inst = 32'h8220000;
      41347: inst = 32'h10408000;
      41348: inst = 32'hc405674;
      41349: inst = 32'h8220000;
      41350: inst = 32'h10408000;
      41351: inst = 32'hc405675;
      41352: inst = 32'h8220000;
      41353: inst = 32'h10408000;
      41354: inst = 32'hc405679;
      41355: inst = 32'h8220000;
      41356: inst = 32'h10408000;
      41357: inst = 32'hc40567a;
      41358: inst = 32'h8220000;
      41359: inst = 32'h10408000;
      41360: inst = 32'hc40567b;
      41361: inst = 32'h8220000;
      41362: inst = 32'h10408000;
      41363: inst = 32'hc40567c;
      41364: inst = 32'h8220000;
      41365: inst = 32'h10408000;
      41366: inst = 32'hc40567d;
      41367: inst = 32'h8220000;
      41368: inst = 32'h10408000;
      41369: inst = 32'hc40567e;
      41370: inst = 32'h8220000;
      41371: inst = 32'h10408000;
      41372: inst = 32'hc40567f;
      41373: inst = 32'h8220000;
      41374: inst = 32'h10408000;
      41375: inst = 32'hc405680;
      41376: inst = 32'h8220000;
      41377: inst = 32'h10408000;
      41378: inst = 32'hc405681;
      41379: inst = 32'h8220000;
      41380: inst = 32'h10408000;
      41381: inst = 32'hc405682;
      41382: inst = 32'h8220000;
      41383: inst = 32'h10408000;
      41384: inst = 32'hc405683;
      41385: inst = 32'h8220000;
      41386: inst = 32'h10408000;
      41387: inst = 32'hc405684;
      41388: inst = 32'h8220000;
      41389: inst = 32'h10408000;
      41390: inst = 32'hc405685;
      41391: inst = 32'h8220000;
      41392: inst = 32'h10408000;
      41393: inst = 32'hc405686;
      41394: inst = 32'h8220000;
      41395: inst = 32'h10408000;
      41396: inst = 32'hc405687;
      41397: inst = 32'h8220000;
      41398: inst = 32'h10408000;
      41399: inst = 32'hc405688;
      41400: inst = 32'h8220000;
      41401: inst = 32'h10408000;
      41402: inst = 32'hc405689;
      41403: inst = 32'h8220000;
      41404: inst = 32'h10408000;
      41405: inst = 32'hc40568a;
      41406: inst = 32'h8220000;
      41407: inst = 32'h10408000;
      41408: inst = 32'hc40568b;
      41409: inst = 32'h8220000;
      41410: inst = 32'h10408000;
      41411: inst = 32'hc40568c;
      41412: inst = 32'h8220000;
      41413: inst = 32'h10408000;
      41414: inst = 32'hc40568d;
      41415: inst = 32'h8220000;
      41416: inst = 32'h10408000;
      41417: inst = 32'hc40568e;
      41418: inst = 32'h8220000;
      41419: inst = 32'h10408000;
      41420: inst = 32'hc40568f;
      41421: inst = 32'h8220000;
      41422: inst = 32'h10408000;
      41423: inst = 32'hc405690;
      41424: inst = 32'h8220000;
      41425: inst = 32'h10408000;
      41426: inst = 32'hc405691;
      41427: inst = 32'h8220000;
      41428: inst = 32'h10408000;
      41429: inst = 32'hc405692;
      41430: inst = 32'h8220000;
      41431: inst = 32'h10408000;
      41432: inst = 32'hc405693;
      41433: inst = 32'h8220000;
      41434: inst = 32'h10408000;
      41435: inst = 32'hc405694;
      41436: inst = 32'h8220000;
      41437: inst = 32'h10408000;
      41438: inst = 32'hc405695;
      41439: inst = 32'h8220000;
      41440: inst = 32'h10408000;
      41441: inst = 32'hc405696;
      41442: inst = 32'h8220000;
      41443: inst = 32'h10408000;
      41444: inst = 32'hc405697;
      41445: inst = 32'h8220000;
      41446: inst = 32'h10408000;
      41447: inst = 32'hc405698;
      41448: inst = 32'h8220000;
      41449: inst = 32'h10408000;
      41450: inst = 32'hc405699;
      41451: inst = 32'h8220000;
      41452: inst = 32'h10408000;
      41453: inst = 32'hc40569a;
      41454: inst = 32'h8220000;
      41455: inst = 32'h10408000;
      41456: inst = 32'hc40569b;
      41457: inst = 32'h8220000;
      41458: inst = 32'h10408000;
      41459: inst = 32'hc40569c;
      41460: inst = 32'h8220000;
      41461: inst = 32'h10408000;
      41462: inst = 32'hc40569d;
      41463: inst = 32'h8220000;
      41464: inst = 32'h10408000;
      41465: inst = 32'hc40569e;
      41466: inst = 32'h8220000;
      41467: inst = 32'h10408000;
      41468: inst = 32'hc40569f;
      41469: inst = 32'h8220000;
      41470: inst = 32'h10408000;
      41471: inst = 32'hc4056a0;
      41472: inst = 32'h8220000;
      41473: inst = 32'h10408000;
      41474: inst = 32'hc4056a1;
      41475: inst = 32'h8220000;
      41476: inst = 32'h10408000;
      41477: inst = 32'hc4056a2;
      41478: inst = 32'h8220000;
      41479: inst = 32'h10408000;
      41480: inst = 32'hc4056a3;
      41481: inst = 32'h8220000;
      41482: inst = 32'h10408000;
      41483: inst = 32'hc4056a4;
      41484: inst = 32'h8220000;
      41485: inst = 32'h10408000;
      41486: inst = 32'hc4056a5;
      41487: inst = 32'h8220000;
      41488: inst = 32'h10408000;
      41489: inst = 32'hc4056a6;
      41490: inst = 32'h8220000;
      41491: inst = 32'h10408000;
      41492: inst = 32'hc4056a7;
      41493: inst = 32'h8220000;
      41494: inst = 32'h10408000;
      41495: inst = 32'hc4056a8;
      41496: inst = 32'h8220000;
      41497: inst = 32'h10408000;
      41498: inst = 32'hc4056a9;
      41499: inst = 32'h8220000;
      41500: inst = 32'h10408000;
      41501: inst = 32'hc4056aa;
      41502: inst = 32'h8220000;
      41503: inst = 32'h10408000;
      41504: inst = 32'hc4056ab;
      41505: inst = 32'h8220000;
      41506: inst = 32'h10408000;
      41507: inst = 32'hc4056ac;
      41508: inst = 32'h8220000;
      41509: inst = 32'h10408000;
      41510: inst = 32'hc4056ad;
      41511: inst = 32'h8220000;
      41512: inst = 32'h10408000;
      41513: inst = 32'hc4056ae;
      41514: inst = 32'h8220000;
      41515: inst = 32'h10408000;
      41516: inst = 32'hc4056af;
      41517: inst = 32'h8220000;
      41518: inst = 32'h10408000;
      41519: inst = 32'hc4056b0;
      41520: inst = 32'h8220000;
      41521: inst = 32'h10408000;
      41522: inst = 32'hc4056b1;
      41523: inst = 32'h8220000;
      41524: inst = 32'h10408000;
      41525: inst = 32'hc4056bc;
      41526: inst = 32'h8220000;
      41527: inst = 32'h10408000;
      41528: inst = 32'hc405711;
      41529: inst = 32'h8220000;
      41530: inst = 32'h10408000;
      41531: inst = 32'hc40571c;
      41532: inst = 32'h8220000;
      41533: inst = 32'h10408000;
      41534: inst = 32'hc405771;
      41535: inst = 32'h8220000;
      41536: inst = 32'h10408000;
      41537: inst = 32'hc40577c;
      41538: inst = 32'h8220000;
      41539: inst = 32'h10408000;
      41540: inst = 32'hc4057d1;
      41541: inst = 32'h8220000;
      41542: inst = 32'h10408000;
      41543: inst = 32'hc4057dc;
      41544: inst = 32'h8220000;
      41545: inst = 32'hc20cba6;
      41546: inst = 32'h10408000;
      41547: inst = 32'hc403fe4;
      41548: inst = 32'h8220000;
      41549: inst = 32'h10408000;
      41550: inst = 32'hc403fec;
      41551: inst = 32'h8220000;
      41552: inst = 32'h10408000;
      41553: inst = 32'hc4040ac;
      41554: inst = 32'h8220000;
      41555: inst = 32'h10408000;
      41556: inst = 32'hc40410c;
      41557: inst = 32'h8220000;
      41558: inst = 32'h10408000;
      41559: inst = 32'hc40416c;
      41560: inst = 32'h8220000;
      41561: inst = 32'h10408000;
      41562: inst = 32'hc4041c4;
      41563: inst = 32'h8220000;
      41564: inst = 32'h10408000;
      41565: inst = 32'hc404224;
      41566: inst = 32'h8220000;
      41567: inst = 32'h10408000;
      41568: inst = 32'hc404284;
      41569: inst = 32'h8220000;
      41570: inst = 32'h10408000;
      41571: inst = 32'hc40428c;
      41572: inst = 32'h8220000;
      41573: inst = 32'h10408000;
      41574: inst = 32'hc4042e4;
      41575: inst = 32'h8220000;
      41576: inst = 32'h10408000;
      41577: inst = 32'hc4042ec;
      41578: inst = 32'h8220000;
      41579: inst = 32'h10408000;
      41580: inst = 32'hc404344;
      41581: inst = 32'h8220000;
      41582: inst = 32'h10408000;
      41583: inst = 32'hc40434c;
      41584: inst = 32'h8220000;
      41585: inst = 32'h10408000;
      41586: inst = 32'hc4054d2;
      41587: inst = 32'h8220000;
      41588: inst = 32'hc20cb44;
      41589: inst = 32'h10408000;
      41590: inst = 32'hc403fe5;
      41591: inst = 32'h8220000;
      41592: inst = 32'h10408000;
      41593: inst = 32'hc403fe6;
      41594: inst = 32'h8220000;
      41595: inst = 32'h10408000;
      41596: inst = 32'hc403fe7;
      41597: inst = 32'h8220000;
      41598: inst = 32'h10408000;
      41599: inst = 32'hc403fe8;
      41600: inst = 32'h8220000;
      41601: inst = 32'h10408000;
      41602: inst = 32'hc403fe9;
      41603: inst = 32'h8220000;
      41604: inst = 32'h10408000;
      41605: inst = 32'hc403fea;
      41606: inst = 32'h8220000;
      41607: inst = 32'h10408000;
      41608: inst = 32'hc403feb;
      41609: inst = 32'h8220000;
      41610: inst = 32'h10408000;
      41611: inst = 32'hc404104;
      41612: inst = 32'h8220000;
      41613: inst = 32'h10408000;
      41614: inst = 32'hc4043a6;
      41615: inst = 32'h8220000;
      41616: inst = 32'h10408000;
      41617: inst = 32'hc4043a7;
      41618: inst = 32'h8220000;
      41619: inst = 32'h10408000;
      41620: inst = 32'hc4043a8;
      41621: inst = 32'h8220000;
      41622: inst = 32'h10408000;
      41623: inst = 32'hc4043a9;
      41624: inst = 32'h8220000;
      41625: inst = 32'h10408000;
      41626: inst = 32'hc4043aa;
      41627: inst = 32'h8220000;
      41628: inst = 32'h10408000;
      41629: inst = 32'hc4043ab;
      41630: inst = 32'h8220000;
      41631: inst = 32'h10408000;
      41632: inst = 32'hc405354;
      41633: inst = 32'h8220000;
      41634: inst = 32'h10408000;
      41635: inst = 32'hc4053b2;
      41636: inst = 32'h8220000;
      41637: inst = 32'h10408000;
      41638: inst = 32'hc405532;
      41639: inst = 32'h8220000;
      41640: inst = 32'hc20a5f0;
      41641: inst = 32'h10408000;
      41642: inst = 32'hc403fed;
      41643: inst = 32'h8220000;
      41644: inst = 32'hc203d29;
      41645: inst = 32'h10408000;
      41646: inst = 32'hc403fee;
      41647: inst = 32'h8220000;
      41648: inst = 32'hc203ca9;
      41649: inst = 32'h10408000;
      41650: inst = 32'hc403fef;
      41651: inst = 32'h8220000;
      41652: inst = 32'hc20448a;
      41653: inst = 32'h10408000;
      41654: inst = 32'hc403ff0;
      41655: inst = 32'h8220000;
      41656: inst = 32'hc20636f;
      41657: inst = 32'h10408000;
      41658: inst = 32'hc403ff1;
      41659: inst = 32'h8220000;
      41660: inst = 32'h10408000;
      41661: inst = 32'hc403ff7;
      41662: inst = 32'h8220000;
      41663: inst = 32'h10408000;
      41664: inst = 32'hc404053;
      41665: inst = 32'h8220000;
      41666: inst = 32'h10408000;
      41667: inst = 32'hc404675;
      41668: inst = 32'h8220000;
      41669: inst = 32'h10408000;
      41670: inst = 32'hc404677;
      41671: inst = 32'h8220000;
      41672: inst = 32'h10408000;
      41673: inst = 32'hc4046ca;
      41674: inst = 32'h8220000;
      41675: inst = 32'h10408000;
      41676: inst = 32'hc4046d5;
      41677: inst = 32'h8220000;
      41678: inst = 32'h10408000;
      41679: inst = 32'hc404732;
      41680: inst = 32'h8220000;
      41681: inst = 32'hc2053ac;
      41682: inst = 32'h10408000;
      41683: inst = 32'hc403ff2;
      41684: inst = 32'h8220000;
      41685: inst = 32'hc203427;
      41686: inst = 32'h10408000;
      41687: inst = 32'hc403ff3;
      41688: inst = 32'h8220000;
      41689: inst = 32'hc20638f;
      41690: inst = 32'h10408000;
      41691: inst = 32'hc403ff4;
      41692: inst = 32'h8220000;
      41693: inst = 32'hc204bac;
      41694: inst = 32'h10408000;
      41695: inst = 32'hc403ff6;
      41696: inst = 32'h8220000;
      41697: inst = 32'h10408000;
      41698: inst = 32'hc40404e;
      41699: inst = 32'h8220000;
      41700: inst = 32'hc204549;
      41701: inst = 32'h10408000;
      41702: inst = 32'hc403ffa;
      41703: inst = 32'h8220000;
      41704: inst = 32'hc20546c;
      41705: inst = 32'h10408000;
      41706: inst = 32'hc403ffb;
      41707: inst = 32'h8220000;
      41708: inst = 32'hc20544d;
      41709: inst = 32'h10408000;
      41710: inst = 32'hc403ffc;
      41711: inst = 32'h8220000;
      41712: inst = 32'hc20cb86;
      41713: inst = 32'h10408000;
      41714: inst = 32'hc404044;
      41715: inst = 32'h8220000;
      41716: inst = 32'hc20dba5;
      41717: inst = 32'h10408000;
      41718: inst = 32'hc404045;
      41719: inst = 32'h8220000;
      41720: inst = 32'h10408000;
      41721: inst = 32'hc4041c6;
      41722: inst = 32'h8220000;
      41723: inst = 32'h10408000;
      41724: inst = 32'hc4041c7;
      41725: inst = 32'h8220000;
      41726: inst = 32'h10408000;
      41727: inst = 32'hc40428a;
      41728: inst = 32'h8220000;
      41729: inst = 32'h10408000;
      41730: inst = 32'hc404345;
      41731: inst = 32'h8220000;
      41732: inst = 32'h10408000;
      41733: inst = 32'hc4053b4;
      41734: inst = 32'h8220000;
      41735: inst = 32'h10408000;
      41736: inst = 32'hc405713;
      41737: inst = 32'h8220000;
      41738: inst = 32'hc20dbc5;
      41739: inst = 32'h10408000;
      41740: inst = 32'hc404046;
      41741: inst = 32'h8220000;
      41742: inst = 32'h10408000;
      41743: inst = 32'hc404047;
      41744: inst = 32'h8220000;
      41745: inst = 32'h10408000;
      41746: inst = 32'hc4040a9;
      41747: inst = 32'h8220000;
      41748: inst = 32'h10408000;
      41749: inst = 32'hc4040aa;
      41750: inst = 32'h8220000;
      41751: inst = 32'h10408000;
      41752: inst = 32'hc4040ab;
      41753: inst = 32'h8220000;
      41754: inst = 32'h10408000;
      41755: inst = 32'hc404109;
      41756: inst = 32'h8220000;
      41757: inst = 32'h10408000;
      41758: inst = 32'hc40410a;
      41759: inst = 32'h8220000;
      41760: inst = 32'h10408000;
      41761: inst = 32'hc40410b;
      41762: inst = 32'h8220000;
      41763: inst = 32'h10408000;
      41764: inst = 32'hc404169;
      41765: inst = 32'h8220000;
      41766: inst = 32'h10408000;
      41767: inst = 32'hc4041c8;
      41768: inst = 32'h8220000;
      41769: inst = 32'h10408000;
      41770: inst = 32'hc4041c9;
      41771: inst = 32'h8220000;
      41772: inst = 32'h10408000;
      41773: inst = 32'hc404226;
      41774: inst = 32'h8220000;
      41775: inst = 32'h10408000;
      41776: inst = 32'hc404227;
      41777: inst = 32'h8220000;
      41778: inst = 32'h10408000;
      41779: inst = 32'hc404228;
      41780: inst = 32'h8220000;
      41781: inst = 32'h10408000;
      41782: inst = 32'hc404286;
      41783: inst = 32'h8220000;
      41784: inst = 32'h10408000;
      41785: inst = 32'hc404287;
      41786: inst = 32'h8220000;
      41787: inst = 32'h10408000;
      41788: inst = 32'hc404288;
      41789: inst = 32'h8220000;
      41790: inst = 32'h10408000;
      41791: inst = 32'hc404289;
      41792: inst = 32'h8220000;
      41793: inst = 32'h10408000;
      41794: inst = 32'hc4042e6;
      41795: inst = 32'h8220000;
      41796: inst = 32'h10408000;
      41797: inst = 32'hc4042e7;
      41798: inst = 32'h8220000;
      41799: inst = 32'h10408000;
      41800: inst = 32'hc4042e8;
      41801: inst = 32'h8220000;
      41802: inst = 32'h10408000;
      41803: inst = 32'hc4042e9;
      41804: inst = 32'h8220000;
      41805: inst = 32'h10408000;
      41806: inst = 32'hc4042ea;
      41807: inst = 32'h8220000;
      41808: inst = 32'h10408000;
      41809: inst = 32'hc4042eb;
      41810: inst = 32'h8220000;
      41811: inst = 32'h10408000;
      41812: inst = 32'hc405594;
      41813: inst = 32'h8220000;
      41814: inst = 32'h10408000;
      41815: inst = 32'hc4055f4;
      41816: inst = 32'h8220000;
      41817: inst = 32'h10408000;
      41818: inst = 32'hc405653;
      41819: inst = 32'h8220000;
      41820: inst = 32'hc20dbc6;
      41821: inst = 32'h10408000;
      41822: inst = 32'hc404048;
      41823: inst = 32'h8220000;
      41824: inst = 32'h10408000;
      41825: inst = 32'hc404049;
      41826: inst = 32'h8220000;
      41827: inst = 32'h10408000;
      41828: inst = 32'hc40404a;
      41829: inst = 32'h8220000;
      41830: inst = 32'h10408000;
      41831: inst = 32'hc404229;
      41832: inst = 32'h8220000;
      41833: inst = 32'h10408000;
      41834: inst = 32'hc404347;
      41835: inst = 32'h8220000;
      41836: inst = 32'h10408000;
      41837: inst = 32'hc404348;
      41838: inst = 32'h8220000;
      41839: inst = 32'h10408000;
      41840: inst = 32'hc404349;
      41841: inst = 32'h8220000;
      41842: inst = 32'h10408000;
      41843: inst = 32'hc40434a;
      41844: inst = 32'h8220000;
      41845: inst = 32'h10408000;
      41846: inst = 32'hc4055f3;
      41847: inst = 32'h8220000;
      41848: inst = 32'hc20e3c6;
      41849: inst = 32'h10408000;
      41850: inst = 32'hc40404b;
      41851: inst = 32'h8220000;
      41852: inst = 32'h10408000;
      41853: inst = 32'hc404346;
      41854: inst = 32'h8220000;
      41855: inst = 32'h10408000;
      41856: inst = 32'hc40434b;
      41857: inst = 32'h8220000;
      41858: inst = 32'h10408000;
      41859: inst = 32'hc405654;
      41860: inst = 32'h8220000;
      41861: inst = 32'hc20cb85;
      41862: inst = 32'h10408000;
      41863: inst = 32'hc40404c;
      41864: inst = 32'h8220000;
      41865: inst = 32'hc206d0b;
      41866: inst = 32'h10408000;
      41867: inst = 32'hc40404d;
      41868: inst = 32'h8220000;
      41869: inst = 32'hc205c2d;
      41870: inst = 32'h10408000;
      41871: inst = 32'hc40404f;
      41872: inst = 32'h8220000;
      41873: inst = 32'hc203d88;
      41874: inst = 32'h10408000;
      41875: inst = 32'hc404050;
      41876: inst = 32'h8220000;
      41877: inst = 32'hc206b6f;
      41878: inst = 32'h10408000;
      41879: inst = 32'hc404051;
      41880: inst = 32'h8220000;
      41881: inst = 32'h10408000;
      41882: inst = 32'hc40466d;
      41883: inst = 32'h8220000;
      41884: inst = 32'h10408000;
      41885: inst = 32'hc4046d7;
      41886: inst = 32'h8220000;
      41887: inst = 32'h10408000;
      41888: inst = 32'hc40472e;
      41889: inst = 32'h8220000;
      41890: inst = 32'hc206b4f;
      41891: inst = 32'h10408000;
      41892: inst = 32'hc404052;
      41893: inst = 32'h8220000;
      41894: inst = 32'h10408000;
      41895: inst = 32'hc4056b6;
      41896: inst = 32'h8220000;
      41897: inst = 32'hc20542d;
      41898: inst = 32'h10408000;
      41899: inst = 32'hc404055;
      41900: inst = 32'h8220000;
      41901: inst = 32'h10408000;
      41902: inst = 32'hc4040b1;
      41903: inst = 32'h8220000;
      41904: inst = 32'hc205bee;
      41905: inst = 32'h10408000;
      41906: inst = 32'hc404056;
      41907: inst = 32'h8220000;
      41908: inst = 32'h10408000;
      41909: inst = 32'hc4040b5;
      41910: inst = 32'h8220000;
      41911: inst = 32'hc2063af;
      41912: inst = 32'h10408000;
      41913: inst = 32'hc404059;
      41914: inst = 32'h8220000;
      41915: inst = 32'hc203d49;
      41916: inst = 32'h10408000;
      41917: inst = 32'hc40405a;
      41918: inst = 32'h8220000;
      41919: inst = 32'hc206b70;
      41920: inst = 32'h10408000;
      41921: inst = 32'hc40405b;
      41922: inst = 32'h8220000;
      41923: inst = 32'h10408000;
      41924: inst = 32'hc404679;
      41925: inst = 32'h8220000;
      41926: inst = 32'h10408000;
      41927: inst = 32'hc40472d;
      41928: inst = 32'h8220000;
      41929: inst = 32'h10408000;
      41930: inst = 32'hc404730;
      41931: inst = 32'h8220000;
      41932: inst = 32'hc20cb64;
      41933: inst = 32'h10408000;
      41934: inst = 32'hc4040a4;
      41935: inst = 32'h8220000;
      41936: inst = 32'h10408000;
      41937: inst = 32'hc404164;
      41938: inst = 32'h8220000;
      41939: inst = 32'hc20dc08;
      41940: inst = 32'h10408000;
      41941: inst = 32'hc4040a5;
      41942: inst = 32'h8220000;
      41943: inst = 32'hc20f77b;
      41944: inst = 32'h10408000;
      41945: inst = 32'hc4040a6;
      41946: inst = 32'h8220000;
      41947: inst = 32'h10408000;
      41948: inst = 32'hc404154;
      41949: inst = 32'h8220000;
      41950: inst = 32'h10408000;
      41951: inst = 32'hc404155;
      41952: inst = 32'h8220000;
      41953: inst = 32'h10408000;
      41954: inst = 32'hc4041b0;
      41955: inst = 32'h8220000;
      41956: inst = 32'h10408000;
      41957: inst = 32'hc4041b7;
      41958: inst = 32'h8220000;
      41959: inst = 32'h10408000;
      41960: inst = 32'hc404274;
      41961: inst = 32'h8220000;
      41962: inst = 32'h10408000;
      41963: inst = 32'hc40427a;
      41964: inst = 32'h8220000;
      41965: inst = 32'h10408000;
      41966: inst = 32'hc404339;
      41967: inst = 32'h8220000;
      41968: inst = 32'h10408000;
      41969: inst = 32'hc4043fa;
      41970: inst = 32'h8220000;
      41971: inst = 32'h10408000;
      41972: inst = 32'hc404453;
      41973: inst = 32'h8220000;
      41974: inst = 32'h10408000;
      41975: inst = 32'hc404458;
      41976: inst = 32'h8220000;
      41977: inst = 32'h10408000;
      41978: inst = 32'hc4044b6;
      41979: inst = 32'h8220000;
      41980: inst = 32'h10408000;
      41981: inst = 32'hc4044ba;
      41982: inst = 32'h8220000;
      41983: inst = 32'h10408000;
      41984: inst = 32'hc404519;
      41985: inst = 32'h8220000;
      41986: inst = 32'h10408000;
      41987: inst = 32'hc4045d3;
      41988: inst = 32'h8220000;
      41989: inst = 32'hc20e48a;
      41990: inst = 32'h10408000;
      41991: inst = 32'hc4040a7;
      41992: inst = 32'h8220000;
      41993: inst = 32'hc20db84;
      41994: inst = 32'h10408000;
      41995: inst = 32'hc4040a8;
      41996: inst = 32'h8220000;
      41997: inst = 32'h10408000;
      41998: inst = 32'hc404108;
      41999: inst = 32'h8220000;
      42000: inst = 32'h10408000;
      42001: inst = 32'hc404168;
      42002: inst = 32'h8220000;
      42003: inst = 32'hc20a5d0;
      42004: inst = 32'h10408000;
      42005: inst = 32'hc4040ad;
      42006: inst = 32'h8220000;
      42007: inst = 32'h10408000;
      42008: inst = 32'hc404231;
      42009: inst = 32'h8220000;
      42010: inst = 32'h10408000;
      42011: inst = 32'hc404290;
      42012: inst = 32'h8220000;
      42013: inst = 32'hc205b6e;
      42014: inst = 32'h10408000;
      42015: inst = 32'hc4040ae;
      42016: inst = 32'h8220000;
      42017: inst = 32'hc204ccb;
      42018: inst = 32'h10408000;
      42019: inst = 32'hc4040b0;
      42020: inst = 32'h8220000;
      42021: inst = 32'h10408000;
      42022: inst = 32'hc4040ba;
      42023: inst = 32'h8220000;
      42024: inst = 32'hc2043aa;
      42025: inst = 32'h10408000;
      42026: inst = 32'hc4040b3;
      42027: inst = 32'h8220000;
      42028: inst = 32'h10408000;
      42029: inst = 32'hc4040b4;
      42030: inst = 32'h8220000;
      42031: inst = 32'hc2063ae;
      42032: inst = 32'h10408000;
      42033: inst = 32'hc4040b6;
      42034: inst = 32'h8220000;
      42035: inst = 32'h10408000;
      42036: inst = 32'hc40466a;
      42037: inst = 32'h8220000;
      42038: inst = 32'h10408000;
      42039: inst = 32'hc4046cd;
      42040: inst = 32'h8220000;
      42041: inst = 32'hc20544c;
      42042: inst = 32'h10408000;
      42043: inst = 32'hc4040b9;
      42044: inst = 32'h8220000;
      42045: inst = 32'h10408000;
      42046: inst = 32'hc4046cc;
      42047: inst = 32'h8220000;
      42048: inst = 32'h10408000;
      42049: inst = 32'hc40472b;
      42050: inst = 32'h8220000;
      42051: inst = 32'hc20dc28;
      42052: inst = 32'h10408000;
      42053: inst = 32'hc404105;
      42054: inst = 32'h8220000;
      42055: inst = 32'h10408000;
      42056: inst = 32'hc405533;
      42057: inst = 32'h8220000;
      42058: inst = 32'hc20ffff;
      42059: inst = 32'h10408000;
      42060: inst = 32'hc404106;
      42061: inst = 32'h8220000;
      42062: inst = 32'h10408000;
      42063: inst = 32'hc40439b;
      42064: inst = 32'h8220000;
      42065: inst = 32'h10408000;
      42066: inst = 32'hc404515;
      42067: inst = 32'h8220000;
      42068: inst = 32'hc20e4cc;
      42069: inst = 32'h10408000;
      42070: inst = 32'hc404107;
      42071: inst = 32'h8220000;
      42072: inst = 32'h10408000;
      42073: inst = 32'hc404167;
      42074: inst = 32'h8220000;
      42075: inst = 32'hc20ce94;
      42076: inst = 32'h10408000;
      42077: inst = 32'hc40410d;
      42078: inst = 32'h8220000;
      42079: inst = 32'hc20c632;
      42080: inst = 32'h10408000;
      42081: inst = 32'hc404113;
      42082: inst = 32'h8220000;
      42083: inst = 32'hc204ca9;
      42084: inst = 32'h10408000;
      42085: inst = 32'hc404114;
      42086: inst = 32'h8220000;
      42087: inst = 32'hc207e0d;
      42088: inst = 32'h10408000;
      42089: inst = 32'hc404116;
      42090: inst = 32'h8220000;
      42091: inst = 32'hc20d694;
      42092: inst = 32'h10408000;
      42093: inst = 32'hc404117;
      42094: inst = 32'h8220000;
      42095: inst = 32'h10408000;
      42096: inst = 32'hc4047f3;
      42097: inst = 32'h8220000;
      42098: inst = 32'h10408000;
      42099: inst = 32'hc404919;
      42100: inst = 32'h8220000;
      42101: inst = 32'hc20eed7;
      42102: inst = 32'h10408000;
      42103: inst = 32'hc404151;
      42104: inst = 32'h8220000;
      42105: inst = 32'h10408000;
      42106: inst = 32'hc4041b4;
      42107: inst = 32'h8220000;
      42108: inst = 32'h10408000;
      42109: inst = 32'hc404217;
      42110: inst = 32'h8220000;
      42111: inst = 32'h10408000;
      42112: inst = 32'hc404218;
      42113: inst = 32'h8220000;
      42114: inst = 32'h10408000;
      42115: inst = 32'hc404270;
      42116: inst = 32'h8220000;
      42117: inst = 32'h10408000;
      42118: inst = 32'hc404277;
      42119: inst = 32'h8220000;
      42120: inst = 32'h10408000;
      42121: inst = 32'hc4042d0;
      42122: inst = 32'h8220000;
      42123: inst = 32'h10408000;
      42124: inst = 32'hc4042d4;
      42125: inst = 32'h8220000;
      42126: inst = 32'h10408000;
      42127: inst = 32'hc404391;
      42128: inst = 32'h8220000;
      42129: inst = 32'h10408000;
      42130: inst = 32'hc404450;
      42131: inst = 32'h8220000;
      42132: inst = 32'h10408000;
      42133: inst = 32'hc404451;
      42134: inst = 32'h8220000;
      42135: inst = 32'h10408000;
      42136: inst = 32'hc404454;
      42137: inst = 32'h8220000;
      42138: inst = 32'h10408000;
      42139: inst = 32'hc40445b;
      42140: inst = 32'h8220000;
      42141: inst = 32'h10408000;
      42142: inst = 32'hc40451c;
      42143: inst = 32'h8220000;
      42144: inst = 32'h10408000;
      42145: inst = 32'hc4053c8;
      42146: inst = 32'h8220000;
      42147: inst = 32'h10408000;
      42148: inst = 32'hc4053ce;
      42149: inst = 32'h8220000;
      42150: inst = 32'hc20f73a;
      42151: inst = 32'h10408000;
      42152: inst = 32'hc404152;
      42153: inst = 32'h8220000;
      42154: inst = 32'h10408000;
      42155: inst = 32'hc40415b;
      42156: inst = 32'h8220000;
      42157: inst = 32'h10408000;
      42158: inst = 32'hc40415c;
      42159: inst = 32'h8220000;
      42160: inst = 32'h10408000;
      42161: inst = 32'hc40421a;
      42162: inst = 32'h8220000;
      42163: inst = 32'h10408000;
      42164: inst = 32'hc4042d7;
      42165: inst = 32'h8220000;
      42166: inst = 32'h10408000;
      42167: inst = 32'hc4042d8;
      42168: inst = 32'h8220000;
      42169: inst = 32'h10408000;
      42170: inst = 32'hc4042d9;
      42171: inst = 32'h8220000;
      42172: inst = 32'h10408000;
      42173: inst = 32'hc40433b;
      42174: inst = 32'h8220000;
      42175: inst = 32'h10408000;
      42176: inst = 32'hc40439c;
      42177: inst = 32'h8220000;
      42178: inst = 32'h10408000;
      42179: inst = 32'hc4044b3;
      42180: inst = 32'h8220000;
      42181: inst = 32'h10408000;
      42182: inst = 32'hc4044b5;
      42183: inst = 32'h8220000;
      42184: inst = 32'h10408000;
      42185: inst = 32'hc404577;
      42186: inst = 32'h8220000;
      42187: inst = 32'h10408000;
      42188: inst = 32'hc4045d8;
      42189: inst = 32'h8220000;
      42190: inst = 32'h10408000;
      42191: inst = 32'hc4045d9;
      42192: inst = 32'h8220000;
      42193: inst = 32'hc20f75b;
      42194: inst = 32'h10408000;
      42195: inst = 32'hc404153;
      42196: inst = 32'h8220000;
      42197: inst = 32'h10408000;
      42198: inst = 32'hc404157;
      42199: inst = 32'h8220000;
      42200: inst = 32'h10408000;
      42201: inst = 32'hc4041b2;
      42202: inst = 32'h8220000;
      42203: inst = 32'h10408000;
      42204: inst = 32'hc404271;
      42205: inst = 32'h8220000;
      42206: inst = 32'h10408000;
      42207: inst = 32'hc404276;
      42208: inst = 32'h8220000;
      42209: inst = 32'h10408000;
      42210: inst = 32'hc4042dc;
      42211: inst = 32'h8220000;
      42212: inst = 32'h10408000;
      42213: inst = 32'hc404336;
      42214: inst = 32'h8220000;
      42215: inst = 32'h10408000;
      42216: inst = 32'hc404394;
      42217: inst = 32'h8220000;
      42218: inst = 32'h10408000;
      42219: inst = 32'hc4043f0;
      42220: inst = 32'h8220000;
      42221: inst = 32'h10408000;
      42222: inst = 32'hc4043fb;
      42223: inst = 32'h8220000;
      42224: inst = 32'h10408000;
      42225: inst = 32'hc404510;
      42226: inst = 32'h8220000;
      42227: inst = 32'h10408000;
      42228: inst = 32'hc404516;
      42229: inst = 32'h8220000;
      42230: inst = 32'h10408000;
      42231: inst = 32'hc404574;
      42232: inst = 32'h8220000;
      42233: inst = 32'hc20f739;
      42234: inst = 32'h10408000;
      42235: inst = 32'hc404156;
      42236: inst = 32'h8220000;
      42237: inst = 32'h10408000;
      42238: inst = 32'hc4041b6;
      42239: inst = 32'h8220000;
      42240: inst = 32'h10408000;
      42241: inst = 32'hc404213;
      42242: inst = 32'h8220000;
      42243: inst = 32'h10408000;
      42244: inst = 32'hc404399;
      42245: inst = 32'h8220000;
      42246: inst = 32'h10408000;
      42247: inst = 32'hc404517;
      42248: inst = 32'h8220000;
      42249: inst = 32'h10408000;
      42250: inst = 32'hc404576;
      42251: inst = 32'h8220000;
      42252: inst = 32'h10408000;
      42253: inst = 32'hc4045d1;
      42254: inst = 32'h8220000;
      42255: inst = 32'h10408000;
      42256: inst = 32'hc4045dc;
      42257: inst = 32'h8220000;
      42258: inst = 32'hc20ffde;
      42259: inst = 32'h10408000;
      42260: inst = 32'hc404158;
      42261: inst = 32'h8220000;
      42262: inst = 32'h10408000;
      42263: inst = 32'hc4041b9;
      42264: inst = 32'h8220000;
      42265: inst = 32'h10408000;
      42266: inst = 32'hc404392;
      42267: inst = 32'h8220000;
      42268: inst = 32'h10408000;
      42269: inst = 32'hc4043f2;
      42270: inst = 32'h8220000;
      42271: inst = 32'h10408000;
      42272: inst = 32'hc4043f7;
      42273: inst = 32'h8220000;
      42274: inst = 32'h10408000;
      42275: inst = 32'hc4044b9;
      42276: inst = 32'h8220000;
      42277: inst = 32'hc20f75a;
      42278: inst = 32'h10408000;
      42279: inst = 32'hc404159;
      42280: inst = 32'h8220000;
      42281: inst = 32'h10408000;
      42282: inst = 32'hc40415a;
      42283: inst = 32'h8220000;
      42284: inst = 32'h10408000;
      42285: inst = 32'hc404272;
      42286: inst = 32'h8220000;
      42287: inst = 32'h10408000;
      42288: inst = 32'hc404273;
      42289: inst = 32'h8220000;
      42290: inst = 32'h10408000;
      42291: inst = 32'hc404331;
      42292: inst = 32'h8220000;
      42293: inst = 32'h10408000;
      42294: inst = 32'hc4043f3;
      42295: inst = 32'h8220000;
      42296: inst = 32'h10408000;
      42297: inst = 32'hc4043fc;
      42298: inst = 32'h8220000;
      42299: inst = 32'h10408000;
      42300: inst = 32'hc404452;
      42301: inst = 32'h8220000;
      42302: inst = 32'h10408000;
      42303: inst = 32'hc404456;
      42304: inst = 32'h8220000;
      42305: inst = 32'h10408000;
      42306: inst = 32'hc404459;
      42307: inst = 32'h8220000;
      42308: inst = 32'h10408000;
      42309: inst = 32'hc40445a;
      42310: inst = 32'h8220000;
      42311: inst = 32'h10408000;
      42312: inst = 32'hc4044bb;
      42313: inst = 32'h8220000;
      42314: inst = 32'h10408000;
      42315: inst = 32'hc40451a;
      42316: inst = 32'h8220000;
      42317: inst = 32'h10408000;
      42318: inst = 32'hc404570;
      42319: inst = 32'h8220000;
      42320: inst = 32'h10408000;
      42321: inst = 32'hc404573;
      42322: inst = 32'h8220000;
      42323: inst = 32'hc20dbe7;
      42324: inst = 32'h10408000;
      42325: inst = 32'hc404165;
      42326: inst = 32'h8220000;
      42327: inst = 32'hc20f77c;
      42328: inst = 32'h10408000;
      42329: inst = 32'hc404166;
      42330: inst = 32'h8220000;
      42331: inst = 32'h10408000;
      42332: inst = 32'hc4041b8;
      42333: inst = 32'h8220000;
      42334: inst = 32'hc20e3a4;
      42335: inst = 32'h10408000;
      42336: inst = 32'hc40416a;
      42337: inst = 32'h8220000;
      42338: inst = 32'h10408000;
      42339: inst = 32'hc405415;
      42340: inst = 32'h8220000;
      42341: inst = 32'h10408000;
      42342: inst = 32'hc405534;
      42343: inst = 32'h8220000;
      42344: inst = 32'h10408000;
      42345: inst = 32'hc405655;
      42346: inst = 32'h8220000;
      42347: inst = 32'hc20e3c5;
      42348: inst = 32'h10408000;
      42349: inst = 32'hc40416b;
      42350: inst = 32'h8220000;
      42351: inst = 32'h10408000;
      42352: inst = 32'hc40428b;
      42353: inst = 32'h8220000;
      42354: inst = 32'h10408000;
      42355: inst = 32'hc4053b5;
      42356: inst = 32'h8220000;
      42357: inst = 32'h10408000;
      42358: inst = 32'hc405595;
      42359: inst = 32'h8220000;
      42360: inst = 32'h10408000;
      42361: inst = 32'hc4055f5;
      42362: inst = 32'h8220000;
      42363: inst = 32'hc206e0c;
      42364: inst = 32'h10408000;
      42365: inst = 32'hc40416d;
      42366: inst = 32'h8220000;
      42367: inst = 32'hc209e50;
      42368: inst = 32'h10408000;
      42369: inst = 32'hc404176;
      42370: inst = 32'h8220000;
      42371: inst = 32'hc20860e;
      42372: inst = 32'h10408000;
      42373: inst = 32'hc404177;
      42374: inst = 32'h8220000;
      42375: inst = 32'hc20b5f1;
      42376: inst = 32'h10408000;
      42377: inst = 32'hc40417b;
      42378: inst = 32'h8220000;
      42379: inst = 32'hc20ffbd;
      42380: inst = 32'h10408000;
      42381: inst = 32'hc4041b1;
      42382: inst = 32'h8220000;
      42383: inst = 32'h10408000;
      42384: inst = 32'hc404279;
      42385: inst = 32'h8220000;
      42386: inst = 32'h10408000;
      42387: inst = 32'hc404332;
      42388: inst = 32'h8220000;
      42389: inst = 32'h10408000;
      42390: inst = 32'hc404396;
      42391: inst = 32'h8220000;
      42392: inst = 32'h10408000;
      42393: inst = 32'hc404457;
      42394: inst = 32'h8220000;
      42395: inst = 32'h10408000;
      42396: inst = 32'hc40445c;
      42397: inst = 32'h8220000;
      42398: inst = 32'h10408000;
      42399: inst = 32'hc4044bc;
      42400: inst = 32'h8220000;
      42401: inst = 32'hc20f6f8;
      42402: inst = 32'h10408000;
      42403: inst = 32'hc4041b3;
      42404: inst = 32'h8220000;
      42405: inst = 32'h10408000;
      42406: inst = 32'hc404215;
      42407: inst = 32'h8220000;
      42408: inst = 32'h10408000;
      42409: inst = 32'hc40421b;
      42410: inst = 32'h8220000;
      42411: inst = 32'h10408000;
      42412: inst = 32'hc4043f5;
      42413: inst = 32'h8220000;
      42414: inst = 32'h10408000;
      42415: inst = 32'hc4043f8;
      42416: inst = 32'h8220000;
      42417: inst = 32'h10408000;
      42418: inst = 32'hc404572;
      42419: inst = 32'h8220000;
      42420: inst = 32'hc20f719;
      42421: inst = 32'h10408000;
      42422: inst = 32'hc4041ba;
      42423: inst = 32'h8220000;
      42424: inst = 32'h10408000;
      42425: inst = 32'hc4041bb;
      42426: inst = 32'h8220000;
      42427: inst = 32'h10408000;
      42428: inst = 32'hc404335;
      42429: inst = 32'h8220000;
      42430: inst = 32'h10408000;
      42431: inst = 32'hc404337;
      42432: inst = 32'h8220000;
      42433: inst = 32'h10408000;
      42434: inst = 32'hc40433a;
      42435: inst = 32'h8220000;
      42436: inst = 32'h10408000;
      42437: inst = 32'hc404393;
      42438: inst = 32'h8220000;
      42439: inst = 32'h10408000;
      42440: inst = 32'hc4043f4;
      42441: inst = 32'h8220000;
      42442: inst = 32'h10408000;
      42443: inst = 32'hc4044b8;
      42444: inst = 32'h8220000;
      42445: inst = 32'h10408000;
      42446: inst = 32'hc404511;
      42447: inst = 32'h8220000;
      42448: inst = 32'h10408000;
      42449: inst = 32'hc404518;
      42450: inst = 32'h8220000;
      42451: inst = 32'h10408000;
      42452: inst = 32'hc40451b;
      42453: inst = 32'h8220000;
      42454: inst = 32'h10408000;
      42455: inst = 32'hc404575;
      42456: inst = 32'h8220000;
      42457: inst = 32'hc20ffbe;
      42458: inst = 32'h10408000;
      42459: inst = 32'hc4041bc;
      42460: inst = 32'h8220000;
      42461: inst = 32'h10408000;
      42462: inst = 32'hc404275;
      42463: inst = 32'h8220000;
      42464: inst = 32'hc20db85;
      42465: inst = 32'h10408000;
      42466: inst = 32'hc4041c5;
      42467: inst = 32'h8220000;
      42468: inst = 32'h10408000;
      42469: inst = 32'hc404225;
      42470: inst = 32'h8220000;
      42471: inst = 32'h10408000;
      42472: inst = 32'hc404285;
      42473: inst = 32'h8220000;
      42474: inst = 32'h10408000;
      42475: inst = 32'hc4042e5;
      42476: inst = 32'h8220000;
      42477: inst = 32'hc20c44c;
      42478: inst = 32'h10408000;
      42479: inst = 32'hc4041ca;
      42480: inst = 32'h8220000;
      42481: inst = 32'hc20cbe8;
      42482: inst = 32'h10408000;
      42483: inst = 32'hc4041cb;
      42484: inst = 32'h8220000;
      42485: inst = 32'hc20cba5;
      42486: inst = 32'h10408000;
      42487: inst = 32'hc4041cc;
      42488: inst = 32'h8220000;
      42489: inst = 32'h10408000;
      42490: inst = 32'hc40422c;
      42491: inst = 32'h8220000;
      42492: inst = 32'hc20c633;
      42493: inst = 32'h10408000;
      42494: inst = 32'hc4041d0;
      42495: inst = 32'h8220000;
      42496: inst = 32'hc205cca;
      42497: inst = 32'h10408000;
      42498: inst = 32'hc4041d1;
      42499: inst = 32'h8220000;
      42500: inst = 32'hc20e6b6;
      42501: inst = 32'h10408000;
      42502: inst = 32'hc4041d6;
      42503: inst = 32'h8220000;
      42504: inst = 32'h10408000;
      42505: inst = 32'hc40478f;
      42506: inst = 32'h8220000;
      42507: inst = 32'h10408000;
      42508: inst = 32'hc4047eb;
      42509: inst = 32'h8220000;
      42510: inst = 32'h10408000;
      42511: inst = 32'hc4047f2;
      42512: inst = 32'h8220000;
      42513: inst = 32'h10408000;
      42514: inst = 32'hc4048b6;
      42515: inst = 32'h8220000;
      42516: inst = 32'hc2055ca;
      42517: inst = 32'h10408000;
      42518: inst = 32'hc4041d7;
      42519: inst = 32'h8220000;
      42520: inst = 32'hc20de95;
      42521: inst = 32'h10408000;
      42522: inst = 32'hc4041d8;
      42523: inst = 32'h8220000;
      42524: inst = 32'h10408000;
      42525: inst = 32'hc40429b;
      42526: inst = 32'h8220000;
      42527: inst = 32'h10408000;
      42528: inst = 32'hc404792;
      42529: inst = 32'h8220000;
      42530: inst = 32'h10408000;
      42531: inst = 32'hc404798;
      42532: inst = 32'h8220000;
      42533: inst = 32'h10408000;
      42534: inst = 32'hc4047f5;
      42535: inst = 32'h8220000;
      42536: inst = 32'h10408000;
      42537: inst = 32'hc404857;
      42538: inst = 32'h8220000;
      42539: inst = 32'h10408000;
      42540: inst = 32'hc404915;
      42541: inst = 32'h8220000;
      42542: inst = 32'hc2054c9;
      42543: inst = 32'h10408000;
      42544: inst = 32'hc4041db;
      42545: inst = 32'h8220000;
      42546: inst = 32'h10408000;
      42547: inst = 32'hc404230;
      42548: inst = 32'h8220000;
      42549: inst = 32'hc20de75;
      42550: inst = 32'h10408000;
      42551: inst = 32'hc4041dc;
      42552: inst = 32'h8220000;
      42553: inst = 32'hc20f718;
      42554: inst = 32'h10408000;
      42555: inst = 32'hc404210;
      42556: inst = 32'h8220000;
      42557: inst = 32'h10408000;
      42558: inst = 32'hc404278;
      42559: inst = 32'h8220000;
      42560: inst = 32'hc20ff9d;
      42561: inst = 32'h10408000;
      42562: inst = 32'hc404211;
      42563: inst = 32'h8220000;
      42564: inst = 32'h10408000;
      42565: inst = 32'hc404219;
      42566: inst = 32'h8220000;
      42567: inst = 32'h10408000;
      42568: inst = 32'hc4042d6;
      42569: inst = 32'h8220000;
      42570: inst = 32'hc20ff9c;
      42571: inst = 32'h10408000;
      42572: inst = 32'hc404212;
      42573: inst = 32'h8220000;
      42574: inst = 32'h10408000;
      42575: inst = 32'hc404216;
      42576: inst = 32'h8220000;
      42577: inst = 32'h10408000;
      42578: inst = 32'hc40421c;
      42579: inst = 32'h8220000;
      42580: inst = 32'h10408000;
      42581: inst = 32'hc40427b;
      42582: inst = 32'h8220000;
      42583: inst = 32'h10408000;
      42584: inst = 32'hc4042d1;
      42585: inst = 32'h8220000;
      42586: inst = 32'h10408000;
      42587: inst = 32'hc4042d5;
      42588: inst = 32'h8220000;
      42589: inst = 32'h10408000;
      42590: inst = 32'hc40433c;
      42591: inst = 32'h8220000;
      42592: inst = 32'h10408000;
      42593: inst = 32'hc404395;
      42594: inst = 32'h8220000;
      42595: inst = 32'h10408000;
      42596: inst = 32'hc404397;
      42597: inst = 32'h8220000;
      42598: inst = 32'h10408000;
      42599: inst = 32'hc404398;
      42600: inst = 32'h8220000;
      42601: inst = 32'h10408000;
      42602: inst = 32'hc40439a;
      42603: inst = 32'h8220000;
      42604: inst = 32'h10408000;
      42605: inst = 32'hc4043f1;
      42606: inst = 32'h8220000;
      42607: inst = 32'h10408000;
      42608: inst = 32'hc404514;
      42609: inst = 32'h8220000;
      42610: inst = 32'h10408000;
      42611: inst = 32'hc4045d2;
      42612: inst = 32'h8220000;
      42613: inst = 32'hc20a46f;
      42614: inst = 32'h10408000;
      42615: inst = 32'hc40422a;
      42616: inst = 32'h8220000;
      42617: inst = 32'hc20d3c7;
      42618: inst = 32'h10408000;
      42619: inst = 32'hc40422b;
      42620: inst = 32'h8220000;
      42621: inst = 32'h10408000;
      42622: inst = 32'hc405475;
      42623: inst = 32'h8220000;
      42624: inst = 32'hc20ce53;
      42625: inst = 32'h10408000;
      42626: inst = 32'hc40422f;
      42627: inst = 32'h8220000;
      42628: inst = 32'hc207d4d;
      42629: inst = 32'h10408000;
      42630: inst = 32'hc40423b;
      42631: inst = 32'h8220000;
      42632: inst = 32'h10408000;
      42633: inst = 32'hc40423c;
      42634: inst = 32'h8220000;
      42635: inst = 32'hc20ff7c;
      42636: inst = 32'h10408000;
      42637: inst = 32'hc40427c;
      42638: inst = 32'h8220000;
      42639: inst = 32'h10408000;
      42640: inst = 32'hc4042d2;
      42641: inst = 32'h8220000;
      42642: inst = 32'h10408000;
      42643: inst = 32'hc404338;
      42644: inst = 32'h8220000;
      42645: inst = 32'h10408000;
      42646: inst = 32'hc4043f6;
      42647: inst = 32'h8220000;
      42648: inst = 32'h10408000;
      42649: inst = 32'hc4044b4;
      42650: inst = 32'h8220000;
      42651: inst = 32'h10408000;
      42652: inst = 32'hc404571;
      42653: inst = 32'h8220000;
      42654: inst = 32'h10408000;
      42655: inst = 32'hc404578;
      42656: inst = 32'h8220000;
      42657: inst = 32'h10408000;
      42658: inst = 32'hc404579;
      42659: inst = 32'h8220000;
      42660: inst = 32'hc20be12;
      42661: inst = 32'h10408000;
      42662: inst = 32'hc40428f;
      42663: inst = 32'h8220000;
      42664: inst = 32'hc209db0;
      42665: inst = 32'h10408000;
      42666: inst = 32'hc40429c;
      42667: inst = 32'h8220000;
      42668: inst = 32'hc20cb65;
      42669: inst = 32'h10408000;
      42670: inst = 32'hc4043a4;
      42671: inst = 32'h8220000;
      42672: inst = 32'h10408000;
      42673: inst = 32'hc4043ac;
      42674: inst = 32'h8220000;
      42675: inst = 32'hc20cb43;
      42676: inst = 32'h10408000;
      42677: inst = 32'hc4043a5;
      42678: inst = 32'h8220000;
      42679: inst = 32'h10408000;
      42680: inst = 32'hc405355;
      42681: inst = 32'h8220000;
      42682: inst = 32'h10408000;
      42683: inst = 32'hc405712;
      42684: inst = 32'h8220000;
      42685: inst = 32'hc205bce;
      42686: inst = 32'h10408000;
      42687: inst = 32'hc40466b;
      42688: inst = 32'h8220000;
      42689: inst = 32'h10408000;
      42690: inst = 32'hc404670;
      42691: inst = 32'h8220000;
      42692: inst = 32'h10408000;
      42693: inst = 32'hc404674;
      42694: inst = 32'h8220000;
      42695: inst = 32'h10408000;
      42696: inst = 32'hc4046d2;
      42697: inst = 32'h8220000;
      42698: inst = 32'h10408000;
      42699: inst = 32'hc404735;
      42700: inst = 32'h8220000;
      42701: inst = 32'h10408000;
      42702: inst = 32'hc404739;
      42703: inst = 32'h8220000;
      42704: inst = 32'hc205c2c;
      42705: inst = 32'h10408000;
      42706: inst = 32'hc40466c;
      42707: inst = 32'h8220000;
      42708: inst = 32'hc2063ce;
      42709: inst = 32'h10408000;
      42710: inst = 32'hc404671;
      42711: inst = 32'h8220000;
      42712: inst = 32'hc205bed;
      42713: inst = 32'h10408000;
      42714: inst = 32'hc404672;
      42715: inst = 32'h8220000;
      42716: inst = 32'h10408000;
      42717: inst = 32'hc404678;
      42718: inst = 32'h8220000;
      42719: inst = 32'h10408000;
      42720: inst = 32'hc4046d3;
      42721: inst = 32'h8220000;
      42722: inst = 32'h10408000;
      42723: inst = 32'hc4046d8;
      42724: inst = 32'h8220000;
      42725: inst = 32'h10408000;
      42726: inst = 32'hc404733;
      42727: inst = 32'h8220000;
      42728: inst = 32'hc204c8a;
      42729: inst = 32'h10408000;
      42730: inst = 32'hc4046cb;
      42731: inst = 32'h8220000;
      42732: inst = 32'h10408000;
      42733: inst = 32'hc404734;
      42734: inst = 32'h8220000;
      42735: inst = 32'hc20542c;
      42736: inst = 32'h10408000;
      42737: inst = 32'hc4046d4;
      42738: inst = 32'h8220000;
      42739: inst = 32'h10408000;
      42740: inst = 32'hc40472c;
      42741: inst = 32'h8220000;
      42742: inst = 32'hc205c0d;
      42743: inst = 32'h10408000;
      42744: inst = 32'hc4046d9;
      42745: inst = 32'h8220000;
      42746: inst = 32'h10408000;
      42747: inst = 32'hc404731;
      42748: inst = 32'h8220000;
      42749: inst = 32'hc20e6b5;
      42750: inst = 32'h10408000;
      42751: inst = 32'hc40478b;
      42752: inst = 32'h8220000;
      42753: inst = 32'h10408000;
      42754: inst = 32'hc4048b9;
      42755: inst = 32'h8220000;
      42756: inst = 32'hc20ae51;
      42757: inst = 32'h10408000;
      42758: inst = 32'hc40478c;
      42759: inst = 32'h8220000;
      42760: inst = 32'hc20960e;
      42761: inst = 32'h10408000;
      42762: inst = 32'hc40478d;
      42763: inst = 32'h8220000;
      42764: inst = 32'hc20c673;
      42765: inst = 32'h10408000;
      42766: inst = 32'hc40478e;
      42767: inst = 32'h8220000;
      42768: inst = 32'h10408000;
      42769: inst = 32'hc404793;
      42770: inst = 32'h8220000;
      42771: inst = 32'h10408000;
      42772: inst = 32'hc404854;
      42773: inst = 32'h8220000;
      42774: inst = 32'hc20be52;
      42775: inst = 32'h10408000;
      42776: inst = 32'hc404790;
      42777: inst = 32'h8220000;
      42778: inst = 32'h10408000;
      42779: inst = 32'hc404858;
      42780: inst = 32'h8220000;
      42781: inst = 32'h10408000;
      42782: inst = 32'hc404859;
      42783: inst = 32'h8220000;
      42784: inst = 32'hc209e2f;
      42785: inst = 32'h10408000;
      42786: inst = 32'hc404791;
      42787: inst = 32'h8220000;
      42788: inst = 32'h10408000;
      42789: inst = 32'hc404794;
      42790: inst = 32'h8220000;
      42791: inst = 32'hc20ae30;
      42792: inst = 32'h10408000;
      42793: inst = 32'hc4047ec;
      42794: inst = 32'h8220000;
      42795: inst = 32'h10408000;
      42796: inst = 32'hc4047f1;
      42797: inst = 32'h8220000;
      42798: inst = 32'hc20ce73;
      42799: inst = 32'h10408000;
      42800: inst = 32'hc4047ed;
      42801: inst = 32'h8220000;
      42802: inst = 32'h10408000;
      42803: inst = 32'hc4048b4;
      42804: inst = 32'h8220000;
      42805: inst = 32'hc208e0e;
      42806: inst = 32'h10408000;
      42807: inst = 32'hc4047f0;
      42808: inst = 32'h8220000;
      42809: inst = 32'h10408000;
      42810: inst = 32'hc404855;
      42811: inst = 32'h8220000;
      42812: inst = 32'hc2085ed;
      42813: inst = 32'h10408000;
      42814: inst = 32'hc4047f4;
      42815: inst = 32'h8220000;
      42816: inst = 32'h10408000;
      42817: inst = 32'hc4048b8;
      42818: inst = 32'h8220000;
      42819: inst = 32'hc20b651;
      42820: inst = 32'h10408000;
      42821: inst = 32'hc4047f8;
      42822: inst = 32'h8220000;
      42823: inst = 32'h10408000;
      42824: inst = 32'hc404914;
      42825: inst = 32'h8220000;
      42826: inst = 32'hc20c672;
      42827: inst = 32'h10408000;
      42828: inst = 32'hc4047f9;
      42829: inst = 32'h8220000;
      42830: inst = 32'h10408000;
      42831: inst = 32'hc404856;
      42832: inst = 32'h8220000;
      42833: inst = 32'h10408000;
      42834: inst = 32'hc4048b7;
      42835: inst = 32'h8220000;
      42836: inst = 32'hc209e0f;
      42837: inst = 32'h10408000;
      42838: inst = 32'hc4048b5;
      42839: inst = 32'h8220000;
      42840: inst = 32'h10408000;
      42841: inst = 32'hc404918;
      42842: inst = 32'h8220000;
      42843: inst = 32'hc20de94;
      42844: inst = 32'h10408000;
      42845: inst = 32'hc404917;
      42846: inst = 32'h8220000;
      42847: inst = 32'hc20c2e2;
      42848: inst = 32'h10408000;
      42849: inst = 32'hc405352;
      42850: inst = 32'h8220000;
      42851: inst = 32'hc20cb23;
      42852: inst = 32'h10408000;
      42853: inst = 32'hc405353;
      42854: inst = 32'h8220000;
      42855: inst = 32'h10408000;
      42856: inst = 32'hc405356;
      42857: inst = 32'h8220000;
      42858: inst = 32'h10408000;
      42859: inst = 32'hc405357;
      42860: inst = 32'h8220000;
      42861: inst = 32'h10408000;
      42862: inst = 32'hc405358;
      42863: inst = 32'h8220000;
      42864: inst = 32'h10408000;
      42865: inst = 32'hc405359;
      42866: inst = 32'h8220000;
      42867: inst = 32'h10408000;
      42868: inst = 32'hc40535a;
      42869: inst = 32'h8220000;
      42870: inst = 32'h10408000;
      42871: inst = 32'hc405592;
      42872: inst = 32'h8220000;
      42873: inst = 32'h10408000;
      42874: inst = 32'hc4055f2;
      42875: inst = 32'h8220000;
      42876: inst = 32'h10408000;
      42877: inst = 32'hc405652;
      42878: inst = 32'h8220000;
      42879: inst = 32'h10408000;
      42880: inst = 32'hc4056b2;
      42881: inst = 32'h8220000;
      42882: inst = 32'hc20c323;
      42883: inst = 32'h10408000;
      42884: inst = 32'hc40535b;
      42885: inst = 32'h8220000;
      42886: inst = 32'h10408000;
      42887: inst = 32'hc4057d2;
      42888: inst = 32'h8220000;
      42889: inst = 32'hc20e407;
      42890: inst = 32'h10408000;
      42891: inst = 32'hc4053b3;
      42892: inst = 32'h8220000;
      42893: inst = 32'hc207d9a;
      42894: inst = 32'h10408000;
      42895: inst = 32'hc4053b6;
      42896: inst = 32'h8220000;
      42897: inst = 32'hc2065fe;
      42898: inst = 32'h10408000;
      42899: inst = 32'hc4053b7;
      42900: inst = 32'h8220000;
      42901: inst = 32'hc2065fd;
      42902: inst = 32'h10408000;
      42903: inst = 32'hc4053b8;
      42904: inst = 32'h8220000;
      42905: inst = 32'h10408000;
      42906: inst = 32'hc4053b9;
      42907: inst = 32'h8220000;
      42908: inst = 32'hc20661e;
      42909: inst = 32'h10408000;
      42910: inst = 32'hc4053ba;
      42911: inst = 32'h8220000;
      42912: inst = 32'hc20bb86;
      42913: inst = 32'h10408000;
      42914: inst = 32'hc4053bb;
      42915: inst = 32'h8220000;
      42916: inst = 32'h10408000;
      42917: inst = 32'hc4054db;
      42918: inst = 32'h8220000;
      42919: inst = 32'hc20e6fa;
      42920: inst = 32'h10408000;
      42921: inst = 32'hc4053c9;
      42922: inst = 32'h8220000;
      42923: inst = 32'h10408000;
      42924: inst = 32'hc4053cd;
      42925: inst = 32'h8220000;
      42926: inst = 32'h10408000;
      42927: inst = 32'hc4055a7;
      42928: inst = 32'h8220000;
      42929: inst = 32'hc20e6fb;
      42930: inst = 32'h10408000;
      42931: inst = 32'hc4053ca;
      42932: inst = 32'h8220000;
      42933: inst = 32'h10408000;
      42934: inst = 32'hc4053cc;
      42935: inst = 32'h8220000;
      42936: inst = 32'h10408000;
      42937: inst = 32'hc405487;
      42938: inst = 32'h8220000;
      42939: inst = 32'h10408000;
      42940: inst = 32'hc40548f;
      42941: inst = 32'h8220000;
      42942: inst = 32'h10408000;
      42943: inst = 32'hc405547;
      42944: inst = 32'h8220000;
      42945: inst = 32'h10408000;
      42946: inst = 32'hc40554f;
      42947: inst = 32'h8220000;
      42948: inst = 32'hc20defb;
      42949: inst = 32'h10408000;
      42950: inst = 32'hc4053cb;
      42951: inst = 32'h8220000;
      42952: inst = 32'h10408000;
      42953: inst = 32'hc405428;
      42954: inst = 32'h8220000;
      42955: inst = 32'h10408000;
      42956: inst = 32'hc405429;
      42957: inst = 32'h8220000;
      42958: inst = 32'h10408000;
      42959: inst = 32'hc40542a;
      42960: inst = 32'h8220000;
      42961: inst = 32'h10408000;
      42962: inst = 32'hc40542b;
      42963: inst = 32'h8220000;
      42964: inst = 32'h10408000;
      42965: inst = 32'hc40542c;
      42966: inst = 32'h8220000;
      42967: inst = 32'h10408000;
      42968: inst = 32'hc40542d;
      42969: inst = 32'h8220000;
      42970: inst = 32'h10408000;
      42971: inst = 32'hc40542e;
      42972: inst = 32'h8220000;
      42973: inst = 32'h10408000;
      42974: inst = 32'hc405488;
      42975: inst = 32'h8220000;
      42976: inst = 32'h10408000;
      42977: inst = 32'hc405489;
      42978: inst = 32'h8220000;
      42979: inst = 32'h10408000;
      42980: inst = 32'hc40548a;
      42981: inst = 32'h8220000;
      42982: inst = 32'h10408000;
      42983: inst = 32'hc40548b;
      42984: inst = 32'h8220000;
      42985: inst = 32'h10408000;
      42986: inst = 32'hc40548c;
      42987: inst = 32'h8220000;
      42988: inst = 32'h10408000;
      42989: inst = 32'hc40548d;
      42990: inst = 32'h8220000;
      42991: inst = 32'h10408000;
      42992: inst = 32'hc40548e;
      42993: inst = 32'h8220000;
      42994: inst = 32'h10408000;
      42995: inst = 32'hc4054e7;
      42996: inst = 32'h8220000;
      42997: inst = 32'h10408000;
      42998: inst = 32'hc4054ea;
      42999: inst = 32'h8220000;
      43000: inst = 32'h10408000;
      43001: inst = 32'hc4054ed;
      43002: inst = 32'h8220000;
      43003: inst = 32'h10408000;
      43004: inst = 32'hc4054ee;
      43005: inst = 32'h8220000;
      43006: inst = 32'h10408000;
      43007: inst = 32'hc4054ef;
      43008: inst = 32'h8220000;
      43009: inst = 32'h10408000;
      43010: inst = 32'hc40554a;
      43011: inst = 32'h8220000;
      43012: inst = 32'h10408000;
      43013: inst = 32'hc40554d;
      43014: inst = 32'h8220000;
      43015: inst = 32'h10408000;
      43016: inst = 32'hc40554e;
      43017: inst = 32'h8220000;
      43018: inst = 32'h10408000;
      43019: inst = 32'hc4055a8;
      43020: inst = 32'h8220000;
      43021: inst = 32'h10408000;
      43022: inst = 32'hc4055a9;
      43023: inst = 32'h8220000;
      43024: inst = 32'h10408000;
      43025: inst = 32'hc4055aa;
      43026: inst = 32'h8220000;
      43027: inst = 32'h10408000;
      43028: inst = 32'hc4055ab;
      43029: inst = 32'h8220000;
      43030: inst = 32'h10408000;
      43031: inst = 32'hc4055ac;
      43032: inst = 32'h8220000;
      43033: inst = 32'h10408000;
      43034: inst = 32'hc4055ad;
      43035: inst = 32'h8220000;
      43036: inst = 32'h10408000;
      43037: inst = 32'hc4055ae;
      43038: inst = 32'h8220000;
      43039: inst = 32'h10408000;
      43040: inst = 32'hc405609;
      43041: inst = 32'h8220000;
      43042: inst = 32'h10408000;
      43043: inst = 32'hc40560b;
      43044: inst = 32'h8220000;
      43045: inst = 32'h10408000;
      43046: inst = 32'hc405669;
      43047: inst = 32'h8220000;
      43048: inst = 32'hc20cbc7;
      43049: inst = 32'h10408000;
      43050: inst = 32'hc405412;
      43051: inst = 32'h8220000;
      43052: inst = 32'h10408000;
      43053: inst = 32'hc405472;
      43054: inst = 32'h8220000;
      43055: inst = 32'hc20edb1;
      43056: inst = 32'h10408000;
      43057: inst = 32'hc405413;
      43058: inst = 32'h8220000;
      43059: inst = 32'hc20db43;
      43060: inst = 32'h10408000;
      43061: inst = 32'hc405414;
      43062: inst = 32'h8220000;
      43063: inst = 32'hc207d78;
      43064: inst = 32'h10408000;
      43065: inst = 32'hc405416;
      43066: inst = 32'h8220000;
      43067: inst = 32'hc206dbc;
      43068: inst = 32'h10408000;
      43069: inst = 32'hc405417;
      43070: inst = 32'h8220000;
      43071: inst = 32'h10408000;
      43072: inst = 32'hc405477;
      43073: inst = 32'h8220000;
      43074: inst = 32'hc206dbb;
      43075: inst = 32'h10408000;
      43076: inst = 32'hc405418;
      43077: inst = 32'h8220000;
      43078: inst = 32'h10408000;
      43079: inst = 32'hc405419;
      43080: inst = 32'h8220000;
      43081: inst = 32'h10408000;
      43082: inst = 32'hc405478;
      43083: inst = 32'h8220000;
      43084: inst = 32'h10408000;
      43085: inst = 32'hc405479;
      43086: inst = 32'h8220000;
      43087: inst = 32'hc206ddc;
      43088: inst = 32'h10408000;
      43089: inst = 32'hc40541a;
      43090: inst = 32'h8220000;
      43091: inst = 32'h10408000;
      43092: inst = 32'hc40547a;
      43093: inst = 32'h8220000;
      43094: inst = 32'hc20bb66;
      43095: inst = 32'h10408000;
      43096: inst = 32'hc40541b;
      43097: inst = 32'h8220000;
      43098: inst = 32'h10408000;
      43099: inst = 32'hc40547b;
      43100: inst = 32'h8220000;
      43101: inst = 32'h10408000;
      43102: inst = 32'hc40559b;
      43103: inst = 32'h8220000;
      43104: inst = 32'hc20eed8;
      43105: inst = 32'h10408000;
      43106: inst = 32'hc405427;
      43107: inst = 32'h8220000;
      43108: inst = 32'h10408000;
      43109: inst = 32'hc40542f;
      43110: inst = 32'h8220000;
      43111: inst = 32'hc20edd2;
      43112: inst = 32'h10408000;
      43113: inst = 32'hc405473;
      43114: inst = 32'h8220000;
      43115: inst = 32'hc20db42;
      43116: inst = 32'h10408000;
      43117: inst = 32'hc405474;
      43118: inst = 32'h8220000;
      43119: inst = 32'hc207d79;
      43120: inst = 32'h10408000;
      43121: inst = 32'hc405476;
      43122: inst = 32'h8220000;
      43123: inst = 32'hc20e590;
      43124: inst = 32'h10408000;
      43125: inst = 32'hc4054d3;
      43126: inst = 32'h8220000;
      43127: inst = 32'hc20e363;
      43128: inst = 32'h10408000;
      43129: inst = 32'hc4054d4;
      43130: inst = 32'h8220000;
      43131: inst = 32'hc20d3a6;
      43132: inst = 32'h10408000;
      43133: inst = 32'hc4054d5;
      43134: inst = 32'h8220000;
      43135: inst = 32'hc207dba;
      43136: inst = 32'h10408000;
      43137: inst = 32'hc4054d6;
      43138: inst = 32'h8220000;
      43139: inst = 32'hc2075fd;
      43140: inst = 32'h10408000;
      43141: inst = 32'hc4054d7;
      43142: inst = 32'h8220000;
      43143: inst = 32'h10408000;
      43144: inst = 32'hc4054d8;
      43145: inst = 32'h8220000;
      43146: inst = 32'h10408000;
      43147: inst = 32'hc4054d9;
      43148: inst = 32'h8220000;
      43149: inst = 32'hc206e1e;
      43150: inst = 32'h10408000;
      43151: inst = 32'hc4054da;
      43152: inst = 32'h8220000;
      43153: inst = 32'hc204a69;
      43154: inst = 32'h10408000;
      43155: inst = 32'hc4054e8;
      43156: inst = 32'h8220000;
      43157: inst = 32'h10408000;
      43158: inst = 32'hc4054e9;
      43159: inst = 32'h8220000;
      43160: inst = 32'h10408000;
      43161: inst = 32'hc4054eb;
      43162: inst = 32'h8220000;
      43163: inst = 32'h10408000;
      43164: inst = 32'hc4054ec;
      43165: inst = 32'h8220000;
      43166: inst = 32'h10408000;
      43167: inst = 32'hc405548;
      43168: inst = 32'h8220000;
      43169: inst = 32'h10408000;
      43170: inst = 32'hc405549;
      43171: inst = 32'h8220000;
      43172: inst = 32'h10408000;
      43173: inst = 32'hc40554b;
      43174: inst = 32'h8220000;
      43175: inst = 32'h10408000;
      43176: inst = 32'hc40554c;
      43177: inst = 32'h8220000;
      43178: inst = 32'h10408000;
      43179: inst = 32'hc405608;
      43180: inst = 32'h8220000;
      43181: inst = 32'h10408000;
      43182: inst = 32'hc40560a;
      43183: inst = 32'h8220000;
      43184: inst = 32'h10408000;
      43185: inst = 32'hc40560c;
      43186: inst = 32'h8220000;
      43187: inst = 32'h10408000;
      43188: inst = 32'hc405668;
      43189: inst = 32'h8220000;
      43190: inst = 32'h10408000;
      43191: inst = 32'hc40566a;
      43192: inst = 32'h8220000;
      43193: inst = 32'hc20eba3;
      43194: inst = 32'h10408000;
      43195: inst = 32'hc405535;
      43196: inst = 32'h8220000;
      43197: inst = 32'hc207411;
      43198: inst = 32'h10408000;
      43199: inst = 32'hc405536;
      43200: inst = 32'h8220000;
      43201: inst = 32'hc205bf2;
      43202: inst = 32'h10408000;
      43203: inst = 32'hc405537;
      43204: inst = 32'h8220000;
      43205: inst = 32'h10408000;
      43206: inst = 32'hc40553a;
      43207: inst = 32'h8220000;
      43208: inst = 32'hc205c12;
      43209: inst = 32'h10408000;
      43210: inst = 32'hc405538;
      43211: inst = 32'h8220000;
      43212: inst = 32'h10408000;
      43213: inst = 32'hc405539;
      43214: inst = 32'h8220000;
      43215: inst = 32'h10408000;
      43216: inst = 32'hc4055f9;
      43217: inst = 32'h8220000;
      43218: inst = 32'hc20bb25;
      43219: inst = 32'h10408000;
      43220: inst = 32'hc40553b;
      43221: inst = 32'h8220000;
      43222: inst = 32'h10408000;
      43223: inst = 32'hc4056bb;
      43224: inst = 32'h8220000;
      43225: inst = 32'h10408000;
      43226: inst = 32'hc40571b;
      43227: inst = 32'h8220000;
      43228: inst = 32'h10408000;
      43229: inst = 32'hc40577b;
      43230: inst = 32'h8220000;
      43231: inst = 32'hc20dba4;
      43232: inst = 32'h10408000;
      43233: inst = 32'hc405593;
      43234: inst = 32'h8220000;
      43235: inst = 32'h10408000;
      43236: inst = 32'hc4056b4;
      43237: inst = 32'h8220000;
      43238: inst = 32'hc206288;
      43239: inst = 32'h10408000;
      43240: inst = 32'hc405596;
      43241: inst = 32'h8220000;
      43242: inst = 32'hc205bb1;
      43243: inst = 32'h10408000;
      43244: inst = 32'hc405597;
      43245: inst = 32'h8220000;
      43246: inst = 32'hc2052ec;
      43247: inst = 32'h10408000;
      43248: inst = 32'hc405598;
      43249: inst = 32'h8220000;
      43250: inst = 32'hc20532d;
      43251: inst = 32'h10408000;
      43252: inst = 32'hc405599;
      43253: inst = 32'h8220000;
      43254: inst = 32'hc205390;
      43255: inst = 32'h10408000;
      43256: inst = 32'hc40559a;
      43257: inst = 32'h8220000;
      43258: inst = 32'hc20e6d9;
      43259: inst = 32'h10408000;
      43260: inst = 32'hc4055af;
      43261: inst = 32'h8220000;
      43262: inst = 32'hc2062ea;
      43263: inst = 32'h10408000;
      43264: inst = 32'hc4055f6;
      43265: inst = 32'h8220000;
      43266: inst = 32'hc2064f8;
      43267: inst = 32'h10408000;
      43268: inst = 32'hc4055f7;
      43269: inst = 32'h8220000;
      43270: inst = 32'hc205bd1;
      43271: inst = 32'h10408000;
      43272: inst = 32'hc4055f8;
      43273: inst = 32'h8220000;
      43274: inst = 32'hc2064d6;
      43275: inst = 32'h10408000;
      43276: inst = 32'hc4055fa;
      43277: inst = 32'h8220000;
      43278: inst = 32'hc20bba7;
      43279: inst = 32'h10408000;
      43280: inst = 32'hc4055fb;
      43281: inst = 32'h8220000;
      43282: inst = 32'hc20eeb7;
      43283: inst = 32'h10408000;
      43284: inst = 32'hc405607;
      43285: inst = 32'h8220000;
      43286: inst = 32'hc20d699;
      43287: inst = 32'h10408000;
      43288: inst = 32'hc40560d;
      43289: inst = 32'h8220000;
      43290: inst = 32'hc20b553;
      43291: inst = 32'h10408000;
      43292: inst = 32'hc40560e;
      43293: inst = 32'h8220000;
      43294: inst = 32'hc2083cd;
      43295: inst = 32'h10408000;
      43296: inst = 32'hc40560f;
      43297: inst = 32'h8220000;
      43298: inst = 32'hc20736c;
      43299: inst = 32'h10408000;
      43300: inst = 32'hc405610;
      43301: inst = 32'h8220000;
      43302: inst = 32'hc20a4d0;
      43303: inst = 32'h10408000;
      43304: inst = 32'hc405611;
      43305: inst = 32'h8220000;
      43306: inst = 32'hc20de55;
      43307: inst = 32'h10408000;
      43308: inst = 32'hc405612;
      43309: inst = 32'h8220000;
      43310: inst = 32'hc2062eb;
      43311: inst = 32'h10408000;
      43312: inst = 32'hc405656;
      43313: inst = 32'h8220000;
      43314: inst = 32'hc206496;
      43315: inst = 32'h10408000;
      43316: inst = 32'hc405657;
      43317: inst = 32'h8220000;
      43318: inst = 32'hc205bb0;
      43319: inst = 32'h10408000;
      43320: inst = 32'hc405658;
      43321: inst = 32'h8220000;
      43322: inst = 32'hc2063f2;
      43323: inst = 32'h10408000;
      43324: inst = 32'hc405659;
      43325: inst = 32'h8220000;
      43326: inst = 32'hc206475;
      43327: inst = 32'h10408000;
      43328: inst = 32'hc40565a;
      43329: inst = 32'h8220000;
      43330: inst = 32'hc20bb87;
      43331: inst = 32'h10408000;
      43332: inst = 32'hc40565b;
      43333: inst = 32'h8220000;
      43334: inst = 32'hc209492;
      43335: inst = 32'h10408000;
      43336: inst = 32'hc40566b;
      43337: inst = 32'h8220000;
      43338: inst = 32'hc204228;
      43339: inst = 32'h10408000;
      43340: inst = 32'hc40566c;
      43341: inst = 32'h8220000;
      43342: inst = 32'h10408000;
      43343: inst = 32'hc405760;
      43344: inst = 32'h8220000;
      43345: inst = 32'hc20632c;
      43346: inst = 32'h10408000;
      43347: inst = 32'hc40566d;
      43348: inst = 32'h8220000;
      43349: inst = 32'hc20a4d1;
      43350: inst = 32'h10408000;
      43351: inst = 32'hc40566e;
      43352: inst = 32'h8220000;
      43353: inst = 32'hc20cdf4;
      43354: inst = 32'h10408000;
      43355: inst = 32'hc40566f;
      43356: inst = 32'h8220000;
      43357: inst = 32'hc20c593;
      43358: inst = 32'h10408000;
      43359: inst = 32'hc405670;
      43360: inst = 32'h8220000;
      43361: inst = 32'hc20944f;
      43362: inst = 32'h10408000;
      43363: inst = 32'hc405671;
      43364: inst = 32'h8220000;
      43365: inst = 32'hc20734c;
      43366: inst = 32'h10408000;
      43367: inst = 32'hc405672;
      43368: inst = 32'h8220000;
      43369: inst = 32'hc20a4b0;
      43370: inst = 32'h10408000;
      43371: inst = 32'hc405673;
      43372: inst = 32'h8220000;
      43373: inst = 32'hc20e3e6;
      43374: inst = 32'h10408000;
      43375: inst = 32'hc4056b3;
      43376: inst = 32'h8220000;
      43377: inst = 32'hc209ac5;
      43378: inst = 32'h10408000;
      43379: inst = 32'hc4056b5;
      43380: inst = 32'h8220000;
      43381: inst = 32'hc206350;
      43382: inst = 32'h10408000;
      43383: inst = 32'hc4056ba;
      43384: inst = 32'h8220000;
      43385: inst = 32'h10408000;
      43386: inst = 32'hc40571a;
      43387: inst = 32'h8220000;
      43388: inst = 32'h10408000;
      43389: inst = 32'hc405776;
      43390: inst = 32'h8220000;
      43391: inst = 32'hc2052ac;
      43392: inst = 32'h10408000;
      43393: inst = 32'hc4056ca;
      43394: inst = 32'h8220000;
      43395: inst = 32'h10408000;
      43396: inst = 32'hc4056d0;
      43397: inst = 32'h8220000;
      43398: inst = 32'h10408000;
      43399: inst = 32'hc4057bf;
      43400: inst = 32'h8220000;
      43401: inst = 32'hc204a6a;
      43402: inst = 32'h10408000;
      43403: inst = 32'hc4056cb;
      43404: inst = 32'h8220000;
      43405: inst = 32'h10408000;
      43406: inst = 32'hc4056cc;
      43407: inst = 32'h8220000;
      43408: inst = 32'h10408000;
      43409: inst = 32'hc4056cd;
      43410: inst = 32'h8220000;
      43411: inst = 32'h10408000;
      43412: inst = 32'hc4056ce;
      43413: inst = 32'h8220000;
      43414: inst = 32'h10408000;
      43415: inst = 32'hc4057c0;
      43416: inst = 32'h8220000;
      43417: inst = 32'hc20528b;
      43418: inst = 32'h10408000;
      43419: inst = 32'hc4056cf;
      43420: inst = 32'h8220000;
      43421: inst = 32'hc205acd;
      43422: inst = 32'h10408000;
      43423: inst = 32'hc4056d1;
      43424: inst = 32'h8220000;
      43425: inst = 32'hc205aed;
      43426: inst = 32'h10408000;
      43427: inst = 32'hc4056d2;
      43428: inst = 32'h8220000;
      43429: inst = 32'h10408000;
      43430: inst = 32'hc40575f;
      43431: inst = 32'h8220000;
      43432: inst = 32'hc20632f;
      43433: inst = 32'h10408000;
      43434: inst = 32'hc4056d3;
      43435: inst = 32'h8220000;
      43436: inst = 32'h10408000;
      43437: inst = 32'hc405715;
      43438: inst = 32'h8220000;
      43439: inst = 32'hc20634f;
      43440: inst = 32'h10408000;
      43441: inst = 32'hc4056fe;
      43442: inst = 32'h8220000;
      43443: inst = 32'hc204208;
      43444: inst = 32'h10408000;
      43445: inst = 32'hc4056ff;
      43446: inst = 32'h8220000;
      43447: inst = 32'h10408000;
      43448: inst = 32'hc405700;
      43449: inst = 32'h8220000;
      43450: inst = 32'hc209ae6;
      43451: inst = 32'h10408000;
      43452: inst = 32'hc405714;
      43453: inst = 32'h8220000;
      43454: inst = 32'hc206370;
      43455: inst = 32'h10408000;
      43456: inst = 32'hc405716;
      43457: inst = 32'h8220000;
      43458: inst = 32'h10408000;
      43459: inst = 32'hc405777;
      43460: inst = 32'h8220000;
      43461: inst = 32'h10408000;
      43462: inst = 32'hc405778;
      43463: inst = 32'h8220000;
      43464: inst = 32'h10408000;
      43465: inst = 32'hc405779;
      43466: inst = 32'h8220000;
      43467: inst = 32'hc20c303;
      43468: inst = 32'h10408000;
      43469: inst = 32'hc405772;
      43470: inst = 32'h8220000;
      43471: inst = 32'hc20aaa2;
      43472: inst = 32'h10408000;
      43473: inst = 32'hc405773;
      43474: inst = 32'h8220000;
      43475: inst = 32'hc2072ea;
      43476: inst = 32'h10408000;
      43477: inst = 32'hc405774;
      43478: inst = 32'h8220000;
      43479: inst = 32'hc205b72;
      43480: inst = 32'h10408000;
      43481: inst = 32'hc405775;
      43482: inst = 32'h8220000;
      43483: inst = 32'hc206371;
      43484: inst = 32'h10408000;
      43485: inst = 32'hc40577a;
      43486: inst = 32'h8220000;
      43487: inst = 32'hc20bae3;
      43488: inst = 32'h10408000;
      43489: inst = 32'hc4057d3;
      43490: inst = 32'h8220000;
      43491: inst = 32'hc20bb04;
      43492: inst = 32'h10408000;
      43493: inst = 32'hc4057d4;
      43494: inst = 32'h8220000;
      43495: inst = 32'hc20b325;
      43496: inst = 32'h10408000;
      43497: inst = 32'hc4057d5;
      43498: inst = 32'h8220000;
      43499: inst = 32'h10408000;
      43500: inst = 32'hc4057d6;
      43501: inst = 32'h8220000;
      43502: inst = 32'h10408000;
      43503: inst = 32'hc4057d7;
      43504: inst = 32'h8220000;
      43505: inst = 32'h10408000;
      43506: inst = 32'hc4057d8;
      43507: inst = 32'h8220000;
      43508: inst = 32'h10408000;
      43509: inst = 32'hc4057d9;
      43510: inst = 32'h8220000;
      43511: inst = 32'h10408000;
      43512: inst = 32'hc4057da;
      43513: inst = 32'h8220000;
      43514: inst = 32'hc20c344;
      43515: inst = 32'h10408000;
      43516: inst = 32'hc4057db;
      43517: inst = 32'h8220000;
      43518: inst = 32'h58000000;
      43519: inst = 32'h11800000;
      43520: inst = 32'hd800000;
      43521: inst = 32'h11a00000;
      43522: inst = 32'hda00000;
      43523: inst = 32'h25ad5800;
      43524: inst = 32'h15ca6800;
      43525: inst = 32'h21c00001;
      43526: inst = 32'h59200000;
      43527: inst = 32'h298c0001;
      43528: inst = 32'h13e00000;
      43529: inst = 32'hfe0aa03;
      43530: inst = 32'h5be00000;
      43531: inst = 32'h11800000;
      43532: inst = 32'hd800000;
      43533: inst = 32'h258c5800;
      43534: inst = 32'h15aa6000;
      43535: inst = 32'h13e00000;
      43536: inst = 32'hfe0aa16;
      43537: inst = 32'h21a00001;
      43538: inst = 32'h5be00000;
      43539: inst = 32'h13e00000;
      43540: inst = 32'hfe0aa0d;
      43541: inst = 32'h5be00000;
      43542: inst = 32'h2d8c5800;
      43543: inst = 32'h2d8a6000;
      43544: inst = 32'h59200000;
      43545: inst = 32'h11800000;
      43546: inst = 32'hd800000;
      43547: inst = 32'h29ab0000;
      43548: inst = 32'h31ad0001;
      43549: inst = 32'h258c5000;
      43550: inst = 32'h21a00000;
      43551: inst = 32'h59200000;
      43552: inst = 32'h13e00000;
      43553: inst = 32'hfe0aa1c;
      43554: inst = 32'h5be00000;
      43555: inst = 32'hc20ea25;
      43556: inst = 32'h10408000;
      43557: inst = 32'hc404a05;
      43558: inst = 32'h8220000;
      43559: inst = 32'h10408000;
      43560: inst = 32'hc404a06;
      43561: inst = 32'h8220000;
      43562: inst = 32'h10408000;
      43563: inst = 32'hc404a07;
      43564: inst = 32'h8220000;
      43565: inst = 32'h10408000;
      43566: inst = 32'hc404a08;
      43567: inst = 32'h8220000;
      43568: inst = 32'h10408000;
      43569: inst = 32'hc404a09;
      43570: inst = 32'h8220000;
      43571: inst = 32'h10408000;
      43572: inst = 32'hc404a0a;
      43573: inst = 32'h8220000;
      43574: inst = 32'h10408000;
      43575: inst = 32'hc404a0b;
      43576: inst = 32'h8220000;
      43577: inst = 32'h10408000;
      43578: inst = 32'hc404a0c;
      43579: inst = 32'h8220000;
      43580: inst = 32'h10408000;
      43581: inst = 32'hc404a0d;
      43582: inst = 32'h8220000;
      43583: inst = 32'h10408000;
      43584: inst = 32'hc404a0e;
      43585: inst = 32'h8220000;
      43586: inst = 32'h10408000;
      43587: inst = 32'hc404a0f;
      43588: inst = 32'h8220000;
      43589: inst = 32'h10408000;
      43590: inst = 32'hc404a10;
      43591: inst = 32'h8220000;
      43592: inst = 32'h10408000;
      43593: inst = 32'hc404a12;
      43594: inst = 32'h8220000;
      43595: inst = 32'h10408000;
      43596: inst = 32'hc404a13;
      43597: inst = 32'h8220000;
      43598: inst = 32'h10408000;
      43599: inst = 32'hc404a1b;
      43600: inst = 32'h8220000;
      43601: inst = 32'h10408000;
      43602: inst = 32'hc404a1c;
      43603: inst = 32'h8220000;
      43604: inst = 32'h10408000;
      43605: inst = 32'hc404a1f;
      43606: inst = 32'h8220000;
      43607: inst = 32'h10408000;
      43608: inst = 32'hc404a20;
      43609: inst = 32'h8220000;
      43610: inst = 32'h10408000;
      43611: inst = 32'hc404a21;
      43612: inst = 32'h8220000;
      43613: inst = 32'h10408000;
      43614: inst = 32'hc404a22;
      43615: inst = 32'h8220000;
      43616: inst = 32'h10408000;
      43617: inst = 32'hc404a23;
      43618: inst = 32'h8220000;
      43619: inst = 32'h10408000;
      43620: inst = 32'hc404a24;
      43621: inst = 32'h8220000;
      43622: inst = 32'h10408000;
      43623: inst = 32'hc404a25;
      43624: inst = 32'h8220000;
      43625: inst = 32'h10408000;
      43626: inst = 32'hc404a26;
      43627: inst = 32'h8220000;
      43628: inst = 32'h10408000;
      43629: inst = 32'hc404a27;
      43630: inst = 32'h8220000;
      43631: inst = 32'h10408000;
      43632: inst = 32'hc404a28;
      43633: inst = 32'h8220000;
      43634: inst = 32'h10408000;
      43635: inst = 32'hc404a2b;
      43636: inst = 32'h8220000;
      43637: inst = 32'h10408000;
      43638: inst = 32'hc404a2c;
      43639: inst = 32'h8220000;
      43640: inst = 32'h10408000;
      43641: inst = 32'hc404a2d;
      43642: inst = 32'h8220000;
      43643: inst = 32'h10408000;
      43644: inst = 32'hc404a2e;
      43645: inst = 32'h8220000;
      43646: inst = 32'h10408000;
      43647: inst = 32'hc404a2f;
      43648: inst = 32'h8220000;
      43649: inst = 32'h10408000;
      43650: inst = 32'hc404a30;
      43651: inst = 32'h8220000;
      43652: inst = 32'h10408000;
      43653: inst = 32'hc404a31;
      43654: inst = 32'h8220000;
      43655: inst = 32'h10408000;
      43656: inst = 32'hc404a32;
      43657: inst = 32'h8220000;
      43658: inst = 32'h10408000;
      43659: inst = 32'hc404a33;
      43660: inst = 32'h8220000;
      43661: inst = 32'h10408000;
      43662: inst = 32'hc404a34;
      43663: inst = 32'h8220000;
      43664: inst = 32'h10408000;
      43665: inst = 32'hc404a38;
      43666: inst = 32'h8220000;
      43667: inst = 32'h10408000;
      43668: inst = 32'hc404a39;
      43669: inst = 32'h8220000;
      43670: inst = 32'h10408000;
      43671: inst = 32'hc404a3a;
      43672: inst = 32'h8220000;
      43673: inst = 32'h10408000;
      43674: inst = 32'hc404a3b;
      43675: inst = 32'h8220000;
      43676: inst = 32'h10408000;
      43677: inst = 32'hc404a3c;
      43678: inst = 32'h8220000;
      43679: inst = 32'h10408000;
      43680: inst = 32'hc404a3d;
      43681: inst = 32'h8220000;
      43682: inst = 32'h10408000;
      43683: inst = 32'hc404a3e;
      43684: inst = 32'h8220000;
      43685: inst = 32'h10408000;
      43686: inst = 32'hc404a3f;
      43687: inst = 32'h8220000;
      43688: inst = 32'h10408000;
      43689: inst = 32'hc404a40;
      43690: inst = 32'h8220000;
      43691: inst = 32'h10408000;
      43692: inst = 32'hc404a42;
      43693: inst = 32'h8220000;
      43694: inst = 32'h10408000;
      43695: inst = 32'hc404a43;
      43696: inst = 32'h8220000;
      43697: inst = 32'h10408000;
      43698: inst = 32'hc404a44;
      43699: inst = 32'h8220000;
      43700: inst = 32'h10408000;
      43701: inst = 32'hc404a45;
      43702: inst = 32'h8220000;
      43703: inst = 32'h10408000;
      43704: inst = 32'hc404a46;
      43705: inst = 32'h8220000;
      43706: inst = 32'h10408000;
      43707: inst = 32'hc404a47;
      43708: inst = 32'h8220000;
      43709: inst = 32'h10408000;
      43710: inst = 32'hc404a48;
      43711: inst = 32'h8220000;
      43712: inst = 32'h10408000;
      43713: inst = 32'hc404a49;
      43714: inst = 32'h8220000;
      43715: inst = 32'h10408000;
      43716: inst = 32'hc404a4a;
      43717: inst = 32'h8220000;
      43718: inst = 32'h10408000;
      43719: inst = 32'hc404a4b;
      43720: inst = 32'h8220000;
      43721: inst = 32'h10408000;
      43722: inst = 32'hc404a4c;
      43723: inst = 32'h8220000;
      43724: inst = 32'h10408000;
      43725: inst = 32'hc404a4d;
      43726: inst = 32'h8220000;
      43727: inst = 32'h10408000;
      43728: inst = 32'hc404a4f;
      43729: inst = 32'h8220000;
      43730: inst = 32'h10408000;
      43731: inst = 32'hc404a50;
      43732: inst = 32'h8220000;
      43733: inst = 32'h10408000;
      43734: inst = 32'hc404a51;
      43735: inst = 32'h8220000;
      43736: inst = 32'h10408000;
      43737: inst = 32'hc404a52;
      43738: inst = 32'h8220000;
      43739: inst = 32'h10408000;
      43740: inst = 32'hc404a53;
      43741: inst = 32'h8220000;
      43742: inst = 32'h10408000;
      43743: inst = 32'hc404a54;
      43744: inst = 32'h8220000;
      43745: inst = 32'h10408000;
      43746: inst = 32'hc404a55;
      43747: inst = 32'h8220000;
      43748: inst = 32'h10408000;
      43749: inst = 32'hc404a56;
      43750: inst = 32'h8220000;
      43751: inst = 32'h10408000;
      43752: inst = 32'hc404a57;
      43753: inst = 32'h8220000;
      43754: inst = 32'h10408000;
      43755: inst = 32'hc404a58;
      43756: inst = 32'h8220000;
      43757: inst = 32'h10408000;
      43758: inst = 32'hc404a59;
      43759: inst = 32'h8220000;
      43760: inst = 32'h10408000;
      43761: inst = 32'hc404a5a;
      43762: inst = 32'h8220000;
      43763: inst = 32'h10408000;
      43764: inst = 32'hc404a66;
      43765: inst = 32'h8220000;
      43766: inst = 32'h10408000;
      43767: inst = 32'hc404a67;
      43768: inst = 32'h8220000;
      43769: inst = 32'h10408000;
      43770: inst = 32'hc404a68;
      43771: inst = 32'h8220000;
      43772: inst = 32'h10408000;
      43773: inst = 32'hc404a69;
      43774: inst = 32'h8220000;
      43775: inst = 32'h10408000;
      43776: inst = 32'hc404a6a;
      43777: inst = 32'h8220000;
      43778: inst = 32'h10408000;
      43779: inst = 32'hc404a6b;
      43780: inst = 32'h8220000;
      43781: inst = 32'h10408000;
      43782: inst = 32'hc404a6c;
      43783: inst = 32'h8220000;
      43784: inst = 32'h10408000;
      43785: inst = 32'hc404a6d;
      43786: inst = 32'h8220000;
      43787: inst = 32'h10408000;
      43788: inst = 32'hc404a6e;
      43789: inst = 32'h8220000;
      43790: inst = 32'h10408000;
      43791: inst = 32'hc404a6f;
      43792: inst = 32'h8220000;
      43793: inst = 32'h10408000;
      43794: inst = 32'hc404a70;
      43795: inst = 32'h8220000;
      43796: inst = 32'h10408000;
      43797: inst = 32'hc404a72;
      43798: inst = 32'h8220000;
      43799: inst = 32'h10408000;
      43800: inst = 32'hc404a73;
      43801: inst = 32'h8220000;
      43802: inst = 32'h10408000;
      43803: inst = 32'hc404a7b;
      43804: inst = 32'h8220000;
      43805: inst = 32'h10408000;
      43806: inst = 32'hc404a7c;
      43807: inst = 32'h8220000;
      43808: inst = 32'h10408000;
      43809: inst = 32'hc404a7f;
      43810: inst = 32'h8220000;
      43811: inst = 32'h10408000;
      43812: inst = 32'hc404a80;
      43813: inst = 32'h8220000;
      43814: inst = 32'h10408000;
      43815: inst = 32'hc404a81;
      43816: inst = 32'h8220000;
      43817: inst = 32'h10408000;
      43818: inst = 32'hc404a82;
      43819: inst = 32'h8220000;
      43820: inst = 32'h10408000;
      43821: inst = 32'hc404a83;
      43822: inst = 32'h8220000;
      43823: inst = 32'h10408000;
      43824: inst = 32'hc404a84;
      43825: inst = 32'h8220000;
      43826: inst = 32'h10408000;
      43827: inst = 32'hc404a85;
      43828: inst = 32'h8220000;
      43829: inst = 32'h10408000;
      43830: inst = 32'hc404a86;
      43831: inst = 32'h8220000;
      43832: inst = 32'h10408000;
      43833: inst = 32'hc404a87;
      43834: inst = 32'h8220000;
      43835: inst = 32'h10408000;
      43836: inst = 32'hc404a88;
      43837: inst = 32'h8220000;
      43838: inst = 32'h10408000;
      43839: inst = 32'hc404a8b;
      43840: inst = 32'h8220000;
      43841: inst = 32'h10408000;
      43842: inst = 32'hc404a8c;
      43843: inst = 32'h8220000;
      43844: inst = 32'h10408000;
      43845: inst = 32'hc404a8d;
      43846: inst = 32'h8220000;
      43847: inst = 32'h10408000;
      43848: inst = 32'hc404a8e;
      43849: inst = 32'h8220000;
      43850: inst = 32'h10408000;
      43851: inst = 32'hc404a8f;
      43852: inst = 32'h8220000;
      43853: inst = 32'h10408000;
      43854: inst = 32'hc404a90;
      43855: inst = 32'h8220000;
      43856: inst = 32'h10408000;
      43857: inst = 32'hc404a91;
      43858: inst = 32'h8220000;
      43859: inst = 32'h10408000;
      43860: inst = 32'hc404a92;
      43861: inst = 32'h8220000;
      43862: inst = 32'h10408000;
      43863: inst = 32'hc404a93;
      43864: inst = 32'h8220000;
      43865: inst = 32'h10408000;
      43866: inst = 32'hc404a94;
      43867: inst = 32'h8220000;
      43868: inst = 32'h10408000;
      43869: inst = 32'hc404a97;
      43870: inst = 32'h8220000;
      43871: inst = 32'h10408000;
      43872: inst = 32'hc404a98;
      43873: inst = 32'h8220000;
      43874: inst = 32'h10408000;
      43875: inst = 32'hc404a99;
      43876: inst = 32'h8220000;
      43877: inst = 32'h10408000;
      43878: inst = 32'hc404a9a;
      43879: inst = 32'h8220000;
      43880: inst = 32'h10408000;
      43881: inst = 32'hc404a9b;
      43882: inst = 32'h8220000;
      43883: inst = 32'h10408000;
      43884: inst = 32'hc404a9c;
      43885: inst = 32'h8220000;
      43886: inst = 32'h10408000;
      43887: inst = 32'hc404a9d;
      43888: inst = 32'h8220000;
      43889: inst = 32'h10408000;
      43890: inst = 32'hc404a9e;
      43891: inst = 32'h8220000;
      43892: inst = 32'h10408000;
      43893: inst = 32'hc404a9f;
      43894: inst = 32'h8220000;
      43895: inst = 32'h10408000;
      43896: inst = 32'hc404aa0;
      43897: inst = 32'h8220000;
      43898: inst = 32'h10408000;
      43899: inst = 32'hc404aa3;
      43900: inst = 32'h8220000;
      43901: inst = 32'h10408000;
      43902: inst = 32'hc404aa4;
      43903: inst = 32'h8220000;
      43904: inst = 32'h10408000;
      43905: inst = 32'hc404aa5;
      43906: inst = 32'h8220000;
      43907: inst = 32'h10408000;
      43908: inst = 32'hc404aa6;
      43909: inst = 32'h8220000;
      43910: inst = 32'h10408000;
      43911: inst = 32'hc404aa7;
      43912: inst = 32'h8220000;
      43913: inst = 32'h10408000;
      43914: inst = 32'hc404aa8;
      43915: inst = 32'h8220000;
      43916: inst = 32'h10408000;
      43917: inst = 32'hc404aa9;
      43918: inst = 32'h8220000;
      43919: inst = 32'h10408000;
      43920: inst = 32'hc404aaa;
      43921: inst = 32'h8220000;
      43922: inst = 32'h10408000;
      43923: inst = 32'hc404aab;
      43924: inst = 32'h8220000;
      43925: inst = 32'h10408000;
      43926: inst = 32'hc404aac;
      43927: inst = 32'h8220000;
      43928: inst = 32'h10408000;
      43929: inst = 32'hc404aad;
      43930: inst = 32'h8220000;
      43931: inst = 32'h10408000;
      43932: inst = 32'hc404ab0;
      43933: inst = 32'h8220000;
      43934: inst = 32'h10408000;
      43935: inst = 32'hc404ab1;
      43936: inst = 32'h8220000;
      43937: inst = 32'h10408000;
      43938: inst = 32'hc404ab2;
      43939: inst = 32'h8220000;
      43940: inst = 32'h10408000;
      43941: inst = 32'hc404ab3;
      43942: inst = 32'h8220000;
      43943: inst = 32'h10408000;
      43944: inst = 32'hc404ab4;
      43945: inst = 32'h8220000;
      43946: inst = 32'h10408000;
      43947: inst = 32'hc404ab5;
      43948: inst = 32'h8220000;
      43949: inst = 32'h10408000;
      43950: inst = 32'hc404ab6;
      43951: inst = 32'h8220000;
      43952: inst = 32'h10408000;
      43953: inst = 32'hc404ab7;
      43954: inst = 32'h8220000;
      43955: inst = 32'h10408000;
      43956: inst = 32'hc404ab8;
      43957: inst = 32'h8220000;
      43958: inst = 32'h10408000;
      43959: inst = 32'hc404ab9;
      43960: inst = 32'h8220000;
      43961: inst = 32'h10408000;
      43962: inst = 32'hc404aba;
      43963: inst = 32'h8220000;
      43964: inst = 32'h10408000;
      43965: inst = 32'hc404ac7;
      43966: inst = 32'h8220000;
      43967: inst = 32'h10408000;
      43968: inst = 32'hc404ac8;
      43969: inst = 32'h8220000;
      43970: inst = 32'h10408000;
      43971: inst = 32'hc404ac9;
      43972: inst = 32'h8220000;
      43973: inst = 32'h10408000;
      43974: inst = 32'hc404aca;
      43975: inst = 32'h8220000;
      43976: inst = 32'h10408000;
      43977: inst = 32'hc404ad2;
      43978: inst = 32'h8220000;
      43979: inst = 32'h10408000;
      43980: inst = 32'hc404ad3;
      43981: inst = 32'h8220000;
      43982: inst = 32'h10408000;
      43983: inst = 32'hc404adb;
      43984: inst = 32'h8220000;
      43985: inst = 32'h10408000;
      43986: inst = 32'hc404adc;
      43987: inst = 32'h8220000;
      43988: inst = 32'h10408000;
      43989: inst = 32'hc404adf;
      43990: inst = 32'h8220000;
      43991: inst = 32'h10408000;
      43992: inst = 32'hc404ae0;
      43993: inst = 32'h8220000;
      43994: inst = 32'h10408000;
      43995: inst = 32'hc404ae7;
      43996: inst = 32'h8220000;
      43997: inst = 32'h10408000;
      43998: inst = 32'hc404ae8;
      43999: inst = 32'h8220000;
      44000: inst = 32'h10408000;
      44001: inst = 32'hc404aeb;
      44002: inst = 32'h8220000;
      44003: inst = 32'h10408000;
      44004: inst = 32'hc404aec;
      44005: inst = 32'h8220000;
      44006: inst = 32'h10408000;
      44007: inst = 32'hc404af3;
      44008: inst = 32'h8220000;
      44009: inst = 32'h10408000;
      44010: inst = 32'hc404af4;
      44011: inst = 32'h8220000;
      44012: inst = 32'h10408000;
      44013: inst = 32'hc404af6;
      44014: inst = 32'h8220000;
      44015: inst = 32'h10408000;
      44016: inst = 32'hc404af7;
      44017: inst = 32'h8220000;
      44018: inst = 32'h10408000;
      44019: inst = 32'hc404af8;
      44020: inst = 32'h8220000;
      44021: inst = 32'h10408000;
      44022: inst = 32'hc404b04;
      44023: inst = 32'h8220000;
      44024: inst = 32'h10408000;
      44025: inst = 32'hc404b05;
      44026: inst = 32'h8220000;
      44027: inst = 32'h10408000;
      44028: inst = 32'hc404b06;
      44029: inst = 32'h8220000;
      44030: inst = 32'h10408000;
      44031: inst = 32'hc404b07;
      44032: inst = 32'h8220000;
      44033: inst = 32'h10408000;
      44034: inst = 32'hc404b11;
      44035: inst = 32'h8220000;
      44036: inst = 32'h10408000;
      44037: inst = 32'hc404b12;
      44038: inst = 32'h8220000;
      44039: inst = 32'h10408000;
      44040: inst = 32'hc404b13;
      44041: inst = 32'h8220000;
      44042: inst = 32'h10408000;
      44043: inst = 32'hc404b14;
      44044: inst = 32'h8220000;
      44045: inst = 32'h10408000;
      44046: inst = 32'hc404b28;
      44047: inst = 32'h8220000;
      44048: inst = 32'h10408000;
      44049: inst = 32'hc404b29;
      44050: inst = 32'h8220000;
      44051: inst = 32'h10408000;
      44052: inst = 32'hc404b2a;
      44053: inst = 32'h8220000;
      44054: inst = 32'h10408000;
      44055: inst = 32'hc404b32;
      44056: inst = 32'h8220000;
      44057: inst = 32'h10408000;
      44058: inst = 32'hc404b33;
      44059: inst = 32'h8220000;
      44060: inst = 32'h10408000;
      44061: inst = 32'hc404b3b;
      44062: inst = 32'h8220000;
      44063: inst = 32'h10408000;
      44064: inst = 32'hc404b3c;
      44065: inst = 32'h8220000;
      44066: inst = 32'h10408000;
      44067: inst = 32'hc404b3f;
      44068: inst = 32'h8220000;
      44069: inst = 32'h10408000;
      44070: inst = 32'hc404b40;
      44071: inst = 32'h8220000;
      44072: inst = 32'h10408000;
      44073: inst = 32'hc404b47;
      44074: inst = 32'h8220000;
      44075: inst = 32'h10408000;
      44076: inst = 32'hc404b48;
      44077: inst = 32'h8220000;
      44078: inst = 32'h10408000;
      44079: inst = 32'hc404b4b;
      44080: inst = 32'h8220000;
      44081: inst = 32'h10408000;
      44082: inst = 32'hc404b4c;
      44083: inst = 32'h8220000;
      44084: inst = 32'h10408000;
      44085: inst = 32'hc404b53;
      44086: inst = 32'h8220000;
      44087: inst = 32'h10408000;
      44088: inst = 32'hc404b54;
      44089: inst = 32'h8220000;
      44090: inst = 32'h10408000;
      44091: inst = 32'hc404b56;
      44092: inst = 32'h8220000;
      44093: inst = 32'h10408000;
      44094: inst = 32'hc404b57;
      44095: inst = 32'h8220000;
      44096: inst = 32'h10408000;
      44097: inst = 32'hc404b65;
      44098: inst = 32'h8220000;
      44099: inst = 32'h10408000;
      44100: inst = 32'hc404b66;
      44101: inst = 32'h8220000;
      44102: inst = 32'h10408000;
      44103: inst = 32'hc404b67;
      44104: inst = 32'h8220000;
      44105: inst = 32'h10408000;
      44106: inst = 32'hc404b72;
      44107: inst = 32'h8220000;
      44108: inst = 32'h10408000;
      44109: inst = 32'hc404b73;
      44110: inst = 32'h8220000;
      44111: inst = 32'h10408000;
      44112: inst = 32'hc404b74;
      44113: inst = 32'h8220000;
      44114: inst = 32'h10408000;
      44115: inst = 32'hc404b89;
      44116: inst = 32'h8220000;
      44117: inst = 32'h10408000;
      44118: inst = 32'hc404b8a;
      44119: inst = 32'h8220000;
      44120: inst = 32'h10408000;
      44121: inst = 32'hc404b8b;
      44122: inst = 32'h8220000;
      44123: inst = 32'h10408000;
      44124: inst = 32'hc404b92;
      44125: inst = 32'h8220000;
      44126: inst = 32'h10408000;
      44127: inst = 32'hc404b93;
      44128: inst = 32'h8220000;
      44129: inst = 32'h10408000;
      44130: inst = 32'hc404b94;
      44131: inst = 32'h8220000;
      44132: inst = 32'h10408000;
      44133: inst = 32'hc404b9b;
      44134: inst = 32'h8220000;
      44135: inst = 32'h10408000;
      44136: inst = 32'hc404b9c;
      44137: inst = 32'h8220000;
      44138: inst = 32'h10408000;
      44139: inst = 32'hc404b9f;
      44140: inst = 32'h8220000;
      44141: inst = 32'h10408000;
      44142: inst = 32'hc404ba0;
      44143: inst = 32'h8220000;
      44144: inst = 32'h10408000;
      44145: inst = 32'hc404ba7;
      44146: inst = 32'h8220000;
      44147: inst = 32'h10408000;
      44148: inst = 32'hc404bab;
      44149: inst = 32'h8220000;
      44150: inst = 32'h10408000;
      44151: inst = 32'hc404bac;
      44152: inst = 32'h8220000;
      44153: inst = 32'h10408000;
      44154: inst = 32'hc404bb3;
      44155: inst = 32'h8220000;
      44156: inst = 32'h10408000;
      44157: inst = 32'hc404bb6;
      44158: inst = 32'h8220000;
      44159: inst = 32'h10408000;
      44160: inst = 32'hc404bb7;
      44161: inst = 32'h8220000;
      44162: inst = 32'h10408000;
      44163: inst = 32'hc404bb9;
      44164: inst = 32'h8220000;
      44165: inst = 32'h10408000;
      44166: inst = 32'hc404bba;
      44167: inst = 32'h8220000;
      44168: inst = 32'h10408000;
      44169: inst = 32'hc404bbb;
      44170: inst = 32'h8220000;
      44171: inst = 32'h10408000;
      44172: inst = 32'hc404bbc;
      44173: inst = 32'h8220000;
      44174: inst = 32'h10408000;
      44175: inst = 32'hc404bbd;
      44176: inst = 32'h8220000;
      44177: inst = 32'h10408000;
      44178: inst = 32'hc404bc6;
      44179: inst = 32'h8220000;
      44180: inst = 32'h10408000;
      44181: inst = 32'hc404bc7;
      44182: inst = 32'h8220000;
      44183: inst = 32'h10408000;
      44184: inst = 32'hc404bc8;
      44185: inst = 32'h8220000;
      44186: inst = 32'h10408000;
      44187: inst = 32'hc404bd3;
      44188: inst = 32'h8220000;
      44189: inst = 32'h10408000;
      44190: inst = 32'hc404bd4;
      44191: inst = 32'h8220000;
      44192: inst = 32'h10408000;
      44193: inst = 32'hc404bd5;
      44194: inst = 32'h8220000;
      44195: inst = 32'h10408000;
      44196: inst = 32'hc404bea;
      44197: inst = 32'h8220000;
      44198: inst = 32'h10408000;
      44199: inst = 32'hc404beb;
      44200: inst = 32'h8220000;
      44201: inst = 32'h10408000;
      44202: inst = 32'hc404bec;
      44203: inst = 32'h8220000;
      44204: inst = 32'h10408000;
      44205: inst = 32'hc404bf3;
      44206: inst = 32'h8220000;
      44207: inst = 32'h10408000;
      44208: inst = 32'hc404bf4;
      44209: inst = 32'h8220000;
      44210: inst = 32'h10408000;
      44211: inst = 32'hc404bf5;
      44212: inst = 32'h8220000;
      44213: inst = 32'h10408000;
      44214: inst = 32'hc404bfb;
      44215: inst = 32'h8220000;
      44216: inst = 32'h10408000;
      44217: inst = 32'hc404bfc;
      44218: inst = 32'h8220000;
      44219: inst = 32'h10408000;
      44220: inst = 32'hc404bff;
      44221: inst = 32'h8220000;
      44222: inst = 32'h10408000;
      44223: inst = 32'hc404c00;
      44224: inst = 32'h8220000;
      44225: inst = 32'h10408000;
      44226: inst = 32'hc404c0b;
      44227: inst = 32'h8220000;
      44228: inst = 32'h10408000;
      44229: inst = 32'hc404c0c;
      44230: inst = 32'h8220000;
      44231: inst = 32'h10408000;
      44232: inst = 32'hc404c16;
      44233: inst = 32'h8220000;
      44234: inst = 32'h10408000;
      44235: inst = 32'hc404c17;
      44236: inst = 32'h8220000;
      44237: inst = 32'h10408000;
      44238: inst = 32'hc404c19;
      44239: inst = 32'h8220000;
      44240: inst = 32'h10408000;
      44241: inst = 32'hc404c1a;
      44242: inst = 32'h8220000;
      44243: inst = 32'h10408000;
      44244: inst = 32'hc404c1b;
      44245: inst = 32'h8220000;
      44246: inst = 32'h10408000;
      44247: inst = 32'hc404c1c;
      44248: inst = 32'h8220000;
      44249: inst = 32'h10408000;
      44250: inst = 32'hc404c1d;
      44251: inst = 32'h8220000;
      44252: inst = 32'h10408000;
      44253: inst = 32'hc404c27;
      44254: inst = 32'h8220000;
      44255: inst = 32'h10408000;
      44256: inst = 32'hc404c28;
      44257: inst = 32'h8220000;
      44258: inst = 32'h10408000;
      44259: inst = 32'hc404c29;
      44260: inst = 32'h8220000;
      44261: inst = 32'h10408000;
      44262: inst = 32'hc404c34;
      44263: inst = 32'h8220000;
      44264: inst = 32'h10408000;
      44265: inst = 32'hc404c35;
      44266: inst = 32'h8220000;
      44267: inst = 32'h10408000;
      44268: inst = 32'hc404c36;
      44269: inst = 32'h8220000;
      44270: inst = 32'h10408000;
      44271: inst = 32'hc404c4b;
      44272: inst = 32'h8220000;
      44273: inst = 32'h10408000;
      44274: inst = 32'hc404c4c;
      44275: inst = 32'h8220000;
      44276: inst = 32'h10408000;
      44277: inst = 32'hc404c4d;
      44278: inst = 32'h8220000;
      44279: inst = 32'h10408000;
      44280: inst = 32'hc404c54;
      44281: inst = 32'h8220000;
      44282: inst = 32'h10408000;
      44283: inst = 32'hc404c55;
      44284: inst = 32'h8220000;
      44285: inst = 32'h10408000;
      44286: inst = 32'hc404c56;
      44287: inst = 32'h8220000;
      44288: inst = 32'h10408000;
      44289: inst = 32'hc404c5b;
      44290: inst = 32'h8220000;
      44291: inst = 32'h10408000;
      44292: inst = 32'hc404c5c;
      44293: inst = 32'h8220000;
      44294: inst = 32'h10408000;
      44295: inst = 32'hc404c5f;
      44296: inst = 32'h8220000;
      44297: inst = 32'h10408000;
      44298: inst = 32'hc404c60;
      44299: inst = 32'h8220000;
      44300: inst = 32'h10408000;
      44301: inst = 32'hc404c6b;
      44302: inst = 32'h8220000;
      44303: inst = 32'h10408000;
      44304: inst = 32'hc404c6c;
      44305: inst = 32'h8220000;
      44306: inst = 32'h10408000;
      44307: inst = 32'hc404c76;
      44308: inst = 32'h8220000;
      44309: inst = 32'h10408000;
      44310: inst = 32'hc404c77;
      44311: inst = 32'h8220000;
      44312: inst = 32'h10408000;
      44313: inst = 32'hc404c88;
      44314: inst = 32'h8220000;
      44315: inst = 32'h10408000;
      44316: inst = 32'hc404c89;
      44317: inst = 32'h8220000;
      44318: inst = 32'h10408000;
      44319: inst = 32'hc404c8a;
      44320: inst = 32'h8220000;
      44321: inst = 32'h10408000;
      44322: inst = 32'hc404c95;
      44323: inst = 32'h8220000;
      44324: inst = 32'h10408000;
      44325: inst = 32'hc404c96;
      44326: inst = 32'h8220000;
      44327: inst = 32'h10408000;
      44328: inst = 32'hc404c97;
      44329: inst = 32'h8220000;
      44330: inst = 32'h10408000;
      44331: inst = 32'hc404ca5;
      44332: inst = 32'h8220000;
      44333: inst = 32'h10408000;
      44334: inst = 32'hc404ca6;
      44335: inst = 32'h8220000;
      44336: inst = 32'h10408000;
      44337: inst = 32'hc404ca7;
      44338: inst = 32'h8220000;
      44339: inst = 32'h10408000;
      44340: inst = 32'hc404ca8;
      44341: inst = 32'h8220000;
      44342: inst = 32'h10408000;
      44343: inst = 32'hc404ca9;
      44344: inst = 32'h8220000;
      44345: inst = 32'h10408000;
      44346: inst = 32'hc404caa;
      44347: inst = 32'h8220000;
      44348: inst = 32'h10408000;
      44349: inst = 32'hc404cab;
      44350: inst = 32'h8220000;
      44351: inst = 32'h10408000;
      44352: inst = 32'hc404cac;
      44353: inst = 32'h8220000;
      44354: inst = 32'h10408000;
      44355: inst = 32'hc404cad;
      44356: inst = 32'h8220000;
      44357: inst = 32'h10408000;
      44358: inst = 32'hc404cae;
      44359: inst = 32'h8220000;
      44360: inst = 32'h10408000;
      44361: inst = 32'hc404cb5;
      44362: inst = 32'h8220000;
      44363: inst = 32'h10408000;
      44364: inst = 32'hc404cb6;
      44365: inst = 32'h8220000;
      44366: inst = 32'h10408000;
      44367: inst = 32'hc404cb7;
      44368: inst = 32'h8220000;
      44369: inst = 32'h10408000;
      44370: inst = 32'hc404cb8;
      44371: inst = 32'h8220000;
      44372: inst = 32'h10408000;
      44373: inst = 32'hc404cb9;
      44374: inst = 32'h8220000;
      44375: inst = 32'h10408000;
      44376: inst = 32'hc404cba;
      44377: inst = 32'h8220000;
      44378: inst = 32'h10408000;
      44379: inst = 32'hc404cbb;
      44380: inst = 32'h8220000;
      44381: inst = 32'h10408000;
      44382: inst = 32'hc404cbc;
      44383: inst = 32'h8220000;
      44384: inst = 32'h10408000;
      44385: inst = 32'hc404cbf;
      44386: inst = 32'h8220000;
      44387: inst = 32'h10408000;
      44388: inst = 32'hc404cc0;
      44389: inst = 32'h8220000;
      44390: inst = 32'h10408000;
      44391: inst = 32'hc404cc1;
      44392: inst = 32'h8220000;
      44393: inst = 32'h10408000;
      44394: inst = 32'hc404cc2;
      44395: inst = 32'h8220000;
      44396: inst = 32'h10408000;
      44397: inst = 32'hc404cc3;
      44398: inst = 32'h8220000;
      44399: inst = 32'h10408000;
      44400: inst = 32'hc404cc4;
      44401: inst = 32'h8220000;
      44402: inst = 32'h10408000;
      44403: inst = 32'hc404cc5;
      44404: inst = 32'h8220000;
      44405: inst = 32'h10408000;
      44406: inst = 32'hc404cc6;
      44407: inst = 32'h8220000;
      44408: inst = 32'h10408000;
      44409: inst = 32'hc404cc7;
      44410: inst = 32'h8220000;
      44411: inst = 32'h10408000;
      44412: inst = 32'hc404cc8;
      44413: inst = 32'h8220000;
      44414: inst = 32'h10408000;
      44415: inst = 32'hc404ccb;
      44416: inst = 32'h8220000;
      44417: inst = 32'h10408000;
      44418: inst = 32'hc404ccc;
      44419: inst = 32'h8220000;
      44420: inst = 32'h10408000;
      44421: inst = 32'hc404ccd;
      44422: inst = 32'h8220000;
      44423: inst = 32'h10408000;
      44424: inst = 32'hc404cce;
      44425: inst = 32'h8220000;
      44426: inst = 32'h10408000;
      44427: inst = 32'hc404ccf;
      44428: inst = 32'h8220000;
      44429: inst = 32'h10408000;
      44430: inst = 32'hc404cd0;
      44431: inst = 32'h8220000;
      44432: inst = 32'h10408000;
      44433: inst = 32'hc404cd1;
      44434: inst = 32'h8220000;
      44435: inst = 32'h10408000;
      44436: inst = 32'hc404cd2;
      44437: inst = 32'h8220000;
      44438: inst = 32'h10408000;
      44439: inst = 32'hc404cd3;
      44440: inst = 32'h8220000;
      44441: inst = 32'h10408000;
      44442: inst = 32'hc404cd4;
      44443: inst = 32'h8220000;
      44444: inst = 32'h10408000;
      44445: inst = 32'hc404cd5;
      44446: inst = 32'h8220000;
      44447: inst = 32'h10408000;
      44448: inst = 32'hc404cd6;
      44449: inst = 32'h8220000;
      44450: inst = 32'h10408000;
      44451: inst = 32'hc404cd7;
      44452: inst = 32'h8220000;
      44453: inst = 32'h10408000;
      44454: inst = 32'hc404cd8;
      44455: inst = 32'h8220000;
      44456: inst = 32'h10408000;
      44457: inst = 32'hc404cd9;
      44458: inst = 32'h8220000;
      44459: inst = 32'h10408000;
      44460: inst = 32'hc404cda;
      44461: inst = 32'h8220000;
      44462: inst = 32'h10408000;
      44463: inst = 32'hc404cdb;
      44464: inst = 32'h8220000;
      44465: inst = 32'h10408000;
      44466: inst = 32'hc404cdc;
      44467: inst = 32'h8220000;
      44468: inst = 32'h10408000;
      44469: inst = 32'hc404cdd;
      44470: inst = 32'h8220000;
      44471: inst = 32'h10408000;
      44472: inst = 32'hc404cde;
      44473: inst = 32'h8220000;
      44474: inst = 32'h10408000;
      44475: inst = 32'hc404cdf;
      44476: inst = 32'h8220000;
      44477: inst = 32'h10408000;
      44478: inst = 32'hc404ce0;
      44479: inst = 32'h8220000;
      44480: inst = 32'h10408000;
      44481: inst = 32'hc404ce2;
      44482: inst = 32'h8220000;
      44483: inst = 32'h10408000;
      44484: inst = 32'hc404ce3;
      44485: inst = 32'h8220000;
      44486: inst = 32'h10408000;
      44487: inst = 32'hc404ce4;
      44488: inst = 32'h8220000;
      44489: inst = 32'h10408000;
      44490: inst = 32'hc404ce5;
      44491: inst = 32'h8220000;
      44492: inst = 32'h10408000;
      44493: inst = 32'hc404ce6;
      44494: inst = 32'h8220000;
      44495: inst = 32'h10408000;
      44496: inst = 32'hc404ce7;
      44497: inst = 32'h8220000;
      44498: inst = 32'h10408000;
      44499: inst = 32'hc404ce8;
      44500: inst = 32'h8220000;
      44501: inst = 32'h10408000;
      44502: inst = 32'hc404ce9;
      44503: inst = 32'h8220000;
      44504: inst = 32'h10408000;
      44505: inst = 32'hc404cea;
      44506: inst = 32'h8220000;
      44507: inst = 32'h10408000;
      44508: inst = 32'hc404ceb;
      44509: inst = 32'h8220000;
      44510: inst = 32'h10408000;
      44511: inst = 32'hc404cef;
      44512: inst = 32'h8220000;
      44513: inst = 32'h10408000;
      44514: inst = 32'hc404cf0;
      44515: inst = 32'h8220000;
      44516: inst = 32'h10408000;
      44517: inst = 32'hc404cf1;
      44518: inst = 32'h8220000;
      44519: inst = 32'h10408000;
      44520: inst = 32'hc404cf2;
      44521: inst = 32'h8220000;
      44522: inst = 32'h10408000;
      44523: inst = 32'hc404cf3;
      44524: inst = 32'h8220000;
      44525: inst = 32'h10408000;
      44526: inst = 32'hc404cf4;
      44527: inst = 32'h8220000;
      44528: inst = 32'h10408000;
      44529: inst = 32'hc404cf5;
      44530: inst = 32'h8220000;
      44531: inst = 32'h10408000;
      44532: inst = 32'hc404cf6;
      44533: inst = 32'h8220000;
      44534: inst = 32'h10408000;
      44535: inst = 32'hc404cf7;
      44536: inst = 32'h8220000;
      44537: inst = 32'h10408000;
      44538: inst = 32'hc404cf8;
      44539: inst = 32'h8220000;
      44540: inst = 32'h10408000;
      44541: inst = 32'hc404d05;
      44542: inst = 32'h8220000;
      44543: inst = 32'h10408000;
      44544: inst = 32'hc404d06;
      44545: inst = 32'h8220000;
      44546: inst = 32'h10408000;
      44547: inst = 32'hc404d07;
      44548: inst = 32'h8220000;
      44549: inst = 32'h10408000;
      44550: inst = 32'hc404d08;
      44551: inst = 32'h8220000;
      44552: inst = 32'h10408000;
      44553: inst = 32'hc404d09;
      44554: inst = 32'h8220000;
      44555: inst = 32'h10408000;
      44556: inst = 32'hc404d0a;
      44557: inst = 32'h8220000;
      44558: inst = 32'h10408000;
      44559: inst = 32'hc404d0b;
      44560: inst = 32'h8220000;
      44561: inst = 32'h10408000;
      44562: inst = 32'hc404d0c;
      44563: inst = 32'h8220000;
      44564: inst = 32'h10408000;
      44565: inst = 32'hc404d0d;
      44566: inst = 32'h8220000;
      44567: inst = 32'h10408000;
      44568: inst = 32'hc404d0e;
      44569: inst = 32'h8220000;
      44570: inst = 32'h10408000;
      44571: inst = 32'hc404d0f;
      44572: inst = 32'h8220000;
      44573: inst = 32'h10408000;
      44574: inst = 32'hc404d16;
      44575: inst = 32'h8220000;
      44576: inst = 32'h10408000;
      44577: inst = 32'hc404d17;
      44578: inst = 32'h8220000;
      44579: inst = 32'h10408000;
      44580: inst = 32'hc404d18;
      44581: inst = 32'h8220000;
      44582: inst = 32'h10408000;
      44583: inst = 32'hc404d19;
      44584: inst = 32'h8220000;
      44585: inst = 32'h10408000;
      44586: inst = 32'hc404d1a;
      44587: inst = 32'h8220000;
      44588: inst = 32'h10408000;
      44589: inst = 32'hc404d1b;
      44590: inst = 32'h8220000;
      44591: inst = 32'h10408000;
      44592: inst = 32'hc404d1c;
      44593: inst = 32'h8220000;
      44594: inst = 32'h10408000;
      44595: inst = 32'hc404d20;
      44596: inst = 32'h8220000;
      44597: inst = 32'h10408000;
      44598: inst = 32'hc404d21;
      44599: inst = 32'h8220000;
      44600: inst = 32'h10408000;
      44601: inst = 32'hc404d22;
      44602: inst = 32'h8220000;
      44603: inst = 32'h10408000;
      44604: inst = 32'hc404d23;
      44605: inst = 32'h8220000;
      44606: inst = 32'h10408000;
      44607: inst = 32'hc404d24;
      44608: inst = 32'h8220000;
      44609: inst = 32'h10408000;
      44610: inst = 32'hc404d25;
      44611: inst = 32'h8220000;
      44612: inst = 32'h10408000;
      44613: inst = 32'hc404d26;
      44614: inst = 32'h8220000;
      44615: inst = 32'h10408000;
      44616: inst = 32'hc404d27;
      44617: inst = 32'h8220000;
      44618: inst = 32'h10408000;
      44619: inst = 32'hc404d28;
      44620: inst = 32'h8220000;
      44621: inst = 32'h10408000;
      44622: inst = 32'hc404d2c;
      44623: inst = 32'h8220000;
      44624: inst = 32'h10408000;
      44625: inst = 32'hc404d2d;
      44626: inst = 32'h8220000;
      44627: inst = 32'h10408000;
      44628: inst = 32'hc404d2e;
      44629: inst = 32'h8220000;
      44630: inst = 32'h10408000;
      44631: inst = 32'hc404d2f;
      44632: inst = 32'h8220000;
      44633: inst = 32'h10408000;
      44634: inst = 32'hc404d30;
      44635: inst = 32'h8220000;
      44636: inst = 32'h10408000;
      44637: inst = 32'hc404d31;
      44638: inst = 32'h8220000;
      44639: inst = 32'h10408000;
      44640: inst = 32'hc404d32;
      44641: inst = 32'h8220000;
      44642: inst = 32'h10408000;
      44643: inst = 32'hc404d33;
      44644: inst = 32'h8220000;
      44645: inst = 32'h10408000;
      44646: inst = 32'hc404d34;
      44647: inst = 32'h8220000;
      44648: inst = 32'h10408000;
      44649: inst = 32'hc404d35;
      44650: inst = 32'h8220000;
      44651: inst = 32'h10408000;
      44652: inst = 32'hc404d36;
      44653: inst = 32'h8220000;
      44654: inst = 32'h10408000;
      44655: inst = 32'hc404d37;
      44656: inst = 32'h8220000;
      44657: inst = 32'h10408000;
      44658: inst = 32'hc404d38;
      44659: inst = 32'h8220000;
      44660: inst = 32'h10408000;
      44661: inst = 32'hc404d39;
      44662: inst = 32'h8220000;
      44663: inst = 32'h10408000;
      44664: inst = 32'hc404d3a;
      44665: inst = 32'h8220000;
      44666: inst = 32'h10408000;
      44667: inst = 32'hc404d3b;
      44668: inst = 32'h8220000;
      44669: inst = 32'h10408000;
      44670: inst = 32'hc404d3c;
      44671: inst = 32'h8220000;
      44672: inst = 32'h10408000;
      44673: inst = 32'hc404d3d;
      44674: inst = 32'h8220000;
      44675: inst = 32'h10408000;
      44676: inst = 32'hc404d3e;
      44677: inst = 32'h8220000;
      44678: inst = 32'h10408000;
      44679: inst = 32'hc404d3f;
      44680: inst = 32'h8220000;
      44681: inst = 32'h10408000;
      44682: inst = 32'hc404d42;
      44683: inst = 32'h8220000;
      44684: inst = 32'h10408000;
      44685: inst = 32'hc404d43;
      44686: inst = 32'h8220000;
      44687: inst = 32'h10408000;
      44688: inst = 32'hc404d44;
      44689: inst = 32'h8220000;
      44690: inst = 32'h10408000;
      44691: inst = 32'hc404d45;
      44692: inst = 32'h8220000;
      44693: inst = 32'h10408000;
      44694: inst = 32'hc404d46;
      44695: inst = 32'h8220000;
      44696: inst = 32'h10408000;
      44697: inst = 32'hc404d47;
      44698: inst = 32'h8220000;
      44699: inst = 32'h10408000;
      44700: inst = 32'hc404d48;
      44701: inst = 32'h8220000;
      44702: inst = 32'h10408000;
      44703: inst = 32'hc404d49;
      44704: inst = 32'h8220000;
      44705: inst = 32'h10408000;
      44706: inst = 32'hc404d4a;
      44707: inst = 32'h8220000;
      44708: inst = 32'h10408000;
      44709: inst = 32'hc404d4b;
      44710: inst = 32'h8220000;
      44711: inst = 32'h10408000;
      44712: inst = 32'hc404d4c;
      44713: inst = 32'h8220000;
      44714: inst = 32'h10408000;
      44715: inst = 32'hc404d4f;
      44716: inst = 32'h8220000;
      44717: inst = 32'h10408000;
      44718: inst = 32'hc404d50;
      44719: inst = 32'h8220000;
      44720: inst = 32'h10408000;
      44721: inst = 32'hc404d51;
      44722: inst = 32'h8220000;
      44723: inst = 32'h10408000;
      44724: inst = 32'hc404d52;
      44725: inst = 32'h8220000;
      44726: inst = 32'h10408000;
      44727: inst = 32'hc404d53;
      44728: inst = 32'h8220000;
      44729: inst = 32'h10408000;
      44730: inst = 32'hc404d54;
      44731: inst = 32'h8220000;
      44732: inst = 32'h10408000;
      44733: inst = 32'hc404d55;
      44734: inst = 32'h8220000;
      44735: inst = 32'h10408000;
      44736: inst = 32'hc404d56;
      44737: inst = 32'h8220000;
      44738: inst = 32'h10408000;
      44739: inst = 32'hc404d57;
      44740: inst = 32'h8220000;
      44741: inst = 32'h10408000;
      44742: inst = 32'hc404d58;
      44743: inst = 32'h8220000;
      44744: inst = 32'h10408000;
      44745: inst = 32'hc404d59;
      44746: inst = 32'h8220000;
      44747: inst = 32'h58000000;
      44748: inst = 32'hc20ea25;
      44749: inst = 32'h10408000;
      44750: inst = 32'hc404a1d;
      44751: inst = 32'h8220000;
      44752: inst = 32'h10408000;
      44753: inst = 32'hc404a1e;
      44754: inst = 32'h8220000;
      44755: inst = 32'h10408000;
      44756: inst = 32'hc404a1f;
      44757: inst = 32'h8220000;
      44758: inst = 32'h10408000;
      44759: inst = 32'hc404a20;
      44760: inst = 32'h8220000;
      44761: inst = 32'h10408000;
      44762: inst = 32'hc404a21;
      44763: inst = 32'h8220000;
      44764: inst = 32'h10408000;
      44765: inst = 32'hc404a22;
      44766: inst = 32'h8220000;
      44767: inst = 32'h10408000;
      44768: inst = 32'hc404a23;
      44769: inst = 32'h8220000;
      44770: inst = 32'h10408000;
      44771: inst = 32'hc404a24;
      44772: inst = 32'h8220000;
      44773: inst = 32'h10408000;
      44774: inst = 32'hc404a25;
      44775: inst = 32'h8220000;
      44776: inst = 32'h10408000;
      44777: inst = 32'hc404a26;
      44778: inst = 32'h8220000;
      44779: inst = 32'h10408000;
      44780: inst = 32'hc404a27;
      44781: inst = 32'h8220000;
      44782: inst = 32'h10408000;
      44783: inst = 32'hc404a2a;
      44784: inst = 32'h8220000;
      44785: inst = 32'h10408000;
      44786: inst = 32'hc404a2b;
      44787: inst = 32'h8220000;
      44788: inst = 32'h10408000;
      44789: inst = 32'hc404a2c;
      44790: inst = 32'h8220000;
      44791: inst = 32'h10408000;
      44792: inst = 32'hc404a36;
      44793: inst = 32'h8220000;
      44794: inst = 32'h10408000;
      44795: inst = 32'hc404a37;
      44796: inst = 32'h8220000;
      44797: inst = 32'h10408000;
      44798: inst = 32'hc404a3a;
      44799: inst = 32'h8220000;
      44800: inst = 32'h10408000;
      44801: inst = 32'hc404a3b;
      44802: inst = 32'h8220000;
      44803: inst = 32'h10408000;
      44804: inst = 32'hc404a7d;
      44805: inst = 32'h8220000;
      44806: inst = 32'h10408000;
      44807: inst = 32'hc404a7e;
      44808: inst = 32'h8220000;
      44809: inst = 32'h10408000;
      44810: inst = 32'hc404a7f;
      44811: inst = 32'h8220000;
      44812: inst = 32'h10408000;
      44813: inst = 32'hc404a80;
      44814: inst = 32'h8220000;
      44815: inst = 32'h10408000;
      44816: inst = 32'hc404a81;
      44817: inst = 32'h8220000;
      44818: inst = 32'h10408000;
      44819: inst = 32'hc404a82;
      44820: inst = 32'h8220000;
      44821: inst = 32'h10408000;
      44822: inst = 32'hc404a83;
      44823: inst = 32'h8220000;
      44824: inst = 32'h10408000;
      44825: inst = 32'hc404a84;
      44826: inst = 32'h8220000;
      44827: inst = 32'h10408000;
      44828: inst = 32'hc404a85;
      44829: inst = 32'h8220000;
      44830: inst = 32'h10408000;
      44831: inst = 32'hc404a86;
      44832: inst = 32'h8220000;
      44833: inst = 32'h10408000;
      44834: inst = 32'hc404a87;
      44835: inst = 32'h8220000;
      44836: inst = 32'h10408000;
      44837: inst = 32'hc404a8a;
      44838: inst = 32'h8220000;
      44839: inst = 32'h10408000;
      44840: inst = 32'hc404a8b;
      44841: inst = 32'h8220000;
      44842: inst = 32'h10408000;
      44843: inst = 32'hc404a8c;
      44844: inst = 32'h8220000;
      44845: inst = 32'h10408000;
      44846: inst = 32'hc404a8d;
      44847: inst = 32'h8220000;
      44848: inst = 32'h10408000;
      44849: inst = 32'hc404a96;
      44850: inst = 32'h8220000;
      44851: inst = 32'h10408000;
      44852: inst = 32'hc404a97;
      44853: inst = 32'h8220000;
      44854: inst = 32'h10408000;
      44855: inst = 32'hc404a9a;
      44856: inst = 32'h8220000;
      44857: inst = 32'h10408000;
      44858: inst = 32'hc404a9b;
      44859: inst = 32'h8220000;
      44860: inst = 32'h10408000;
      44861: inst = 32'hc404add;
      44862: inst = 32'h8220000;
      44863: inst = 32'h10408000;
      44864: inst = 32'hc404ade;
      44865: inst = 32'h8220000;
      44866: inst = 32'h10408000;
      44867: inst = 32'hc404adf;
      44868: inst = 32'h8220000;
      44869: inst = 32'h10408000;
      44870: inst = 32'hc404aea;
      44871: inst = 32'h8220000;
      44872: inst = 32'h10408000;
      44873: inst = 32'hc404aeb;
      44874: inst = 32'h8220000;
      44875: inst = 32'h10408000;
      44876: inst = 32'hc404aec;
      44877: inst = 32'h8220000;
      44878: inst = 32'h10408000;
      44879: inst = 32'hc404aed;
      44880: inst = 32'h8220000;
      44881: inst = 32'h10408000;
      44882: inst = 32'hc404aee;
      44883: inst = 32'h8220000;
      44884: inst = 32'h10408000;
      44885: inst = 32'hc404af6;
      44886: inst = 32'h8220000;
      44887: inst = 32'h10408000;
      44888: inst = 32'hc404af7;
      44889: inst = 32'h8220000;
      44890: inst = 32'h10408000;
      44891: inst = 32'hc404afa;
      44892: inst = 32'h8220000;
      44893: inst = 32'h10408000;
      44894: inst = 32'hc404afb;
      44895: inst = 32'h8220000;
      44896: inst = 32'h10408000;
      44897: inst = 32'hc404b3d;
      44898: inst = 32'h8220000;
      44899: inst = 32'h10408000;
      44900: inst = 32'hc404b3e;
      44901: inst = 32'h8220000;
      44902: inst = 32'h10408000;
      44903: inst = 32'hc404b4a;
      44904: inst = 32'h8220000;
      44905: inst = 32'h10408000;
      44906: inst = 32'hc404b4c;
      44907: inst = 32'h8220000;
      44908: inst = 32'h10408000;
      44909: inst = 32'hc404b4d;
      44910: inst = 32'h8220000;
      44911: inst = 32'h10408000;
      44912: inst = 32'hc404b4e;
      44913: inst = 32'h8220000;
      44914: inst = 32'h10408000;
      44915: inst = 32'hc404b4f;
      44916: inst = 32'h8220000;
      44917: inst = 32'h10408000;
      44918: inst = 32'hc404b56;
      44919: inst = 32'h8220000;
      44920: inst = 32'h10408000;
      44921: inst = 32'hc404b57;
      44922: inst = 32'h8220000;
      44923: inst = 32'h10408000;
      44924: inst = 32'hc404b5a;
      44925: inst = 32'h8220000;
      44926: inst = 32'h10408000;
      44927: inst = 32'hc404b5b;
      44928: inst = 32'h8220000;
      44929: inst = 32'h10408000;
      44930: inst = 32'hc404b9d;
      44931: inst = 32'h8220000;
      44932: inst = 32'h10408000;
      44933: inst = 32'hc404b9e;
      44934: inst = 32'h8220000;
      44935: inst = 32'h10408000;
      44936: inst = 32'hc404ba0;
      44937: inst = 32'h8220000;
      44938: inst = 32'h10408000;
      44939: inst = 32'hc404ba1;
      44940: inst = 32'h8220000;
      44941: inst = 32'h10408000;
      44942: inst = 32'hc404ba2;
      44943: inst = 32'h8220000;
      44944: inst = 32'h10408000;
      44945: inst = 32'hc404ba3;
      44946: inst = 32'h8220000;
      44947: inst = 32'h10408000;
      44948: inst = 32'hc404ba4;
      44949: inst = 32'h8220000;
      44950: inst = 32'h10408000;
      44951: inst = 32'hc404ba5;
      44952: inst = 32'h8220000;
      44953: inst = 32'h10408000;
      44954: inst = 32'hc404baa;
      44955: inst = 32'h8220000;
      44956: inst = 32'h10408000;
      44957: inst = 32'hc404bab;
      44958: inst = 32'h8220000;
      44959: inst = 32'h10408000;
      44960: inst = 32'hc404bac;
      44961: inst = 32'h8220000;
      44962: inst = 32'h10408000;
      44963: inst = 32'hc404bad;
      44964: inst = 32'h8220000;
      44965: inst = 32'h10408000;
      44966: inst = 32'hc404bae;
      44967: inst = 32'h8220000;
      44968: inst = 32'h10408000;
      44969: inst = 32'hc404baf;
      44970: inst = 32'h8220000;
      44971: inst = 32'h10408000;
      44972: inst = 32'hc404bb0;
      44973: inst = 32'h8220000;
      44974: inst = 32'h10408000;
      44975: inst = 32'hc404bb6;
      44976: inst = 32'h8220000;
      44977: inst = 32'h10408000;
      44978: inst = 32'hc404bb7;
      44979: inst = 32'h8220000;
      44980: inst = 32'h10408000;
      44981: inst = 32'hc404bba;
      44982: inst = 32'h8220000;
      44983: inst = 32'h10408000;
      44984: inst = 32'hc404bbb;
      44985: inst = 32'h8220000;
      44986: inst = 32'h10408000;
      44987: inst = 32'hc404bfd;
      44988: inst = 32'h8220000;
      44989: inst = 32'h10408000;
      44990: inst = 32'hc404bfe;
      44991: inst = 32'h8220000;
      44992: inst = 32'h10408000;
      44993: inst = 32'hc404c00;
      44994: inst = 32'h8220000;
      44995: inst = 32'h10408000;
      44996: inst = 32'hc404c01;
      44997: inst = 32'h8220000;
      44998: inst = 32'h10408000;
      44999: inst = 32'hc404c02;
      45000: inst = 32'h8220000;
      45001: inst = 32'h10408000;
      45002: inst = 32'hc404c03;
      45003: inst = 32'h8220000;
      45004: inst = 32'h10408000;
      45005: inst = 32'hc404c04;
      45006: inst = 32'h8220000;
      45007: inst = 32'h10408000;
      45008: inst = 32'hc404c05;
      45009: inst = 32'h8220000;
      45010: inst = 32'h10408000;
      45011: inst = 32'hc404c0a;
      45012: inst = 32'h8220000;
      45013: inst = 32'h10408000;
      45014: inst = 32'hc404c0b;
      45015: inst = 32'h8220000;
      45016: inst = 32'h10408000;
      45017: inst = 32'hc404c0c;
      45018: inst = 32'h8220000;
      45019: inst = 32'h10408000;
      45020: inst = 32'hc404c0e;
      45021: inst = 32'h8220000;
      45022: inst = 32'h10408000;
      45023: inst = 32'hc404c0f;
      45024: inst = 32'h8220000;
      45025: inst = 32'h10408000;
      45026: inst = 32'hc404c10;
      45027: inst = 32'h8220000;
      45028: inst = 32'h10408000;
      45029: inst = 32'hc404c11;
      45030: inst = 32'h8220000;
      45031: inst = 32'h10408000;
      45032: inst = 32'hc404c16;
      45033: inst = 32'h8220000;
      45034: inst = 32'h10408000;
      45035: inst = 32'hc404c17;
      45036: inst = 32'h8220000;
      45037: inst = 32'h10408000;
      45038: inst = 32'hc404c1a;
      45039: inst = 32'h8220000;
      45040: inst = 32'h10408000;
      45041: inst = 32'hc404c1b;
      45042: inst = 32'h8220000;
      45043: inst = 32'h10408000;
      45044: inst = 32'hc404c5d;
      45045: inst = 32'h8220000;
      45046: inst = 32'h10408000;
      45047: inst = 32'hc404c5e;
      45048: inst = 32'h8220000;
      45049: inst = 32'h10408000;
      45050: inst = 32'hc404c6a;
      45051: inst = 32'h8220000;
      45052: inst = 32'h10408000;
      45053: inst = 32'hc404c6b;
      45054: inst = 32'h8220000;
      45055: inst = 32'h10408000;
      45056: inst = 32'hc404c6c;
      45057: inst = 32'h8220000;
      45058: inst = 32'h10408000;
      45059: inst = 32'hc404c6d;
      45060: inst = 32'h8220000;
      45061: inst = 32'h10408000;
      45062: inst = 32'hc404c6e;
      45063: inst = 32'h8220000;
      45064: inst = 32'h10408000;
      45065: inst = 32'hc404c6f;
      45066: inst = 32'h8220000;
      45067: inst = 32'h10408000;
      45068: inst = 32'hc404c70;
      45069: inst = 32'h8220000;
      45070: inst = 32'h10408000;
      45071: inst = 32'hc404c71;
      45072: inst = 32'h8220000;
      45073: inst = 32'h10408000;
      45074: inst = 32'hc404c72;
      45075: inst = 32'h8220000;
      45076: inst = 32'h10408000;
      45077: inst = 32'hc404c76;
      45078: inst = 32'h8220000;
      45079: inst = 32'h10408000;
      45080: inst = 32'hc404c77;
      45081: inst = 32'h8220000;
      45082: inst = 32'h10408000;
      45083: inst = 32'hc404c7a;
      45084: inst = 32'h8220000;
      45085: inst = 32'h10408000;
      45086: inst = 32'hc404c7b;
      45087: inst = 32'h8220000;
      45088: inst = 32'h10408000;
      45089: inst = 32'hc404cbd;
      45090: inst = 32'h8220000;
      45091: inst = 32'h10408000;
      45092: inst = 32'hc404cbe;
      45093: inst = 32'h8220000;
      45094: inst = 32'h10408000;
      45095: inst = 32'hc404cca;
      45096: inst = 32'h8220000;
      45097: inst = 32'h10408000;
      45098: inst = 32'hc404ccb;
      45099: inst = 32'h8220000;
      45100: inst = 32'h10408000;
      45101: inst = 32'hc404cd0;
      45102: inst = 32'h8220000;
      45103: inst = 32'h10408000;
      45104: inst = 32'hc404cd1;
      45105: inst = 32'h8220000;
      45106: inst = 32'h10408000;
      45107: inst = 32'hc404cd2;
      45108: inst = 32'h8220000;
      45109: inst = 32'h10408000;
      45110: inst = 32'hc404cd3;
      45111: inst = 32'h8220000;
      45112: inst = 32'h10408000;
      45113: inst = 32'hc404cd6;
      45114: inst = 32'h8220000;
      45115: inst = 32'h10408000;
      45116: inst = 32'hc404cd7;
      45117: inst = 32'h8220000;
      45118: inst = 32'h10408000;
      45119: inst = 32'hc404cda;
      45120: inst = 32'h8220000;
      45121: inst = 32'h10408000;
      45122: inst = 32'hc404cdb;
      45123: inst = 32'h8220000;
      45124: inst = 32'h10408000;
      45125: inst = 32'hc404cdc;
      45126: inst = 32'h8220000;
      45127: inst = 32'h10408000;
      45128: inst = 32'hc404cdd;
      45129: inst = 32'h8220000;
      45130: inst = 32'h10408000;
      45131: inst = 32'hc404cde;
      45132: inst = 32'h8220000;
      45133: inst = 32'h10408000;
      45134: inst = 32'hc404cdf;
      45135: inst = 32'h8220000;
      45136: inst = 32'h10408000;
      45137: inst = 32'hc404ce0;
      45138: inst = 32'h8220000;
      45139: inst = 32'h10408000;
      45140: inst = 32'hc404ce1;
      45141: inst = 32'h8220000;
      45142: inst = 32'h10408000;
      45143: inst = 32'hc404ce2;
      45144: inst = 32'h8220000;
      45145: inst = 32'h10408000;
      45146: inst = 32'hc404d1d;
      45147: inst = 32'h8220000;
      45148: inst = 32'h10408000;
      45149: inst = 32'hc404d1e;
      45150: inst = 32'h8220000;
      45151: inst = 32'h10408000;
      45152: inst = 32'hc404d2a;
      45153: inst = 32'h8220000;
      45154: inst = 32'h10408000;
      45155: inst = 32'hc404d2b;
      45156: inst = 32'h8220000;
      45157: inst = 32'h10408000;
      45158: inst = 32'hc404d31;
      45159: inst = 32'h8220000;
      45160: inst = 32'h10408000;
      45161: inst = 32'hc404d32;
      45162: inst = 32'h8220000;
      45163: inst = 32'h10408000;
      45164: inst = 32'hc404d33;
      45165: inst = 32'h8220000;
      45166: inst = 32'h10408000;
      45167: inst = 32'hc404d34;
      45168: inst = 32'h8220000;
      45169: inst = 32'h10408000;
      45170: inst = 32'hc404d36;
      45171: inst = 32'h8220000;
      45172: inst = 32'h10408000;
      45173: inst = 32'hc404d37;
      45174: inst = 32'h8220000;
      45175: inst = 32'h10408000;
      45176: inst = 32'hc404d3a;
      45177: inst = 32'h8220000;
      45178: inst = 32'h10408000;
      45179: inst = 32'hc404d3b;
      45180: inst = 32'h8220000;
      45181: inst = 32'h10408000;
      45182: inst = 32'hc404d3c;
      45183: inst = 32'h8220000;
      45184: inst = 32'h10408000;
      45185: inst = 32'hc404d3d;
      45186: inst = 32'h8220000;
      45187: inst = 32'h10408000;
      45188: inst = 32'hc404d3e;
      45189: inst = 32'h8220000;
      45190: inst = 32'h10408000;
      45191: inst = 32'hc404d3f;
      45192: inst = 32'h8220000;
      45193: inst = 32'h10408000;
      45194: inst = 32'hc404d40;
      45195: inst = 32'h8220000;
      45196: inst = 32'h10408000;
      45197: inst = 32'hc404d41;
      45198: inst = 32'h8220000;
      45199: inst = 32'h10408000;
      45200: inst = 32'hc404d42;
      45201: inst = 32'h8220000;
      45202: inst = 32'h58000000;
      45203: inst = 32'h10608000;
      45204: inst = 32'hc600000;
      45205: inst = 32'hc20aaaa;
      45206: inst = 32'h4c210000;
      45207: inst = 32'h8230000;
      45208: inst = 32'h104000fe;
      45209: inst = 32'hc40502a;
      45210: inst = 32'h30420001;
      45211: inst = 32'h13e00000;
      45212: inst = 32'hfe0b09a;
      45213: inst = 32'h1c400000;
      45214: inst = 32'h5be00000;
      45215: inst = 32'h13e00000;
      45216: inst = 32'hfe0b096;
      45217: inst = 32'h5be00000;
    endcase
  end
endmodule
